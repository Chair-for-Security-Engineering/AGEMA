module Reg1(x, y);
 input [275:0] x;
 output [274:0] y;

  assign y[0] = x[145];
  register_stage #(.WIDTH(274)) inst_0(.clk(x[136]), .D({x[146],x[147],x[137],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[185],x[186],x[187],x[188],x[189],x[190],x[191],x[192],x[193],x[194],x[195],x[196],x[197],x[198],x[199],x[200],x[201],x[202],x[203],x[204],x[205],x[206],x[207],x[208],x[209],x[210],x[211],x[212],x[213],x[214],x[215],x[216],x[217],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[238],x[239],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[247],x[248],x[249],x[250],x[251],x[252],x[253],x[254],x[255],x[256],x[257],x[258],x[259],x[260],x[261],x[262],x[263],x[264],x[265],x[266],x[267],x[268],x[269],x[270],x[271],x[272],x[273],x[274],x[275]}), .Q({y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194],y[195],y[196],y[197],y[198],y[199],y[200],y[201],y[202],y[203],y[204],y[205],y[206],y[207],y[208],y[209],y[210],y[211],y[212],y[213],y[214],y[215],y[216],y[217],y[218],y[219],y[220],y[221],y[222],y[223],y[224],y[225],y[226],y[227],y[228],y[229],y[230],y[231],y[232],y[233],y[234],y[235],y[236],y[237],y[238],y[239],y[240],y[241],y[242],y[243],y[244],y[245],y[246],y[247],y[248],y[249],y[250],y[251],y[252],y[253],y[254],y[255],y[256],y[257],y[258],y[259],y[260],y[261],y[262],y[263],y[264],y[265],y[266],y[267],y[268],y[269],y[270],y[271],y[272],y[273],y[274]}));
endmodule

module Reg2(x, y);
 input [550:0] x;
 output [549:0] y;

  assign y[0] = x[289];
  assign y[1] = x[290];
  register_stage #(.WIDTH(548)) inst_0(.clk(x[272]), .D({x[291],x[292],x[293],x[294],x[273],x[274],x[256],x[257],x[258],x[259],x[260],x[261],x[262],x[263],x[264],x[265],x[266],x[267],x[268],x[269],x[270],x[271],x[275],x[276],x[277],x[278],x[279],x[280],x[281],x[282],x[283],x[284],x[285],x[286],x[287],x[288],x[0],x[1],x[2],x[3],x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[185],x[186],x[187],x[188],x[189],x[190],x[191],x[192],x[193],x[194],x[195],x[196],x[197],x[198],x[199],x[200],x[201],x[202],x[203],x[204],x[205],x[206],x[207],x[208],x[209],x[210],x[211],x[212],x[213],x[214],x[215],x[216],x[217],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[238],x[239],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[247],x[248],x[249],x[250],x[251],x[252],x[253],x[254],x[255],x[295],x[296],x[297],x[298],x[299],x[300],x[301],x[302],x[303],x[304],x[305],x[306],x[307],x[308],x[309],x[310],x[311],x[312],x[313],x[314],x[315],x[316],x[317],x[318],x[319],x[320],x[321],x[322],x[323],x[324],x[325],x[326],x[327],x[328],x[329],x[330],x[331],x[332],x[333],x[334],x[335],x[336],x[337],x[338],x[339],x[340],x[341],x[342],x[343],x[344],x[345],x[346],x[347],x[348],x[349],x[350],x[351],x[352],x[353],x[354],x[355],x[356],x[357],x[358],x[359],x[360],x[361],x[362],x[363],x[364],x[365],x[366],x[367],x[368],x[369],x[370],x[371],x[372],x[373],x[374],x[375],x[376],x[377],x[378],x[379],x[380],x[381],x[382],x[383],x[384],x[385],x[386],x[387],x[388],x[389],x[390],x[391],x[392],x[393],x[394],x[395],x[396],x[397],x[398],x[399],x[400],x[401],x[402],x[403],x[404],x[405],x[406],x[407],x[408],x[409],x[410],x[411],x[412],x[413],x[414],x[415],x[416],x[417],x[418],x[419],x[420],x[421],x[422],x[423],x[424],x[425],x[426],x[427],x[428],x[429],x[430],x[431],x[432],x[433],x[434],x[435],x[436],x[437],x[438],x[439],x[440],x[441],x[442],x[443],x[444],x[445],x[446],x[447],x[448],x[449],x[450],x[451],x[452],x[453],x[454],x[455],x[456],x[457],x[458],x[459],x[460],x[461],x[462],x[463],x[464],x[465],x[466],x[467],x[468],x[469],x[470],x[471],x[472],x[473],x[474],x[475],x[476],x[477],x[478],x[479],x[480],x[481],x[482],x[483],x[484],x[485],x[486],x[487],x[488],x[489],x[490],x[491],x[492],x[493],x[494],x[495],x[496],x[497],x[498],x[499],x[500],x[501],x[502],x[503],x[504],x[505],x[506],x[507],x[508],x[509],x[510],x[511],x[512],x[513],x[514],x[515],x[516],x[517],x[518],x[519],x[520],x[521],x[522],x[523],x[524],x[525],x[526],x[527],x[528],x[529],x[530],x[531],x[532],x[533],x[534],x[535],x[536],x[537],x[538],x[539],x[540],x[541],x[542],x[543],x[544],x[545],x[546],x[547],x[548],x[549],x[550]}), .Q({y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194],y[195],y[196],y[197],y[198],y[199],y[200],y[201],y[202],y[203],y[204],y[205],y[206],y[207],y[208],y[209],y[210],y[211],y[212],y[213],y[214],y[215],y[216],y[217],y[218],y[219],y[220],y[221],y[222],y[223],y[224],y[225],y[226],y[227],y[228],y[229],y[230],y[231],y[232],y[233],y[234],y[235],y[236],y[237],y[238],y[239],y[240],y[241],y[242],y[243],y[244],y[245],y[246],y[247],y[248],y[249],y[250],y[251],y[252],y[253],y[254],y[255],y[256],y[257],y[258],y[259],y[260],y[261],y[262],y[263],y[264],y[265],y[266],y[267],y[268],y[269],y[270],y[271],y[272],y[273],y[274],y[275],y[276],y[277],y[278],y[279],y[280],y[281],y[282],y[283],y[284],y[285],y[286],y[287],y[288],y[289],y[290],y[291],y[292],y[293],y[294],y[295],y[296],y[297],y[298],y[299],y[300],y[301],y[302],y[303],y[304],y[305],y[306],y[307],y[308],y[309],y[310],y[311],y[312],y[313],y[314],y[315],y[316],y[317],y[318],y[319],y[320],y[321],y[322],y[323],y[324],y[325],y[326],y[327],y[328],y[329],y[330],y[331],y[332],y[333],y[334],y[335],y[336],y[337],y[338],y[339],y[340],y[341],y[342],y[343],y[344],y[345],y[346],y[347],y[348],y[349],y[350],y[351],y[352],y[353],y[354],y[355],y[356],y[357],y[358],y[359],y[360],y[361],y[362],y[363],y[364],y[365],y[366],y[367],y[368],y[369],y[370],y[371],y[372],y[373],y[374],y[375],y[376],y[377],y[378],y[379],y[380],y[381],y[382],y[383],y[384],y[385],y[386],y[387],y[388],y[389],y[390],y[391],y[392],y[393],y[394],y[395],y[396],y[397],y[398],y[399],y[400],y[401],y[402],y[403],y[404],y[405],y[406],y[407],y[408],y[409],y[410],y[411],y[412],y[413],y[414],y[415],y[416],y[417],y[418],y[419],y[420],y[421],y[422],y[423],y[424],y[425],y[426],y[427],y[428],y[429],y[430],y[431],y[432],y[433],y[434],y[435],y[436],y[437],y[438],y[439],y[440],y[441],y[442],y[443],y[444],y[445],y[446],y[447],y[448],y[449],y[450],y[451],y[452],y[453],y[454],y[455],y[456],y[457],y[458],y[459],y[460],y[461],y[462],y[463],y[464],y[465],y[466],y[467],y[468],y[469],y[470],y[471],y[472],y[473],y[474],y[475],y[476],y[477],y[478],y[479],y[480],y[481],y[482],y[483],y[484],y[485],y[486],y[487],y[488],y[489],y[490],y[491],y[492],y[493],y[494],y[495],y[496],y[497],y[498],y[499],y[500],y[501],y[502],y[503],y[504],y[505],y[506],y[507],y[508],y[509],y[510],y[511],y[512],y[513],y[514],y[515],y[516],y[517],y[518],y[519],y[520],y[521],y[522],y[523],y[524],y[525],y[526],y[527],y[528],y[529],y[530],y[531],y[532],y[533],y[534],y[535],y[536],y[537],y[538],y[539],y[540],y[541],y[542],y[543],y[544],y[545],y[546],y[547],y[548],y[549]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx6(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx12(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx13(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx195(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx196(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx197(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx198(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx199(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx200(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx201(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx202(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx203(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx204(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx205(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx206(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx207(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx208(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx209(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx210(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx211(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx212(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx213(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx214(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx215(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx216(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx217(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx218(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx219(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx220(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx221(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx222(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx223(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx224(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx225(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx226(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx227(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx228(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx229(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx230(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx231(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx232(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx233(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx234(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx235(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx236(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx237(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx238(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx239(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx240(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx241(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx242(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx243(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx244(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx245(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx246(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx247(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx248(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx249(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx250(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx251(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx252(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx253(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx254(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx255(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx256(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx257(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx258(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx259(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx260(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx261(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx262(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx263(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx264(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx265(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx266(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx267(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx268(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx269(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx270(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx271(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx272(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx273(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx274(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx275(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx276(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx277(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx278(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx279(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx280(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx281(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx282(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx283(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx284(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx285(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx286(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx287(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx288(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx289(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx290(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx291(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx292(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx293(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx294(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx295(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx296(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx297(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx298(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx299(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx300(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx301(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx302(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx303(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx304(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx305(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx306(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx307(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx308(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx309(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx310(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx311(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx312(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx313(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx314(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx315(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx316(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx317(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx318(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx319(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx320(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx321(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx322(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx323(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx324(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx325(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx326(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx327(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx328(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx329(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx330(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx331(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx332(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx333(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx334(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx335(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx336(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx337(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx338(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx339(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx340(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx341(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx342(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx343(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx344(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx345(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx346(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx347(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx348(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx349(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx350(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx351(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx352(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx353(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx354(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx355(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx356(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx357(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx358(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx359(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx360(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx361(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx362(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx363(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx364(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx365(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx366(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx367(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx368(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx369(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx370(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx371(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx372(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx373(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx374(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx375(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx376(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx377(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx378(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx379(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx380(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx381(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx382(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx383(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx384(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx385(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx386(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx387(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx388(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx389(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx390(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx391(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx392(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx393(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx394(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx395(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx396(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx397(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx398(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx399(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx400(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx401(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx402(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx403(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx404(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx405(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx406(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx407(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx408(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx409(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx410(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx411(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx412(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx413(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx414(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx415(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx416(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx417(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx418(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx419(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx420(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx421(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx422(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx423(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx424(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx425(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx426(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx427(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx428(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx429(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx430(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx431(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx432(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx433(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx434(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx435(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx436(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx437(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx438(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx439(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx440(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx441(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx442(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx443(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx444(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx445(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx446(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx447(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx448(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx449(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx450(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx451(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx452(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx453(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx454(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx455(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx456(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx457(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx458(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx459(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx460(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx461(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx462(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx463(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx464(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx465(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx466(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx467(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx468(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx469(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx470(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx471(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx472(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx473(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx474(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx475(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx476(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx477(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx478(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx479(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx480(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx481(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx482(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx483(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx484(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx485(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx486(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx487(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx488(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx489(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx490(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx491(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx492(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx493(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx494(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx495(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx496(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx497(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx498(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx499(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx500(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx501(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx502(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx503(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx504(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx505(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx506(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx507(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx508(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx509(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx510(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx511(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx512(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx513(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx514(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx515(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx516(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx517(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx518(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx519(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx520(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx521(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx522(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx523(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx524(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx525(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx526(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx527(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx528(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx529(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx530(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx531(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx532(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx533(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx534(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx535(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx536(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx537(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx538(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx539(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx540(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx541(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx542(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx543(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx544(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx545(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx546(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx547(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx548(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx549(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [824:0] x;
 output [549:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx4 Fx4_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx5 Fx5_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx6 Fx6_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx7 Fx7_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx11 Fx11_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx12 Fx12_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx13 Fx13_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx14 Fx14_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx18 Fx18_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx19 Fx19_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx20 Fx20_inst(.x({x[31], x[30]}), .y(y[20]));
  Fx21 Fx21_inst(.x({x[32], x[30]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[34], x[33]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[35], x[33]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[37], x[36]}), .y(y[24]));
  Fx25 Fx25_inst(.x({x[38], x[36]}), .y(y[25]));
  Fx26 Fx26_inst(.x({x[40], x[39]}), .y(y[26]));
  Fx27 Fx27_inst(.x({x[41], x[39]}), .y(y[27]));
  Fx28 Fx28_inst(.x({x[43], x[42]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[44], x[42]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[46], x[45]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[47], x[45]}), .y(y[31]));
  Fx32 Fx32_inst(.x({x[49], x[48]}), .y(y[32]));
  Fx33 Fx33_inst(.x({x[50], x[48]}), .y(y[33]));
  Fx34 Fx34_inst(.x({x[52], x[51]}), .y(y[34]));
  Fx35 Fx35_inst(.x({x[53], x[51]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[55], x[54]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[56], x[54]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[58], x[57]}), .y(y[38]));
  Fx39 Fx39_inst(.x({x[59], x[57]}), .y(y[39]));
  Fx40 Fx40_inst(.x({x[61], x[60]}), .y(y[40]));
  Fx41 Fx41_inst(.x({x[62], x[60]}), .y(y[41]));
  Fx42 Fx42_inst(.x({x[64], x[63]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[65], x[63]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[67], x[66]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[68], x[66]}), .y(y[45]));
  Fx46 Fx46_inst(.x({x[70], x[69]}), .y(y[46]));
  Fx47 Fx47_inst(.x({x[71], x[69]}), .y(y[47]));
  Fx48 Fx48_inst(.x({x[73], x[72]}), .y(y[48]));
  Fx49 Fx49_inst(.x({x[74], x[72]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[76], x[75]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[77], x[75]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[79], x[78]}), .y(y[52]));
  Fx53 Fx53_inst(.x({x[80], x[78]}), .y(y[53]));
  Fx54 Fx54_inst(.x({x[82], x[81]}), .y(y[54]));
  Fx55 Fx55_inst(.x({x[83], x[81]}), .y(y[55]));
  Fx56 Fx56_inst(.x({x[85], x[84]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[86], x[84]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[88], x[87]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[89], x[87]}), .y(y[59]));
  Fx60 Fx60_inst(.x({x[91], x[90]}), .y(y[60]));
  Fx61 Fx61_inst(.x({x[92], x[90]}), .y(y[61]));
  Fx62 Fx62_inst(.x({x[94], x[93]}), .y(y[62]));
  Fx63 Fx63_inst(.x({x[95], x[93]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[97], x[96]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[98], x[96]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[100], x[99]}), .y(y[66]));
  Fx67 Fx67_inst(.x({x[101], x[99]}), .y(y[67]));
  Fx68 Fx68_inst(.x({x[103], x[102]}), .y(y[68]));
  Fx69 Fx69_inst(.x({x[104], x[102]}), .y(y[69]));
  Fx70 Fx70_inst(.x({x[106], x[105]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[107], x[105]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[109], x[108]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[110], x[108]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[112], x[111]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[113], x[111]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[115], x[114]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[116], x[114]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[118], x[117]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[119], x[117]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[121], x[120]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[122], x[120]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[124], x[123]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[125], x[123]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[127], x[126]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[128], x[126]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[130], x[129]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[131], x[129]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[133], x[132]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[134], x[132]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[136], x[135]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[137], x[135]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[139], x[138]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[140], x[138]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[142], x[141]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[143], x[141]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[145], x[144]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[146], x[144]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[148], x[147]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[149], x[147]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[151], x[150]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[152], x[150]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[154], x[153]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[155], x[153]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[157], x[156]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[158], x[156]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[160], x[159]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[161], x[159]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[163], x[162]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[164], x[162]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[166], x[165]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[167], x[165]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[169], x[168]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[170], x[168]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[172], x[171]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[173], x[171]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[175], x[174]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[176], x[174]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[178], x[177]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[179], x[177]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[181], x[180]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[182], x[180]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[184], x[183]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[185], x[183]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[187], x[186]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[188], x[186]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[190], x[189]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[191], x[189]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[193], x[192]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[194], x[192]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[196], x[195]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[197], x[195]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[199], x[198]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[200], x[198]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[202], x[201]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[203], x[201]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[205], x[204]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[206], x[204]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[208], x[207]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[209], x[207]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[211], x[210]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[212], x[210]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[214], x[213]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[215], x[213]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[217], x[216]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[218], x[216]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[220], x[219]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[221], x[219]}), .y(y[147]));
  Fx148 Fx148_inst(.x({x[223], x[222]}), .y(y[148]));
  Fx149 Fx149_inst(.x({x[224], x[222]}), .y(y[149]));
  Fx150 Fx150_inst(.x({x[226], x[225]}), .y(y[150]));
  Fx151 Fx151_inst(.x({x[227], x[225]}), .y(y[151]));
  Fx152 Fx152_inst(.x({x[229], x[228]}), .y(y[152]));
  Fx153 Fx153_inst(.x({x[230], x[228]}), .y(y[153]));
  Fx154 Fx154_inst(.x({x[232], x[231]}), .y(y[154]));
  Fx155 Fx155_inst(.x({x[233], x[231]}), .y(y[155]));
  Fx156 Fx156_inst(.x({x[235], x[234]}), .y(y[156]));
  Fx157 Fx157_inst(.x({x[236], x[234]}), .y(y[157]));
  Fx158 Fx158_inst(.x({x[238], x[237]}), .y(y[158]));
  Fx159 Fx159_inst(.x({x[239], x[237]}), .y(y[159]));
  Fx160 Fx160_inst(.x({x[241], x[240]}), .y(y[160]));
  Fx161 Fx161_inst(.x({x[242], x[240]}), .y(y[161]));
  Fx162 Fx162_inst(.x({x[244], x[243]}), .y(y[162]));
  Fx163 Fx163_inst(.x({x[245], x[243]}), .y(y[163]));
  Fx164 Fx164_inst(.x({x[247], x[246]}), .y(y[164]));
  Fx165 Fx165_inst(.x({x[248], x[246]}), .y(y[165]));
  Fx166 Fx166_inst(.x({x[250], x[249]}), .y(y[166]));
  Fx167 Fx167_inst(.x({x[251], x[249]}), .y(y[167]));
  Fx168 Fx168_inst(.x({x[253], x[252]}), .y(y[168]));
  Fx169 Fx169_inst(.x({x[254], x[252]}), .y(y[169]));
  Fx170 Fx170_inst(.x({x[256], x[255]}), .y(y[170]));
  Fx171 Fx171_inst(.x({x[257], x[255]}), .y(y[171]));
  Fx172 Fx172_inst(.x({x[259], x[258]}), .y(y[172]));
  Fx173 Fx173_inst(.x({x[260], x[258]}), .y(y[173]));
  Fx174 Fx174_inst(.x({x[262], x[261]}), .y(y[174]));
  Fx175 Fx175_inst(.x({x[263], x[261]}), .y(y[175]));
  Fx176 Fx176_inst(.x({x[265], x[264]}), .y(y[176]));
  Fx177 Fx177_inst(.x({x[266], x[264]}), .y(y[177]));
  Fx178 Fx178_inst(.x({x[268], x[267]}), .y(y[178]));
  Fx179 Fx179_inst(.x({x[269], x[267]}), .y(y[179]));
  Fx180 Fx180_inst(.x({x[271], x[270]}), .y(y[180]));
  Fx181 Fx181_inst(.x({x[272], x[270]}), .y(y[181]));
  Fx182 Fx182_inst(.x({x[274], x[273]}), .y(y[182]));
  Fx183 Fx183_inst(.x({x[275], x[273]}), .y(y[183]));
  Fx184 Fx184_inst(.x({x[277], x[276]}), .y(y[184]));
  Fx185 Fx185_inst(.x({x[278], x[276]}), .y(y[185]));
  Fx186 Fx186_inst(.x({x[280], x[279]}), .y(y[186]));
  Fx187 Fx187_inst(.x({x[281], x[279]}), .y(y[187]));
  Fx188 Fx188_inst(.x({x[283], x[282]}), .y(y[188]));
  Fx189 Fx189_inst(.x({x[284], x[282]}), .y(y[189]));
  Fx190 Fx190_inst(.x({x[286], x[285]}), .y(y[190]));
  Fx191 Fx191_inst(.x({x[287], x[285]}), .y(y[191]));
  Fx192 Fx192_inst(.x({x[289], x[288]}), .y(y[192]));
  Fx193 Fx193_inst(.x({x[290], x[288]}), .y(y[193]));
  Fx194 Fx194_inst(.x({x[292], x[291]}), .y(y[194]));
  Fx195 Fx195_inst(.x({x[293], x[291]}), .y(y[195]));
  Fx196 Fx196_inst(.x({x[295], x[294]}), .y(y[196]));
  Fx197 Fx197_inst(.x({x[296], x[294]}), .y(y[197]));
  Fx198 Fx198_inst(.x({x[298], x[297]}), .y(y[198]));
  Fx199 Fx199_inst(.x({x[299], x[297]}), .y(y[199]));
  Fx200 Fx200_inst(.x({x[301], x[300]}), .y(y[200]));
  Fx201 Fx201_inst(.x({x[302], x[300]}), .y(y[201]));
  Fx202 Fx202_inst(.x({x[304], x[303]}), .y(y[202]));
  Fx203 Fx203_inst(.x({x[305], x[303]}), .y(y[203]));
  Fx204 Fx204_inst(.x({x[307], x[306]}), .y(y[204]));
  Fx205 Fx205_inst(.x({x[308], x[306]}), .y(y[205]));
  Fx206 Fx206_inst(.x({x[310], x[309]}), .y(y[206]));
  Fx207 Fx207_inst(.x({x[311], x[309]}), .y(y[207]));
  Fx208 Fx208_inst(.x({x[313], x[312]}), .y(y[208]));
  Fx209 Fx209_inst(.x({x[314], x[312]}), .y(y[209]));
  Fx210 Fx210_inst(.x({x[316], x[315]}), .y(y[210]));
  Fx211 Fx211_inst(.x({x[317], x[315]}), .y(y[211]));
  Fx212 Fx212_inst(.x({x[319], x[318]}), .y(y[212]));
  Fx213 Fx213_inst(.x({x[320], x[318]}), .y(y[213]));
  Fx214 Fx214_inst(.x({x[322], x[321]}), .y(y[214]));
  Fx215 Fx215_inst(.x({x[323], x[321]}), .y(y[215]));
  Fx216 Fx216_inst(.x({x[325], x[324]}), .y(y[216]));
  Fx217 Fx217_inst(.x({x[326], x[324]}), .y(y[217]));
  Fx218 Fx218_inst(.x({x[328], x[327]}), .y(y[218]));
  Fx219 Fx219_inst(.x({x[329], x[327]}), .y(y[219]));
  Fx220 Fx220_inst(.x({x[331], x[330]}), .y(y[220]));
  Fx221 Fx221_inst(.x({x[332], x[330]}), .y(y[221]));
  Fx222 Fx222_inst(.x({x[334], x[333]}), .y(y[222]));
  Fx223 Fx223_inst(.x({x[335], x[333]}), .y(y[223]));
  Fx224 Fx224_inst(.x({x[337], x[336]}), .y(y[224]));
  Fx225 Fx225_inst(.x({x[338], x[336]}), .y(y[225]));
  Fx226 Fx226_inst(.x({x[340], x[339]}), .y(y[226]));
  Fx227 Fx227_inst(.x({x[341], x[339]}), .y(y[227]));
  Fx228 Fx228_inst(.x({x[343], x[342]}), .y(y[228]));
  Fx229 Fx229_inst(.x({x[344], x[342]}), .y(y[229]));
  Fx230 Fx230_inst(.x({x[346], x[345]}), .y(y[230]));
  Fx231 Fx231_inst(.x({x[347], x[345]}), .y(y[231]));
  Fx232 Fx232_inst(.x({x[349], x[348]}), .y(y[232]));
  Fx233 Fx233_inst(.x({x[350], x[348]}), .y(y[233]));
  Fx234 Fx234_inst(.x({x[352], x[351]}), .y(y[234]));
  Fx235 Fx235_inst(.x({x[353], x[351]}), .y(y[235]));
  Fx236 Fx236_inst(.x({x[355], x[354]}), .y(y[236]));
  Fx237 Fx237_inst(.x({x[356], x[354]}), .y(y[237]));
  Fx238 Fx238_inst(.x({x[358], x[357]}), .y(y[238]));
  Fx239 Fx239_inst(.x({x[359], x[357]}), .y(y[239]));
  Fx240 Fx240_inst(.x({x[361], x[360]}), .y(y[240]));
  Fx241 Fx241_inst(.x({x[362], x[360]}), .y(y[241]));
  Fx242 Fx242_inst(.x({x[364], x[363]}), .y(y[242]));
  Fx243 Fx243_inst(.x({x[365], x[363]}), .y(y[243]));
  Fx244 Fx244_inst(.x({x[367], x[366]}), .y(y[244]));
  Fx245 Fx245_inst(.x({x[368], x[366]}), .y(y[245]));
  Fx246 Fx246_inst(.x({x[370], x[369]}), .y(y[246]));
  Fx247 Fx247_inst(.x({x[371], x[369]}), .y(y[247]));
  Fx248 Fx248_inst(.x({x[373], x[372]}), .y(y[248]));
  Fx249 Fx249_inst(.x({x[374], x[372]}), .y(y[249]));
  Fx250 Fx250_inst(.x({x[376], x[375]}), .y(y[250]));
  Fx251 Fx251_inst(.x({x[377], x[375]}), .y(y[251]));
  Fx252 Fx252_inst(.x({x[379], x[378]}), .y(y[252]));
  Fx253 Fx253_inst(.x({x[380], x[378]}), .y(y[253]));
  Fx254 Fx254_inst(.x({x[382], x[381]}), .y(y[254]));
  Fx255 Fx255_inst(.x({x[383], x[381]}), .y(y[255]));
  Fx256 Fx256_inst(.x({x[385], x[384]}), .y(y[256]));
  Fx257 Fx257_inst(.x({x[386], x[384]}), .y(y[257]));
  Fx258 Fx258_inst(.x({x[388], x[387]}), .y(y[258]));
  Fx259 Fx259_inst(.x({x[389], x[387]}), .y(y[259]));
  Fx260 Fx260_inst(.x({x[391], x[390]}), .y(y[260]));
  Fx261 Fx261_inst(.x({x[392], x[390]}), .y(y[261]));
  Fx262 Fx262_inst(.x({x[394], x[393]}), .y(y[262]));
  Fx263 Fx263_inst(.x({x[395], x[393]}), .y(y[263]));
  Fx264 Fx264_inst(.x({x[397], x[396]}), .y(y[264]));
  Fx265 Fx265_inst(.x({x[398], x[396]}), .y(y[265]));
  Fx266 Fx266_inst(.x({x[400], x[399]}), .y(y[266]));
  Fx267 Fx267_inst(.x({x[401], x[399]}), .y(y[267]));
  Fx268 Fx268_inst(.x({x[403], x[402]}), .y(y[268]));
  Fx269 Fx269_inst(.x({x[404], x[402]}), .y(y[269]));
  Fx270 Fx270_inst(.x({x[406], x[405]}), .y(y[270]));
  Fx271 Fx271_inst(.x({x[407], x[405]}), .y(y[271]));
  Fx272 Fx272_inst(.x({x[409], x[408]}), .y(y[272]));
  Fx273 Fx273_inst(.x({x[410], x[408]}), .y(y[273]));
  Fx274 Fx274_inst(.x({x[412], x[411]}), .y(y[274]));
  Fx275 Fx275_inst(.x({x[413], x[411]}), .y(y[275]));
  Fx276 Fx276_inst(.x({x[415], x[414]}), .y(y[276]));
  Fx277 Fx277_inst(.x({x[416], x[414]}), .y(y[277]));
  Fx278 Fx278_inst(.x({x[418], x[417]}), .y(y[278]));
  Fx279 Fx279_inst(.x({x[419], x[417]}), .y(y[279]));
  Fx280 Fx280_inst(.x({x[421], x[420]}), .y(y[280]));
  Fx281 Fx281_inst(.x({x[422], x[420]}), .y(y[281]));
  Fx282 Fx282_inst(.x({x[424], x[423]}), .y(y[282]));
  Fx283 Fx283_inst(.x({x[425], x[423]}), .y(y[283]));
  Fx284 Fx284_inst(.x({x[427], x[426]}), .y(y[284]));
  Fx285 Fx285_inst(.x({x[428], x[426]}), .y(y[285]));
  Fx286 Fx286_inst(.x({x[430], x[429]}), .y(y[286]));
  Fx287 Fx287_inst(.x({x[431], x[429]}), .y(y[287]));
  Fx288 Fx288_inst(.x({x[433], x[432]}), .y(y[288]));
  Fx289 Fx289_inst(.x({x[434], x[432]}), .y(y[289]));
  Fx290 Fx290_inst(.x({x[436], x[435]}), .y(y[290]));
  Fx291 Fx291_inst(.x({x[437], x[435]}), .y(y[291]));
  Fx292 Fx292_inst(.x({x[439], x[438]}), .y(y[292]));
  Fx293 Fx293_inst(.x({x[440], x[438]}), .y(y[293]));
  Fx294 Fx294_inst(.x({x[442], x[441]}), .y(y[294]));
  Fx295 Fx295_inst(.x({x[443], x[441]}), .y(y[295]));
  Fx296 Fx296_inst(.x({x[445], x[444]}), .y(y[296]));
  Fx297 Fx297_inst(.x({x[446], x[444]}), .y(y[297]));
  Fx298 Fx298_inst(.x({x[448], x[447]}), .y(y[298]));
  Fx299 Fx299_inst(.x({x[449], x[447]}), .y(y[299]));
  Fx300 Fx300_inst(.x({x[451], x[450]}), .y(y[300]));
  Fx301 Fx301_inst(.x({x[452], x[450]}), .y(y[301]));
  Fx302 Fx302_inst(.x({x[454], x[453]}), .y(y[302]));
  Fx303 Fx303_inst(.x({x[455], x[453]}), .y(y[303]));
  Fx304 Fx304_inst(.x({x[457], x[456]}), .y(y[304]));
  Fx305 Fx305_inst(.x({x[458], x[456]}), .y(y[305]));
  Fx306 Fx306_inst(.x({x[460], x[459]}), .y(y[306]));
  Fx307 Fx307_inst(.x({x[461], x[459]}), .y(y[307]));
  Fx308 Fx308_inst(.x({x[463], x[462]}), .y(y[308]));
  Fx309 Fx309_inst(.x({x[464], x[462]}), .y(y[309]));
  Fx310 Fx310_inst(.x({x[466], x[465]}), .y(y[310]));
  Fx311 Fx311_inst(.x({x[467], x[465]}), .y(y[311]));
  Fx312 Fx312_inst(.x({x[469], x[468]}), .y(y[312]));
  Fx313 Fx313_inst(.x({x[470], x[468]}), .y(y[313]));
  Fx314 Fx314_inst(.x({x[472], x[471]}), .y(y[314]));
  Fx315 Fx315_inst(.x({x[473], x[471]}), .y(y[315]));
  Fx316 Fx316_inst(.x({x[475], x[474]}), .y(y[316]));
  Fx317 Fx317_inst(.x({x[476], x[474]}), .y(y[317]));
  Fx318 Fx318_inst(.x({x[478], x[477]}), .y(y[318]));
  Fx319 Fx319_inst(.x({x[479], x[477]}), .y(y[319]));
  Fx320 Fx320_inst(.x({x[481], x[480]}), .y(y[320]));
  Fx321 Fx321_inst(.x({x[482], x[480]}), .y(y[321]));
  Fx322 Fx322_inst(.x({x[484], x[483]}), .y(y[322]));
  Fx323 Fx323_inst(.x({x[485], x[483]}), .y(y[323]));
  Fx324 Fx324_inst(.x({x[487], x[486]}), .y(y[324]));
  Fx325 Fx325_inst(.x({x[488], x[486]}), .y(y[325]));
  Fx326 Fx326_inst(.x({x[490], x[489]}), .y(y[326]));
  Fx327 Fx327_inst(.x({x[491], x[489]}), .y(y[327]));
  Fx328 Fx328_inst(.x({x[493], x[492]}), .y(y[328]));
  Fx329 Fx329_inst(.x({x[494], x[492]}), .y(y[329]));
  Fx330 Fx330_inst(.x({x[496], x[495]}), .y(y[330]));
  Fx331 Fx331_inst(.x({x[497], x[495]}), .y(y[331]));
  Fx332 Fx332_inst(.x({x[499], x[498]}), .y(y[332]));
  Fx333 Fx333_inst(.x({x[500], x[498]}), .y(y[333]));
  Fx334 Fx334_inst(.x({x[502], x[501]}), .y(y[334]));
  Fx335 Fx335_inst(.x({x[503], x[501]}), .y(y[335]));
  Fx336 Fx336_inst(.x({x[505], x[504]}), .y(y[336]));
  Fx337 Fx337_inst(.x({x[506], x[504]}), .y(y[337]));
  Fx338 Fx338_inst(.x({x[508], x[507]}), .y(y[338]));
  Fx339 Fx339_inst(.x({x[509], x[507]}), .y(y[339]));
  Fx340 Fx340_inst(.x({x[511], x[510]}), .y(y[340]));
  Fx341 Fx341_inst(.x({x[512], x[510]}), .y(y[341]));
  Fx342 Fx342_inst(.x({x[514], x[513]}), .y(y[342]));
  Fx343 Fx343_inst(.x({x[515], x[513]}), .y(y[343]));
  Fx344 Fx344_inst(.x({x[517], x[516]}), .y(y[344]));
  Fx345 Fx345_inst(.x({x[518], x[516]}), .y(y[345]));
  Fx346 Fx346_inst(.x({x[520], x[519]}), .y(y[346]));
  Fx347 Fx347_inst(.x({x[521], x[519]}), .y(y[347]));
  Fx348 Fx348_inst(.x({x[523], x[522]}), .y(y[348]));
  Fx349 Fx349_inst(.x({x[524], x[522]}), .y(y[349]));
  Fx350 Fx350_inst(.x({x[526], x[525]}), .y(y[350]));
  Fx351 Fx351_inst(.x({x[527], x[525]}), .y(y[351]));
  Fx352 Fx352_inst(.x({x[529], x[528]}), .y(y[352]));
  Fx353 Fx353_inst(.x({x[530], x[528]}), .y(y[353]));
  Fx354 Fx354_inst(.x({x[532], x[531]}), .y(y[354]));
  Fx355 Fx355_inst(.x({x[533], x[531]}), .y(y[355]));
  Fx356 Fx356_inst(.x({x[535], x[534]}), .y(y[356]));
  Fx357 Fx357_inst(.x({x[536], x[534]}), .y(y[357]));
  Fx358 Fx358_inst(.x({x[538], x[537]}), .y(y[358]));
  Fx359 Fx359_inst(.x({x[539], x[537]}), .y(y[359]));
  Fx360 Fx360_inst(.x({x[541], x[540]}), .y(y[360]));
  Fx361 Fx361_inst(.x({x[542], x[540]}), .y(y[361]));
  Fx362 Fx362_inst(.x({x[544], x[543]}), .y(y[362]));
  Fx363 Fx363_inst(.x({x[545], x[543]}), .y(y[363]));
  Fx364 Fx364_inst(.x({x[547], x[546]}), .y(y[364]));
  Fx365 Fx365_inst(.x({x[548], x[546]}), .y(y[365]));
  Fx366 Fx366_inst(.x({x[550], x[549]}), .y(y[366]));
  Fx367 Fx367_inst(.x({x[551], x[549]}), .y(y[367]));
  Fx368 Fx368_inst(.x({x[553], x[552]}), .y(y[368]));
  Fx369 Fx369_inst(.x({x[554], x[552]}), .y(y[369]));
  Fx370 Fx370_inst(.x({x[556], x[555]}), .y(y[370]));
  Fx371 Fx371_inst(.x({x[557], x[555]}), .y(y[371]));
  Fx372 Fx372_inst(.x({x[559], x[558]}), .y(y[372]));
  Fx373 Fx373_inst(.x({x[560], x[558]}), .y(y[373]));
  Fx374 Fx374_inst(.x({x[562], x[561]}), .y(y[374]));
  Fx375 Fx375_inst(.x({x[563], x[561]}), .y(y[375]));
  Fx376 Fx376_inst(.x({x[565], x[564]}), .y(y[376]));
  Fx377 Fx377_inst(.x({x[566], x[564]}), .y(y[377]));
  Fx378 Fx378_inst(.x({x[568], x[567]}), .y(y[378]));
  Fx379 Fx379_inst(.x({x[569], x[567]}), .y(y[379]));
  Fx380 Fx380_inst(.x({x[571], x[570]}), .y(y[380]));
  Fx381 Fx381_inst(.x({x[572], x[570]}), .y(y[381]));
  Fx382 Fx382_inst(.x({x[574], x[573]}), .y(y[382]));
  Fx383 Fx383_inst(.x({x[575], x[573]}), .y(y[383]));
  Fx384 Fx384_inst(.x({x[577], x[576]}), .y(y[384]));
  Fx385 Fx385_inst(.x({x[578], x[576]}), .y(y[385]));
  Fx386 Fx386_inst(.x({x[580], x[579]}), .y(y[386]));
  Fx387 Fx387_inst(.x({x[581], x[579]}), .y(y[387]));
  Fx388 Fx388_inst(.x({x[583], x[582]}), .y(y[388]));
  Fx389 Fx389_inst(.x({x[584], x[582]}), .y(y[389]));
  Fx390 Fx390_inst(.x({x[586], x[585]}), .y(y[390]));
  Fx391 Fx391_inst(.x({x[587], x[585]}), .y(y[391]));
  Fx392 Fx392_inst(.x({x[589], x[588]}), .y(y[392]));
  Fx393 Fx393_inst(.x({x[590], x[588]}), .y(y[393]));
  Fx394 Fx394_inst(.x({x[592], x[591]}), .y(y[394]));
  Fx395 Fx395_inst(.x({x[593], x[591]}), .y(y[395]));
  Fx396 Fx396_inst(.x({x[595], x[594]}), .y(y[396]));
  Fx397 Fx397_inst(.x({x[596], x[594]}), .y(y[397]));
  Fx398 Fx398_inst(.x({x[598], x[597]}), .y(y[398]));
  Fx399 Fx399_inst(.x({x[599], x[597]}), .y(y[399]));
  Fx400 Fx400_inst(.x({x[601], x[600]}), .y(y[400]));
  Fx401 Fx401_inst(.x({x[602], x[600]}), .y(y[401]));
  Fx402 Fx402_inst(.x({x[604], x[603]}), .y(y[402]));
  Fx403 Fx403_inst(.x({x[605], x[603]}), .y(y[403]));
  Fx404 Fx404_inst(.x({x[607], x[606]}), .y(y[404]));
  Fx405 Fx405_inst(.x({x[608], x[606]}), .y(y[405]));
  Fx406 Fx406_inst(.x({x[610], x[609]}), .y(y[406]));
  Fx407 Fx407_inst(.x({x[611], x[609]}), .y(y[407]));
  Fx408 Fx408_inst(.x({x[613], x[612]}), .y(y[408]));
  Fx409 Fx409_inst(.x({x[614], x[612]}), .y(y[409]));
  Fx410 Fx410_inst(.x({x[616], x[615]}), .y(y[410]));
  Fx411 Fx411_inst(.x({x[617], x[615]}), .y(y[411]));
  Fx412 Fx412_inst(.x({x[619], x[618]}), .y(y[412]));
  Fx413 Fx413_inst(.x({x[620], x[618]}), .y(y[413]));
  Fx414 Fx414_inst(.x({x[622], x[621]}), .y(y[414]));
  Fx415 Fx415_inst(.x({x[623], x[621]}), .y(y[415]));
  Fx416 Fx416_inst(.x({x[625], x[624]}), .y(y[416]));
  Fx417 Fx417_inst(.x({x[626], x[624]}), .y(y[417]));
  Fx418 Fx418_inst(.x({x[628], x[627]}), .y(y[418]));
  Fx419 Fx419_inst(.x({x[629], x[627]}), .y(y[419]));
  Fx420 Fx420_inst(.x({x[631], x[630]}), .y(y[420]));
  Fx421 Fx421_inst(.x({x[632], x[630]}), .y(y[421]));
  Fx422 Fx422_inst(.x({x[634], x[633]}), .y(y[422]));
  Fx423 Fx423_inst(.x({x[635], x[633]}), .y(y[423]));
  Fx424 Fx424_inst(.x({x[637], x[636]}), .y(y[424]));
  Fx425 Fx425_inst(.x({x[638], x[636]}), .y(y[425]));
  Fx426 Fx426_inst(.x({x[640], x[639]}), .y(y[426]));
  Fx427 Fx427_inst(.x({x[641], x[639]}), .y(y[427]));
  Fx428 Fx428_inst(.x({x[643], x[642]}), .y(y[428]));
  Fx429 Fx429_inst(.x({x[644], x[642]}), .y(y[429]));
  Fx430 Fx430_inst(.x({x[646], x[645]}), .y(y[430]));
  Fx431 Fx431_inst(.x({x[647], x[645]}), .y(y[431]));
  Fx432 Fx432_inst(.x({x[649], x[648]}), .y(y[432]));
  Fx433 Fx433_inst(.x({x[650], x[648]}), .y(y[433]));
  Fx434 Fx434_inst(.x({x[652], x[651]}), .y(y[434]));
  Fx435 Fx435_inst(.x({x[653], x[651]}), .y(y[435]));
  Fx436 Fx436_inst(.x({x[655], x[654]}), .y(y[436]));
  Fx437 Fx437_inst(.x({x[656], x[654]}), .y(y[437]));
  Fx438 Fx438_inst(.x({x[658], x[657]}), .y(y[438]));
  Fx439 Fx439_inst(.x({x[659], x[657]}), .y(y[439]));
  Fx440 Fx440_inst(.x({x[661], x[660]}), .y(y[440]));
  Fx441 Fx441_inst(.x({x[662], x[660]}), .y(y[441]));
  Fx442 Fx442_inst(.x({x[664], x[663]}), .y(y[442]));
  Fx443 Fx443_inst(.x({x[665], x[663]}), .y(y[443]));
  Fx444 Fx444_inst(.x({x[667], x[666]}), .y(y[444]));
  Fx445 Fx445_inst(.x({x[668], x[666]}), .y(y[445]));
  Fx446 Fx446_inst(.x({x[670], x[669]}), .y(y[446]));
  Fx447 Fx447_inst(.x({x[671], x[669]}), .y(y[447]));
  Fx448 Fx448_inst(.x({x[673], x[672]}), .y(y[448]));
  Fx449 Fx449_inst(.x({x[674], x[672]}), .y(y[449]));
  Fx450 Fx450_inst(.x({x[676], x[675]}), .y(y[450]));
  Fx451 Fx451_inst(.x({x[677], x[675]}), .y(y[451]));
  Fx452 Fx452_inst(.x({x[679], x[678]}), .y(y[452]));
  Fx453 Fx453_inst(.x({x[680], x[678]}), .y(y[453]));
  Fx454 Fx454_inst(.x({x[682], x[681]}), .y(y[454]));
  Fx455 Fx455_inst(.x({x[683], x[681]}), .y(y[455]));
  Fx456 Fx456_inst(.x({x[685], x[684]}), .y(y[456]));
  Fx457 Fx457_inst(.x({x[686], x[684]}), .y(y[457]));
  Fx458 Fx458_inst(.x({x[688], x[687]}), .y(y[458]));
  Fx459 Fx459_inst(.x({x[689], x[687]}), .y(y[459]));
  Fx460 Fx460_inst(.x({x[691], x[690]}), .y(y[460]));
  Fx461 Fx461_inst(.x({x[692], x[690]}), .y(y[461]));
  Fx462 Fx462_inst(.x({x[694], x[693]}), .y(y[462]));
  Fx463 Fx463_inst(.x({x[695], x[693]}), .y(y[463]));
  Fx464 Fx464_inst(.x({x[697], x[696]}), .y(y[464]));
  Fx465 Fx465_inst(.x({x[698], x[696]}), .y(y[465]));
  Fx466 Fx466_inst(.x({x[700], x[699]}), .y(y[466]));
  Fx467 Fx467_inst(.x({x[701], x[699]}), .y(y[467]));
  Fx468 Fx468_inst(.x({x[703], x[702]}), .y(y[468]));
  Fx469 Fx469_inst(.x({x[704], x[702]}), .y(y[469]));
  Fx470 Fx470_inst(.x({x[706], x[705]}), .y(y[470]));
  Fx471 Fx471_inst(.x({x[707], x[705]}), .y(y[471]));
  Fx472 Fx472_inst(.x({x[709], x[708]}), .y(y[472]));
  Fx473 Fx473_inst(.x({x[710], x[708]}), .y(y[473]));
  Fx474 Fx474_inst(.x({x[712], x[711]}), .y(y[474]));
  Fx475 Fx475_inst(.x({x[713], x[711]}), .y(y[475]));
  Fx476 Fx476_inst(.x({x[715], x[714]}), .y(y[476]));
  Fx477 Fx477_inst(.x({x[716], x[714]}), .y(y[477]));
  Fx478 Fx478_inst(.x({x[718], x[717]}), .y(y[478]));
  Fx479 Fx479_inst(.x({x[719], x[717]}), .y(y[479]));
  Fx480 Fx480_inst(.x({x[721], x[720]}), .y(y[480]));
  Fx481 Fx481_inst(.x({x[722], x[720]}), .y(y[481]));
  Fx482 Fx482_inst(.x({x[724], x[723]}), .y(y[482]));
  Fx483 Fx483_inst(.x({x[725], x[723]}), .y(y[483]));
  Fx484 Fx484_inst(.x({x[727], x[726]}), .y(y[484]));
  Fx485 Fx485_inst(.x({x[728], x[726]}), .y(y[485]));
  Fx486 Fx486_inst(.x({x[730], x[729]}), .y(y[486]));
  Fx487 Fx487_inst(.x({x[731], x[729]}), .y(y[487]));
  Fx488 Fx488_inst(.x({x[733], x[732]}), .y(y[488]));
  Fx489 Fx489_inst(.x({x[734], x[732]}), .y(y[489]));
  Fx490 Fx490_inst(.x({x[736], x[735]}), .y(y[490]));
  Fx491 Fx491_inst(.x({x[737], x[735]}), .y(y[491]));
  Fx492 Fx492_inst(.x({x[739], x[738]}), .y(y[492]));
  Fx493 Fx493_inst(.x({x[740], x[738]}), .y(y[493]));
  Fx494 Fx494_inst(.x({x[742], x[741]}), .y(y[494]));
  Fx495 Fx495_inst(.x({x[743], x[741]}), .y(y[495]));
  Fx496 Fx496_inst(.x({x[745], x[744]}), .y(y[496]));
  Fx497 Fx497_inst(.x({x[746], x[744]}), .y(y[497]));
  Fx498 Fx498_inst(.x({x[748], x[747]}), .y(y[498]));
  Fx499 Fx499_inst(.x({x[749], x[747]}), .y(y[499]));
  Fx500 Fx500_inst(.x({x[751], x[750]}), .y(y[500]));
  Fx501 Fx501_inst(.x({x[752], x[750]}), .y(y[501]));
  Fx502 Fx502_inst(.x({x[754], x[753]}), .y(y[502]));
  Fx503 Fx503_inst(.x({x[755], x[753]}), .y(y[503]));
  Fx504 Fx504_inst(.x({x[757], x[756]}), .y(y[504]));
  Fx505 Fx505_inst(.x({x[758], x[756]}), .y(y[505]));
  Fx506 Fx506_inst(.x({x[760], x[759]}), .y(y[506]));
  Fx507 Fx507_inst(.x({x[761], x[759]}), .y(y[507]));
  Fx508 Fx508_inst(.x({x[763], x[762]}), .y(y[508]));
  Fx509 Fx509_inst(.x({x[764], x[762]}), .y(y[509]));
  Fx510 Fx510_inst(.x({x[766], x[765]}), .y(y[510]));
  Fx511 Fx511_inst(.x({x[767], x[765]}), .y(y[511]));
  Fx512 Fx512_inst(.x({x[769], x[768]}), .y(y[512]));
  Fx513 Fx513_inst(.x({x[770], x[768]}), .y(y[513]));
  Fx514 Fx514_inst(.x({x[772], x[771]}), .y(y[514]));
  Fx515 Fx515_inst(.x({x[773], x[771]}), .y(y[515]));
  Fx516 Fx516_inst(.x({x[775], x[774]}), .y(y[516]));
  Fx517 Fx517_inst(.x({x[776], x[774]}), .y(y[517]));
  Fx518 Fx518_inst(.x({x[778], x[777]}), .y(y[518]));
  Fx519 Fx519_inst(.x({x[779], x[777]}), .y(y[519]));
  Fx520 Fx520_inst(.x({x[781], x[780]}), .y(y[520]));
  Fx521 Fx521_inst(.x({x[782], x[780]}), .y(y[521]));
  Fx522 Fx522_inst(.x({x[784], x[783]}), .y(y[522]));
  Fx523 Fx523_inst(.x({x[785], x[783]}), .y(y[523]));
  Fx524 Fx524_inst(.x({x[787], x[786]}), .y(y[524]));
  Fx525 Fx525_inst(.x({x[788], x[786]}), .y(y[525]));
  Fx526 Fx526_inst(.x({x[790], x[789]}), .y(y[526]));
  Fx527 Fx527_inst(.x({x[791], x[789]}), .y(y[527]));
  Fx528 Fx528_inst(.x({x[793], x[792]}), .y(y[528]));
  Fx529 Fx529_inst(.x({x[794], x[792]}), .y(y[529]));
  Fx530 Fx530_inst(.x({x[796], x[795]}), .y(y[530]));
  Fx531 Fx531_inst(.x({x[797], x[795]}), .y(y[531]));
  Fx532 Fx532_inst(.x({x[799], x[798]}), .y(y[532]));
  Fx533 Fx533_inst(.x({x[800], x[798]}), .y(y[533]));
  Fx534 Fx534_inst(.x({x[802], x[801]}), .y(y[534]));
  Fx535 Fx535_inst(.x({x[803], x[801]}), .y(y[535]));
  Fx536 Fx536_inst(.x({x[805], x[804]}), .y(y[536]));
  Fx537 Fx537_inst(.x({x[806], x[804]}), .y(y[537]));
  Fx538 Fx538_inst(.x({x[808], x[807]}), .y(y[538]));
  Fx539 Fx539_inst(.x({x[809], x[807]}), .y(y[539]));
  Fx540 Fx540_inst(.x({x[811], x[810]}), .y(y[540]));
  Fx541 Fx541_inst(.x({x[812], x[810]}), .y(y[541]));
  Fx542 Fx542_inst(.x({x[814], x[813]}), .y(y[542]));
  Fx543 Fx543_inst(.x({x[815], x[813]}), .y(y[543]));
  Fx544 Fx544_inst(.x({x[817], x[816]}), .y(y[544]));
  Fx545 Fx545_inst(.x({x[818], x[816]}), .y(y[545]));
  Fx546 Fx546_inst(.x({x[820], x[819]}), .y(y[546]));
  Fx547 Fx547_inst(.x({x[821], x[819]}), .y(y[547]));
  Fx548 Fx548_inst(.x({x[823], x[822]}), .y(y[548]));
  Fx549 Fx549_inst(.x({x[824], x[822]}), .y(y[549]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind66(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind67(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind68(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind69(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind70(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind71(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind72(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind73(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind74(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind75(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind76(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind77(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind78(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind79(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind80(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind81(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind82(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind83(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind84(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind85(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind86(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind87(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind88(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind89(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind90(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind91(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind92(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind93(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind94(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind95(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind96(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind97(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind98(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind99(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind100(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind101(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind102(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind103(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind104(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind105(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind106(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind107(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind108(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind109(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind110(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind111(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind112(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind113(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind114(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind115(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind116(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind117(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind118(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind119(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind120(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind121(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind122(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind123(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind124(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind125(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind126(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind127(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind128(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind129(x, y);
 input [35:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[20] | t[21]);
  assign t[11] = ~(t[22] | t[23]);
  assign t[12] = t[24] ^ x[2];
  assign t[13] = t[25] ^ x[5];
  assign t[14] = t[26] ^ x[8];
  assign t[15] = t[27] ^ x[11];
  assign t[16] = t[28] ^ x[14];
  assign t[17] = t[29] ^ x[17];
  assign t[18] = t[30] ^ x[20];
  assign t[19] = t[31] ^ x[23];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[32] ^ x[26];
  assign t[21] = t[33] ^ x[29];
  assign t[22] = t[34] ^ x[32];
  assign t[23] = t[35] ^ x[35];
  assign t[24] = (x[0] & x[1]);
  assign t[25] = (x[3] & x[4]);
  assign t[26] = (x[6] & x[7]);
  assign t[27] = (x[9] & x[10]);
  assign t[28] = (x[12] & x[13]);
  assign t[29] = (x[15] & x[16]);
  assign t[2] = ~(t[5] | t[6]);
  assign t[30] = (x[18] & x[19]);
  assign t[31] = (x[21] & x[22]);
  assign t[32] = (x[24] & x[25]);
  assign t[33] = (x[27] & x[28]);
  assign t[34] = (x[30] & x[31]);
  assign t[35] = (x[33] & x[34]);
  assign t[3] = ~(t[13] & t[14]);
  assign t[4] = ~(t[15] & t[16]);
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[17] & t[8]);
  assign t[7] = ~(t[18] | t[9]);
  assign t[8] = ~(t[19]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = t[12] & t[0];
endmodule

module R1ind130(x, y);
 input x;
 output y;

  assign y = ~(x);
endmodule

module R1ind131(x, y);
 input [41:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[10] = ~(t[24] | t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[25] & t[26]);
  assign t[15] = ~(t[27] & t[28]);
  assign t[16] = ~(t[10]);
  assign t[17] = ~(t[29] & t[20]);
  assign t[18] = ~(t[30] | t[31]);
  assign t[19] = ~(t[32] | t[33]);
  assign t[1] = ~(t[4]);
  assign t[20] = ~(t[34]);
  assign t[21] = t[35] ^ x[2];
  assign t[22] = t[36] ^ x[5];
  assign t[23] = t[37] ^ x[8];
  assign t[24] = t[38] ^ x[11];
  assign t[25] = t[39] ^ x[14];
  assign t[26] = t[40] ^ x[17];
  assign t[27] = t[41] ^ x[20];
  assign t[28] = t[42] ^ x[23];
  assign t[29] = t[43] ^ x[26];
  assign t[2] = ~(t[22]);
  assign t[30] = t[44] ^ x[29];
  assign t[31] = t[45] ^ x[32];
  assign t[32] = t[46] ^ x[35];
  assign t[33] = t[47] ^ x[38];
  assign t[34] = t[48] ^ x[41];
  assign t[35] = (x[0] & x[1]);
  assign t[36] = (x[3] & x[4]);
  assign t[37] = (x[6] & x[7]);
  assign t[38] = (x[9] & x[10]);
  assign t[39] = (x[12] & x[13]);
  assign t[3] = ~(t[23]);
  assign t[40] = (x[15] & x[16]);
  assign t[41] = (x[18] & x[19]);
  assign t[42] = (x[21] & x[22]);
  assign t[43] = (x[24] & x[25]);
  assign t[44] = (x[27] & x[28]);
  assign t[45] = (x[30] & x[31]);
  assign t[46] = (x[33] & x[34]);
  assign t[47] = (x[36] & x[37]);
  assign t[48] = (x[39] & x[40]);
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[8]);
  assign t[7] = t[21] & t[9];
  assign t[8] = ~(t[21] & t[10]);
  assign t[9] = t[11] & t[12];
  assign y = ~(t[21] & t[0]);
endmodule

module R1ind132(x, y);
 input [38:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = ~(t[23] & t[2]);
  assign t[10] = ~(t[25] & t[12]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] | t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[27] & t[24]);
  assign t[17] = ~(t[28] & t[29]);
  assign t[18] = ~(t[12]);
  assign t[19] = ~(t[30] & t[22]);
  assign t[1] = ~(t[24] & t[3]);
  assign t[20] = ~(t[31] | t[32]);
  assign t[21] = ~(t[33] | t[34]);
  assign t[22] = ~(t[35]);
  assign t[23] = t[36] ^ x[2];
  assign t[24] = t[37] ^ x[5];
  assign t[25] = t[38] ^ x[8];
  assign t[26] = t[39] ^ x[11];
  assign t[27] = t[40] ^ x[14];
  assign t[28] = t[41] ^ x[17];
  assign t[29] = t[42] ^ x[20];
  assign t[2] = ~(t[4] | t[5]);
  assign t[30] = t[43] ^ x[23];
  assign t[31] = t[44] ^ x[26];
  assign t[32] = t[45] ^ x[29];
  assign t[33] = t[46] ^ x[32];
  assign t[34] = t[47] ^ x[35];
  assign t[35] = t[48] ^ x[38];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[6] & x[7]);
  assign t[39] = (x[9] & x[10]);
  assign t[3] = ~(t[6] | t[5]);
  assign t[40] = (x[12] & x[13]);
  assign t[41] = (x[15] & x[16]);
  assign t[42] = (x[18] & x[19]);
  assign t[43] = (x[21] & x[22]);
  assign t[44] = (x[24] & x[25]);
  assign t[45] = (x[27] & x[28]);
  assign t[46] = (x[30] & x[31]);
  assign t[47] = (x[33] & x[34]);
  assign t[48] = (x[36] & x[37]);
  assign t[4] = t[7] & t[8];
  assign t[5] = ~(t[25]);
  assign t[6] = ~(t[4]);
  assign t[7] = ~(t[9]);
  assign t[8] = ~(t[10]);
  assign t[9] = t[25] & t[11];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind133(x, y);
 input [35:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[23] & t[2]);
  assign t[10] = ~(t[25] & t[12]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] | t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] & t[21]);
  assign t[16] = ~(t[27] & t[23]);
  assign t[17] = ~(t[24] & t[28]);
  assign t[18] = ~(t[12]);
  assign t[19] = ~(t[29] & t[22]);
  assign t[1] = ~(t[24] & t[3]);
  assign t[20] = ~(t[30] | t[31]);
  assign t[21] = ~(t[32] | t[33]);
  assign t[22] = ~(t[34]);
  assign t[23] = t[35] ^ x[2];
  assign t[24] = t[36] ^ x[5];
  assign t[25] = t[37] ^ x[8];
  assign t[26] = t[38] ^ x[11];
  assign t[27] = t[39] ^ x[14];
  assign t[28] = t[40] ^ x[17];
  assign t[29] = t[41] ^ x[20];
  assign t[2] = ~(t[4] | t[5]);
  assign t[30] = t[42] ^ x[23];
  assign t[31] = t[43] ^ x[26];
  assign t[32] = t[44] ^ x[29];
  assign t[33] = t[45] ^ x[32];
  assign t[34] = t[46] ^ x[35];
  assign t[35] = (x[0] & x[1]);
  assign t[36] = (x[3] & x[4]);
  assign t[37] = (x[6] & x[7]);
  assign t[38] = (x[9] & x[10]);
  assign t[39] = (x[12] & x[13]);
  assign t[3] = ~(t[6] | t[5]);
  assign t[40] = (x[15] & x[16]);
  assign t[41] = (x[18] & x[19]);
  assign t[42] = (x[21] & x[22]);
  assign t[43] = (x[24] & x[25]);
  assign t[44] = (x[27] & x[28]);
  assign t[45] = (x[30] & x[31]);
  assign t[46] = (x[33] & x[34]);
  assign t[4] = t[7] & t[8];
  assign t[5] = ~(t[25]);
  assign t[6] = ~(t[4]);
  assign t[7] = ~(t[9]);
  assign t[8] = ~(t[10]);
  assign t[9] = t[25] & t[11];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind134(x, y);
 input [41:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[13]);
  assign t[12] = t[29] & t[14];
  assign t[13] = ~(t[29] & t[15]);
  assign t[14] = t[16] & t[17];
  assign t[15] = ~(t[30] | t[18]);
  assign t[16] = ~(t[19] | t[20]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[31] & t[32]);
  assign t[1] = ~(t[26] & t[4]);
  assign t[20] = ~(t[26] & t[33]);
  assign t[21] = ~(t[15]);
  assign t[22] = ~(t[34] & t[25]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = ~(t[39]);
  assign t[26] = t[40] ^ x[2];
  assign t[27] = t[41] ^ x[5];
  assign t[28] = t[42] ^ x[8];
  assign t[29] = t[43] ^ x[11];
  assign t[2] = t[5] ^ t[6];
  assign t[30] = t[44] ^ x[14];
  assign t[31] = t[45] ^ x[17];
  assign t[32] = t[46] ^ x[20];
  assign t[33] = t[47] ^ x[23];
  assign t[34] = t[48] ^ x[26];
  assign t[35] = t[49] ^ x[29];
  assign t[36] = t[50] ^ x[32];
  assign t[37] = t[51] ^ x[35];
  assign t[38] = t[52] ^ x[38];
  assign t[39] = t[53] ^ x[41];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (x[0] & x[1]);
  assign t[41] = (x[3] & x[4]);
  assign t[42] = (x[6] & x[7]);
  assign t[43] = (x[9] & x[10]);
  assign t[44] = (x[12] & x[13]);
  assign t[45] = (x[15] & x[16]);
  assign t[46] = (x[18] & x[19]);
  assign t[47] = (x[21] & x[22]);
  assign t[48] = (x[24] & x[25]);
  assign t[49] = (x[27] & x[28]);
  assign t[4] = ~(t[9] | t[8]);
  assign t[50] = (x[30] & x[31]);
  assign t[51] = (x[33] & x[34]);
  assign t[52] = (x[36] & x[37]);
  assign t[53] = (x[39] & x[40]);
  assign t[5] = ~(t[27]);
  assign t[6] = ~(t[28]);
  assign t[7] = ~(t[9]);
  assign t[8] = ~(t[29]);
  assign t[9] = t[10] & t[11];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind135(x, y);
 input [41:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[10] = ~(t[25] | t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[26] & t[27]);
  assign t[15] = ~(t[28] & t[23]);
  assign t[16] = ~(t[10]);
  assign t[17] = ~(t[29] & t[20]);
  assign t[18] = ~(t[30] | t[31]);
  assign t[19] = ~(t[32] | t[33]);
  assign t[1] = ~(t[4]);
  assign t[20] = ~(t[34]);
  assign t[21] = t[35] ^ x[2];
  assign t[22] = t[36] ^ x[5];
  assign t[23] = t[37] ^ x[8];
  assign t[24] = t[38] ^ x[11];
  assign t[25] = t[39] ^ x[14];
  assign t[26] = t[40] ^ x[17];
  assign t[27] = t[41] ^ x[20];
  assign t[28] = t[42] ^ x[23];
  assign t[29] = t[43] ^ x[26];
  assign t[2] = ~(t[22] ^ t[23]);
  assign t[30] = t[44] ^ x[29];
  assign t[31] = t[45] ^ x[32];
  assign t[32] = t[46] ^ x[35];
  assign t[33] = t[47] ^ x[38];
  assign t[34] = t[48] ^ x[41];
  assign t[35] = (x[0] & x[1]);
  assign t[36] = (x[3] & x[4]);
  assign t[37] = (x[6] & x[7]);
  assign t[38] = (x[9] & x[10]);
  assign t[39] = (x[12] & x[13]);
  assign t[3] = ~(t[24]);
  assign t[40] = (x[15] & x[16]);
  assign t[41] = (x[18] & x[19]);
  assign t[42] = (x[21] & x[22]);
  assign t[43] = (x[24] & x[25]);
  assign t[44] = (x[27] & x[28]);
  assign t[45] = (x[30] & x[31]);
  assign t[46] = (x[33] & x[34]);
  assign t[47] = (x[36] & x[37]);
  assign t[48] = (x[39] & x[40]);
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[8]);
  assign t[7] = t[21] & t[9];
  assign t[8] = ~(t[21] & t[10]);
  assign t[9] = t[11] & t[12];
  assign y = ~(t[21] & t[0]);
endmodule

module R1ind136(x, y);
 input [35:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[10] = ~(t[24] | t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[22] & t[25]);
  assign t[15] = ~(t[26] & t[23]);
  assign t[16] = ~(t[10]);
  assign t[17] = ~(t[27] & t[20]);
  assign t[18] = ~(t[28] | t[29]);
  assign t[19] = ~(t[30] | t[31]);
  assign t[1] = ~(t[4]);
  assign t[20] = ~(t[32]);
  assign t[21] = t[33] ^ x[2];
  assign t[22] = t[34] ^ x[5];
  assign t[23] = t[35] ^ x[8];
  assign t[24] = t[36] ^ x[11];
  assign t[25] = t[37] ^ x[14];
  assign t[26] = t[38] ^ x[17];
  assign t[27] = t[39] ^ x[20];
  assign t[28] = t[40] ^ x[23];
  assign t[29] = t[41] ^ x[26];
  assign t[2] = ~(t[22]);
  assign t[30] = t[42] ^ x[29];
  assign t[31] = t[43] ^ x[32];
  assign t[32] = t[44] ^ x[35];
  assign t[33] = (x[0] & x[1]);
  assign t[34] = (x[3] & x[4]);
  assign t[35] = (x[6] & x[7]);
  assign t[36] = (x[9] & x[10]);
  assign t[37] = (x[12] & x[13]);
  assign t[38] = (x[15] & x[16]);
  assign t[39] = (x[18] & x[19]);
  assign t[3] = ~(t[23]);
  assign t[40] = (x[21] & x[22]);
  assign t[41] = (x[24] & x[25]);
  assign t[42] = (x[27] & x[28]);
  assign t[43] = (x[30] & x[31]);
  assign t[44] = (x[33] & x[34]);
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[8]);
  assign t[7] = t[21] & t[9];
  assign t[8] = ~(t[21] & t[10]);
  assign t[9] = t[11] & t[12];
  assign y = ~(t[21] & t[0]);
endmodule

module R1ind137(x, y);
 input [41:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[27] & t[12];
  assign t[11] = ~(t[27] & t[13]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] | t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[24] & t[29]);
  assign t[18] = ~(t[30] & t[31]);
  assign t[19] = ~(t[13]);
  assign t[1] = ~(t[4] & t[24]);
  assign t[20] = ~(t[32] & t[23]);
  assign t[21] = ~(t[33] | t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[8];
  assign t[27] = t[41] ^ x[11];
  assign t[28] = t[42] ^ x[14];
  assign t[29] = t[43] ^ x[17];
  assign t[2] = t[25] ^ t[26];
  assign t[30] = t[44] ^ x[20];
  assign t[31] = t[45] ^ x[23];
  assign t[32] = t[46] ^ x[26];
  assign t[33] = t[47] ^ x[29];
  assign t[34] = t[48] ^ x[32];
  assign t[35] = t[49] ^ x[35];
  assign t[36] = t[50] ^ x[38];
  assign t[37] = t[51] ^ x[41];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = (x[6] & x[7]);
  assign t[41] = (x[9] & x[10]);
  assign t[42] = (x[12] & x[13]);
  assign t[43] = (x[15] & x[16]);
  assign t[44] = (x[18] & x[19]);
  assign t[45] = (x[21] & x[22]);
  assign t[46] = (x[24] & x[25]);
  assign t[47] = (x[27] & x[28]);
  assign t[48] = (x[30] & x[31]);
  assign t[49] = (x[33] & x[34]);
  assign t[4] = ~(t[7] | t[6]);
  assign t[50] = (x[36] & x[37]);
  assign t[51] = (x[39] & x[40]);
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[27]);
  assign t[7] = t[8] & t[9];
  assign t[8] = ~(t[10]);
  assign t[9] = ~(t[11]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind138(x, y);
 input [41:0] x;
 output y;

 wire [48:0] t;
  assign t[0] = t[1] ? t[3] : t[2];
  assign t[10] = ~(t[24] | t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(t[18] & t[19]);
  assign t[14] = ~(t[25] & t[26]);
  assign t[15] = ~(t[27] & t[28]);
  assign t[16] = ~(t[10]);
  assign t[17] = ~(t[29] & t[20]);
  assign t[18] = ~(t[30] | t[31]);
  assign t[19] = ~(t[32] | t[33]);
  assign t[1] = ~(t[4]);
  assign t[20] = ~(t[34]);
  assign t[21] = t[35] ^ x[2];
  assign t[22] = t[36] ^ x[5];
  assign t[23] = t[37] ^ x[8];
  assign t[24] = t[38] ^ x[11];
  assign t[25] = t[39] ^ x[14];
  assign t[26] = t[40] ^ x[17];
  assign t[27] = t[41] ^ x[20];
  assign t[28] = t[42] ^ x[23];
  assign t[29] = t[43] ^ x[26];
  assign t[2] = ~(t[22]);
  assign t[30] = t[44] ^ x[29];
  assign t[31] = t[45] ^ x[32];
  assign t[32] = t[46] ^ x[35];
  assign t[33] = t[47] ^ x[38];
  assign t[34] = t[48] ^ x[41];
  assign t[35] = (x[0] & x[1]);
  assign t[36] = (x[3] & x[4]);
  assign t[37] = (x[6] & x[7]);
  assign t[38] = (x[9] & x[10]);
  assign t[39] = (x[12] & x[13]);
  assign t[3] = ~(t[23]);
  assign t[40] = (x[15] & x[16]);
  assign t[41] = (x[18] & x[19]);
  assign t[42] = (x[21] & x[22]);
  assign t[43] = (x[24] & x[25]);
  assign t[44] = (x[27] & x[28]);
  assign t[45] = (x[30] & x[31]);
  assign t[46] = (x[33] & x[34]);
  assign t[47] = (x[36] & x[37]);
  assign t[48] = (x[39] & x[40]);
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[7]);
  assign t[6] = ~(t[8]);
  assign t[7] = t[21] & t[9];
  assign t[8] = ~(t[21] & t[10]);
  assign t[9] = t[11] & t[12];
  assign y = ~(t[21] & t[0]);
endmodule

module R1ind139(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind140(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind141(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind142(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind143(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind144(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind145(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind146(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind147(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind148(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind149(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind150(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind151(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind152(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind153(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind154(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind155(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind156(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind157(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind158(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind159(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind160(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind161(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind162(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind163(x, y);
 input [123:0] x;
 output y;

 wire [216:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[73] & t[115];
  assign t[101] = t[166] ^ t[167];
  assign t[102] = t[168] ^ t[169];
  assign t[103] = t[170] ^ t[171];
  assign t[104] = t[172] ^ t[173];
  assign t[105] = t[82] ^ t[85];
  assign t[106] = t[174] ^ t[175];
  assign t[107] = t[116] ^ t[117];
  assign t[108] = t[87] ^ t[118];
  assign t[109] = t[87] & t[118];
  assign t[10] = ~(t[16]);
  assign t[110] = t[53] & t[58];
  assign t[111] = t[119] ^ t[120];
  assign t[112] = t[121] ^ t[122];
  assign t[113] = t[53] ^ t[123];
  assign t[114] = t[70] ^ t[52];
  assign t[115] = t[124] ^ t[120];
  assign t[116] = t[123] & t[85];
  assign t[117] = t[55] & t[125];
  assign t[118] = t[125] ^ t[86];
  assign t[119] = t[126] ^ t[127];
  assign t[11] = t[138] & t[17];
  assign t[120] = t[128] ^ t[110];
  assign t[121] = t[113] & t[114];
  assign t[122] = t[69] & t[52];
  assign t[123] = t[86] ^ t[129];
  assign t[124] = t[130] ^ t[131];
  assign t[125] = t[53] ^ t[66];
  assign t[126] = t[132] ^ t[117];
  assign t[127] = t[71] & t[133];
  assign t[128] = t[37] & t[59];
  assign t[129] = t[49] ^ t[85];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[134] ^ t[122];
  assign t[131] = t[88] & t[70];
  assign t[132] = t[125] ^ t[72];
  assign t[133] = t[85] ^ t[125];
  assign t[134] = t[69] ^ t[52];
  assign t[135] = t[176] ^ x[2];
  assign t[136] = t[177] ^ x[6];
  assign t[137] = t[178] ^ x[9];
  assign t[138] = t[179] ^ x[12];
  assign t[139] = t[180] ^ x[15];
  assign t[13] = ~(t[138]);
  assign t[140] = t[181] ^ x[18];
  assign t[141] = t[182] ^ x[21];
  assign t[142] = t[183] ^ x[24];
  assign t[143] = t[184] ^ x[27];
  assign t[144] = t[185] ^ x[30];
  assign t[145] = t[186] ^ x[33];
  assign t[146] = t[187] ^ x[36];
  assign t[147] = t[188] ^ x[39];
  assign t[148] = t[189] ^ x[42];
  assign t[149] = t[190] ^ x[45];
  assign t[14] = ~(t[20] | t[21]);
  assign t[150] = t[191] ^ x[48];
  assign t[151] = t[192] ^ x[51];
  assign t[152] = t[193] ^ x[54];
  assign t[153] = t[194] ^ x[57];
  assign t[154] = t[195] ^ x[60];
  assign t[155] = t[196] ^ x[63];
  assign t[156] = t[197] ^ x[66];
  assign t[157] = t[198] ^ x[69];
  assign t[158] = t[199] ^ x[72];
  assign t[159] = t[200] ^ x[75];
  assign t[15] = t[22] ^ t[23];
  assign t[160] = t[201] ^ x[78];
  assign t[161] = t[202] ^ x[81];
  assign t[162] = t[203] ^ x[84];
  assign t[163] = t[204] ^ x[87];
  assign t[164] = t[205] ^ x[90];
  assign t[165] = t[206] ^ x[93];
  assign t[166] = t[207] ^ x[96];
  assign t[167] = t[208] ^ x[99];
  assign t[168] = t[209] ^ x[102];
  assign t[169] = t[210] ^ x[105];
  assign t[16] = ~(t[138] & t[24]);
  assign t[170] = t[211] ^ x[108];
  assign t[171] = t[212] ^ x[111];
  assign t[172] = t[213] ^ x[114];
  assign t[173] = t[214] ^ x[117];
  assign t[174] = t[215] ^ x[120];
  assign t[175] = t[216] ^ x[123];
  assign t[176] = (x[0] & x[1]);
  assign t[177] = (x[4] & x[5]);
  assign t[178] = (x[7] & x[8]);
  assign t[179] = (x[10] & x[11]);
  assign t[17] = t[25] & t[26];
  assign t[180] = (x[13] & x[14]);
  assign t[181] = (x[16] & x[17]);
  assign t[182] = (x[19] & x[20]);
  assign t[183] = (x[22] & x[23]);
  assign t[184] = (x[25] & x[26]);
  assign t[185] = (x[28] & x[29]);
  assign t[186] = (x[31] & x[32]);
  assign t[187] = (x[34] & x[35]);
  assign t[188] = (x[37] & x[38]);
  assign t[189] = (x[40] & x[41]);
  assign t[18] = ~(t[139]);
  assign t[190] = (x[43] & x[44]);
  assign t[191] = (x[46] & x[47]);
  assign t[192] = (x[49] & x[50]);
  assign t[193] = (x[52] & x[53]);
  assign t[194] = (x[55] & x[56]);
  assign t[195] = (x[58] & x[59]);
  assign t[196] = (x[61] & x[62]);
  assign t[197] = (x[64] & x[65]);
  assign t[198] = (x[67] & x[68]);
  assign t[199] = (x[70] & x[71]);
  assign t[19] = ~(t[138]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[73] & x[74]);
  assign t[201] = (x[76] & x[77]);
  assign t[202] = (x[79] & x[80]);
  assign t[203] = (x[82] & x[83]);
  assign t[204] = (x[85] & x[86]);
  assign t[205] = (x[88] & x[89]);
  assign t[206] = (x[91] & x[92]);
  assign t[207] = (x[94] & x[95]);
  assign t[208] = (x[97] & x[98]);
  assign t[209] = (x[100] & x[101]);
  assign t[20] = ~(t[140]);
  assign t[210] = (x[103] & x[104]);
  assign t[211] = (x[106] & x[107]);
  assign t[212] = (x[109] & x[110]);
  assign t[213] = (x[112] & x[113]);
  assign t[214] = (x[115] & x[116]);
  assign t[215] = (x[118] & x[119]);
  assign t[216] = (x[121] & x[122]);
  assign t[21] = ~(t[141]);
  assign t[22] = t[27] ^ t[28];
  assign t[23] = t[29] ^ t[30];
  assign t[24] = ~(t[142] | t[31]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = t[36] & t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[6]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = ~(t[143] & t[144]);
  assign t[33] = ~(t[145] & t[146]);
  assign t[34] = ~(t[24]);
  assign t[35] = ~(t[147] & t[46]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = t[49] ^ t[50];
  assign t[38] = t[51] & t[52];
  assign t[39] = t[47] & t[53];
  assign t[3] = ~(t[7]);
  assign t[40] = t[54] & t[55];
  assign t[41] = t[56] ^ t[57];
  assign t[42] = t[47] & t[58];
  assign t[43] = t[36] & t[59];
  assign t[44] = ~(t[148] | t[149]);
  assign t[45] = ~(t[150] | t[151]);
  assign t[46] = ~(t[152]);
  assign t[47] = t[60] ^ t[61];
  assign t[48] = t[62] ^ t[63];
  assign t[49] = t[12] ? t[153] : t[64];
  assign t[4] = t[8] ? t[136] : x[3];
  assign t[50] = t[12] ? t[154] : t[65];
  assign t[51] = t[60] ^ t[62];
  assign t[52] = t[66] ^ t[67];
  assign t[53] = t[68] ^ t[49];
  assign t[54] = t[61] ^ t[63];
  assign t[55] = t[69] ^ t[37];
  assign t[56] = t[62] & t[70];
  assign t[57] = t[63] & t[71];
  assign t[58] = t[66] ^ t[72];
  assign t[59] = t[53] ^ t[67];
  assign t[5] = ~(t[9] ^ t[137]);
  assign t[60] = t[73] ^ t[74];
  assign t[61] = t[75] ^ t[76];
  assign t[62] = t[77] ^ t[78];
  assign t[63] = t[79] ^ t[80];
  assign t[64] = t[155] ^ t[156];
  assign t[65] = t[157] ^ t[158];
  assign t[66] = t[81] ^ t[82];
  assign t[67] = t[83] ^ t[50];
  assign t[68] = t[12] ? t[159] : t[84];
  assign t[69] = t[68] ^ t[82];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[85] ^ t[86];
  assign t[71] = t[87] ^ t[88];
  assign t[72] = t[89] ^ t[50];
  assign t[73] = t[90] ^ t[91];
  assign t[74] = t[92] & t[93];
  assign t[75] = t[94] ^ t[95];
  assign t[76] = t[96] & t[97];
  assign t[77] = t[93] & t[98];
  assign t[78] = t[93] ^ t[99];
  assign t[79] = t[97] & t[100];
  assign t[7] = ~(t[12]);
  assign t[80] = t[97] ^ t[99];
  assign t[81] = t[12] ? t[160] : t[101];
  assign t[82] = t[12] ? t[161] : t[102];
  assign t[83] = t[12] ? t[162] : t[103];
  assign t[84] = t[163] ^ t[137];
  assign t[85] = t[12] ? t[164] : t[104];
  assign t[86] = t[89] ^ t[83];
  assign t[87] = t[68] ^ t[50];
  assign t[88] = t[86] ^ t[105];
  assign t[89] = t[12] ? t[165] : t[106];
  assign t[8] = ~(t[13]);
  assign t[90] = t[107] ^ t[108];
  assign t[91] = t[109] ^ t[110];
  assign t[92] = t[75] ^ t[99];
  assign t[93] = t[111] ^ t[73];
  assign t[94] = t[112] ^ t[91];
  assign t[95] = t[113] ^ t[114];
  assign t[96] = t[73] ^ t[99];
  assign t[97] = t[115] ^ t[75];
  assign t[98] = t[111] & t[75];
  assign t[99] = t[115] & t[111];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = t[0] ? t[1] : t[135];
endmodule

module R1ind164(x, y);
 input [123:0] x;
 output y;

 wire [215:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[166] ^ t[136];
  assign t[101] = t[167] ^ t[168];
  assign t[102] = t[169] ^ t[170];
  assign t[103] = t[171] ^ t[172];
  assign t[104] = t[78] ^ t[63];
  assign t[105] = t[80] ^ t[79];
  assign t[106] = t[79] ^ t[63];
  assign t[107] = t[105] & t[122];
  assign t[108] = t[105] ^ t[63];
  assign t[109] = t[173] ^ t[174];
  assign t[10] = ~(t[16]);
  assign t[110] = t[123] ^ t[124];
  assign t[111] = t[50] & t[125];
  assign t[112] = t[54] & t[60];
  assign t[113] = t[52] & t[59];
  assign t[114] = t[126] ^ t[124];
  assign t[115] = t[52] ^ t[127];
  assign t[116] = t[125] ^ t[128];
  assign t[117] = t[129] ^ t[130];
  assign t[118] = t[49] ^ t[131];
  assign t[119] = t[49] & t[131];
  assign t[11] = t[137] & t[17];
  assign t[120] = t[132] ^ t[130];
  assign t[121] = t[37] & t[73];
  assign t[122] = t[80] & t[78];
  assign t[123] = t[92] ^ t[128];
  assign t[124] = t[92] & t[128];
  assign t[125] = t[86] ^ t[66];
  assign t[126] = t[115] & t[116];
  assign t[127] = t[66] ^ t[133];
  assign t[128] = t[72] ^ t[76];
  assign t[129] = t[127] & t[86];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[74] & t[56];
  assign t[131] = t[56] ^ t[66];
  assign t[132] = t[56] ^ t[75];
  assign t[133] = t[70] ^ t[86];
  assign t[134] = t[175] ^ x[2];
  assign t[135] = t[176] ^ x[6];
  assign t[136] = t[177] ^ x[9];
  assign t[137] = t[178] ^ x[12];
  assign t[138] = t[179] ^ x[15];
  assign t[139] = t[180] ^ x[18];
  assign t[13] = ~(t[137]);
  assign t[140] = t[181] ^ x[21];
  assign t[141] = t[182] ^ x[24];
  assign t[142] = t[183] ^ x[27];
  assign t[143] = t[184] ^ x[30];
  assign t[144] = t[185] ^ x[33];
  assign t[145] = t[186] ^ x[36];
  assign t[146] = t[187] ^ x[39];
  assign t[147] = t[188] ^ x[42];
  assign t[148] = t[189] ^ x[45];
  assign t[149] = t[190] ^ x[48];
  assign t[14] = ~(t[20] | t[21]);
  assign t[150] = t[191] ^ x[51];
  assign t[151] = t[192] ^ x[54];
  assign t[152] = t[193] ^ x[57];
  assign t[153] = t[194] ^ x[60];
  assign t[154] = t[195] ^ x[63];
  assign t[155] = t[196] ^ x[66];
  assign t[156] = t[197] ^ x[69];
  assign t[157] = t[198] ^ x[72];
  assign t[158] = t[199] ^ x[75];
  assign t[159] = t[200] ^ x[78];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[201] ^ x[81];
  assign t[161] = t[202] ^ x[84];
  assign t[162] = t[203] ^ x[87];
  assign t[163] = t[204] ^ x[90];
  assign t[164] = t[205] ^ x[93];
  assign t[165] = t[206] ^ x[96];
  assign t[166] = t[207] ^ x[99];
  assign t[167] = t[208] ^ x[102];
  assign t[168] = t[209] ^ x[105];
  assign t[169] = t[210] ^ x[108];
  assign t[16] = ~(t[137] & t[24]);
  assign t[170] = t[211] ^ x[111];
  assign t[171] = t[212] ^ x[114];
  assign t[172] = t[213] ^ x[117];
  assign t[173] = t[214] ^ x[120];
  assign t[174] = t[215] ^ x[123];
  assign t[175] = (x[0] & x[1]);
  assign t[176] = (x[4] & x[5]);
  assign t[177] = (x[7] & x[8]);
  assign t[178] = (x[10] & x[11]);
  assign t[179] = (x[13] & x[14]);
  assign t[17] = t[25] & t[26];
  assign t[180] = (x[16] & x[17]);
  assign t[181] = (x[19] & x[20]);
  assign t[182] = (x[22] & x[23]);
  assign t[183] = (x[25] & x[26]);
  assign t[184] = (x[28] & x[29]);
  assign t[185] = (x[31] & x[32]);
  assign t[186] = (x[34] & x[35]);
  assign t[187] = (x[37] & x[38]);
  assign t[188] = (x[40] & x[41]);
  assign t[189] = (x[43] & x[44]);
  assign t[18] = ~(t[138]);
  assign t[190] = (x[46] & x[47]);
  assign t[191] = (x[49] & x[50]);
  assign t[192] = (x[52] & x[53]);
  assign t[193] = (x[55] & x[56]);
  assign t[194] = (x[58] & x[59]);
  assign t[195] = (x[61] & x[62]);
  assign t[196] = (x[64] & x[65]);
  assign t[197] = (x[67] & x[68]);
  assign t[198] = (x[70] & x[71]);
  assign t[199] = (x[73] & x[74]);
  assign t[19] = ~(t[137]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[76] & x[77]);
  assign t[201] = (x[79] & x[80]);
  assign t[202] = (x[82] & x[83]);
  assign t[203] = (x[85] & x[86]);
  assign t[204] = (x[88] & x[89]);
  assign t[205] = (x[91] & x[92]);
  assign t[206] = (x[94] & x[95]);
  assign t[207] = (x[97] & x[98]);
  assign t[208] = (x[100] & x[101]);
  assign t[209] = (x[103] & x[104]);
  assign t[20] = ~(t[139]);
  assign t[210] = (x[106] & x[107]);
  assign t[211] = (x[109] & x[110]);
  assign t[212] = (x[112] & x[113]);
  assign t[213] = (x[115] & x[116]);
  assign t[214] = (x[118] & x[119]);
  assign t[215] = (x[121] & x[122]);
  assign t[21] = ~(t[140]);
  assign t[22] = t[27] ^ t[28];
  assign t[23] = t[29] ^ t[30];
  assign t[24] = ~(t[141] | t[31]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = t[36] & t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[6]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = ~(t[142] & t[143]);
  assign t[33] = ~(t[144] & t[145]);
  assign t[34] = ~(t[24]);
  assign t[35] = ~(t[146] & t[46]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = t[49] ^ t[50];
  assign t[38] = t[51] & t[52];
  assign t[39] = t[53] & t[54];
  assign t[3] = ~(t[7]);
  assign t[40] = t[55] & t[56];
  assign t[41] = t[57] ^ t[58];
  assign t[42] = t[51] & t[59];
  assign t[43] = t[53] & t[60];
  assign t[44] = ~(t[147] | t[148]);
  assign t[45] = ~(t[149] | t[150]);
  assign t[46] = ~(t[151]);
  assign t[47] = t[61] & t[62];
  assign t[48] = t[61] ^ t[63];
  assign t[49] = t[64] ^ t[65];
  assign t[4] = t[8] ? t[135] : x[3];
  assign t[50] = t[66] ^ t[67];
  assign t[51] = t[68] ^ t[69];
  assign t[52] = t[64] ^ t[70];
  assign t[53] = t[51] ^ t[71];
  assign t[54] = t[70] ^ t[65];
  assign t[55] = t[69] ^ t[36];
  assign t[56] = t[52] ^ t[72];
  assign t[57] = t[36] & t[73];
  assign t[58] = t[55] & t[74];
  assign t[59] = t[72] ^ t[75];
  assign t[5] = ~(t[9] ^ t[136]);
  assign t[60] = t[52] ^ t[76];
  assign t[61] = t[77] ^ t[78];
  assign t[62] = t[79] & t[77];
  assign t[63] = t[77] & t[80];
  assign t[64] = t[12] ? t[152] : t[81];
  assign t[65] = t[12] ? t[153] : t[82];
  assign t[66] = t[83] ^ t[84];
  assign t[67] = t[85] ^ t[86];
  assign t[68] = t[79] ^ t[87];
  assign t[69] = t[78] ^ t[88];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[12] ? t[154] : t[89];
  assign t[71] = t[90] ^ t[36];
  assign t[72] = t[91] ^ t[85];
  assign t[73] = t[86] ^ t[56];
  assign t[74] = t[92] ^ t[54];
  assign t[75] = t[83] ^ t[65];
  assign t[76] = t[84] ^ t[65];
  assign t[77] = t[93] ^ t[94];
  assign t[78] = t[95] ^ t[96];
  assign t[79] = t[97] ^ t[98];
  assign t[7] = ~(t[12]);
  assign t[80] = t[99] ^ t[94];
  assign t[81] = t[155] ^ t[156];
  assign t[82] = t[157] ^ t[158];
  assign t[83] = t[12] ? t[159] : t[100];
  assign t[84] = t[12] ? t[160] : t[101];
  assign t[85] = t[12] ? t[161] : t[102];
  assign t[86] = t[12] ? t[162] : t[103];
  assign t[87] = t[104] & t[105];
  assign t[88] = t[106] & t[61];
  assign t[89] = t[163] ^ t[164];
  assign t[8] = ~(t[13]);
  assign t[90] = t[107] ^ t[108];
  assign t[91] = t[12] ? t[165] : t[109];
  assign t[92] = t[64] ^ t[85];
  assign t[93] = t[110] ^ t[111];
  assign t[94] = t[112] ^ t[113];
  assign t[95] = t[114] ^ t[98];
  assign t[96] = t[115] ^ t[116];
  assign t[97] = t[117] ^ t[118];
  assign t[98] = t[119] ^ t[113];
  assign t[99] = t[120] ^ t[121];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = t[0] ? t[1] : t[134];
endmodule

module R1ind165(x, y);
 input [120:0] x;
 output y;

 wire [211:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[35] & t[49];
  assign t[101] = t[58] & t[57];
  assign t[102] = t[111] ^ t[86];
  assign t[103] = t[53] ^ t[112];
  assign t[104] = t[68] ^ t[79];
  assign t[105] = t[170] ^ t[171];
  assign t[106] = t[113] ^ t[114];
  assign t[107] = t[115] ^ t[101];
  assign t[108] = t[116] ^ t[117];
  assign t[109] = t[70] & t[73];
  assign t[10] = ~(t[16]);
  assign t[110] = t[118] & t[65];
  assign t[111] = t[119] ^ t[120];
  assign t[112] = t[121] ^ t[122];
  assign t[113] = t[123] ^ t[110];
  assign t[114] = t[124] & t[125];
  assign t[115] = t[126] & t[127];
  assign t[116] = t[128] ^ t[120];
  assign t[117] = t[129] & t[121];
  assign t[118] = t[51] ^ t[126];
  assign t[119] = t[53] & t[112];
  assign t[11] = t[135] & t[17];
  assign t[120] = t[51] & t[122];
  assign t[121] = t[73] ^ t[66];
  assign t[122] = t[74] ^ t[130];
  assign t[123] = t[65] ^ t[75];
  assign t[124] = t[35] ^ t[129];
  assign t[125] = t[73] ^ t[65];
  assign t[126] = t[76] ^ t[48];
  assign t[127] = t[58] ^ t[130];
  assign t[128] = t[51] ^ t[122];
  assign t[129] = t[66] ^ t[131];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[83] ^ t[48];
  assign t[131] = t[67] ^ t[73];
  assign t[132] = t[172] ^ x[2];
  assign t[133] = t[173] ^ x[6];
  assign t[134] = t[174] ^ x[9];
  assign t[135] = t[175] ^ x[12];
  assign t[136] = t[176] ^ x[15];
  assign t[137] = t[177] ^ x[18];
  assign t[138] = t[178] ^ x[21];
  assign t[139] = t[179] ^ x[24];
  assign t[13] = ~(t[135]);
  assign t[140] = t[180] ^ x[27];
  assign t[141] = t[181] ^ x[30];
  assign t[142] = t[182] ^ x[33];
  assign t[143] = t[183] ^ x[36];
  assign t[144] = t[184] ^ x[39];
  assign t[145] = t[185] ^ x[42];
  assign t[146] = t[186] ^ x[45];
  assign t[147] = t[187] ^ x[48];
  assign t[148] = t[188] ^ x[51];
  assign t[149] = t[189] ^ x[54];
  assign t[14] = t[136] & t[137];
  assign t[150] = t[190] ^ x[57];
  assign t[151] = t[191] ^ x[60];
  assign t[152] = t[192] ^ x[63];
  assign t[153] = t[193] ^ x[66];
  assign t[154] = t[194] ^ x[69];
  assign t[155] = t[195] ^ x[72];
  assign t[156] = t[196] ^ x[75];
  assign t[157] = t[197] ^ x[78];
  assign t[158] = t[198] ^ x[81];
  assign t[159] = t[199] ^ x[84];
  assign t[15] = ~(t[20] ^ t[21]);
  assign t[160] = t[200] ^ x[87];
  assign t[161] = t[201] ^ x[90];
  assign t[162] = t[202] ^ x[93];
  assign t[163] = t[203] ^ x[96];
  assign t[164] = t[204] ^ x[99];
  assign t[165] = t[205] ^ x[102];
  assign t[166] = t[206] ^ x[105];
  assign t[167] = t[207] ^ x[108];
  assign t[168] = t[208] ^ x[111];
  assign t[169] = t[209] ^ x[114];
  assign t[16] = ~(t[135] & t[22]);
  assign t[170] = t[210] ^ x[117];
  assign t[171] = t[211] ^ x[120];
  assign t[172] = (x[0] & x[1]);
  assign t[173] = (x[4] & x[5]);
  assign t[174] = (x[7] & x[8]);
  assign t[175] = (x[10] & x[11]);
  assign t[176] = (x[13] & x[14]);
  assign t[177] = (x[16] & x[17]);
  assign t[178] = (x[19] & x[20]);
  assign t[179] = (x[22] & x[23]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[25] & x[26]);
  assign t[181] = (x[28] & x[29]);
  assign t[182] = (x[31] & x[32]);
  assign t[183] = (x[34] & x[35]);
  assign t[184] = (x[37] & x[38]);
  assign t[185] = (x[40] & x[41]);
  assign t[186] = (x[43] & x[44]);
  assign t[187] = (x[46] & x[47]);
  assign t[188] = (x[49] & x[50]);
  assign t[189] = (x[52] & x[53]);
  assign t[18] = ~(t[138]);
  assign t[190] = (x[55] & x[56]);
  assign t[191] = (x[58] & x[59]);
  assign t[192] = (x[61] & x[62]);
  assign t[193] = (x[64] & x[65]);
  assign t[194] = (x[67] & x[68]);
  assign t[195] = (x[70] & x[71]);
  assign t[196] = (x[73] & x[74]);
  assign t[197] = (x[76] & x[77]);
  assign t[198] = (x[79] & x[80]);
  assign t[199] = (x[82] & x[83]);
  assign t[19] = ~(t[135]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[85] & x[86]);
  assign t[201] = (x[88] & x[89]);
  assign t[202] = (x[91] & x[92]);
  assign t[203] = (x[94] & x[95]);
  assign t[204] = (x[97] & x[98]);
  assign t[205] = (x[100] & x[101]);
  assign t[206] = (x[103] & x[104]);
  assign t[207] = (x[106] & x[107]);
  assign t[208] = (x[109] & x[110]);
  assign t[209] = (x[112] & x[113]);
  assign t[20] = t[25] ^ t[26];
  assign t[210] = (x[115] & x[116]);
  assign t[211] = (x[118] & x[119]);
  assign t[21] = t[27] ^ t[28];
  assign t[22] = ~(t[139] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = t[34] & t[35];
  assign t[26] = t[36] ^ t[37];
  assign t[27] = t[38] ^ t[39];
  assign t[28] = t[40] ^ t[41];
  assign t[29] = ~(t[42] & t[43]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[140] & t[136]);
  assign t[31] = ~(t[141] & t[142]);
  assign t[32] = ~(t[22]);
  assign t[33] = ~(t[143] & t[44]);
  assign t[34] = t[45] ^ t[46];
  assign t[35] = t[47] ^ t[48];
  assign t[36] = t[34] & t[49];
  assign t[37] = t[50] & t[51];
  assign t[38] = t[52] & t[53];
  assign t[39] = t[54] ^ t[55];
  assign t[3] = ~(t[7]);
  assign t[40] = t[56] & t[57];
  assign t[41] = t[56] & t[58];
  assign t[42] = ~(t[144] | t[145]);
  assign t[43] = ~(t[146] | t[147]);
  assign t[44] = ~(t[148]);
  assign t[45] = t[59] ^ t[60];
  assign t[46] = t[61] ^ t[62];
  assign t[47] = t[12] ? t[149] : t[63];
  assign t[48] = t[12] ? t[150] : t[64];
  assign t[49] = t[65] ^ t[66];
  assign t[4] = t[8] ? t[133] : x[3];
  assign t[50] = t[52] ^ t[45];
  assign t[51] = t[47] ^ t[67];
  assign t[52] = t[68] ^ t[69];
  assign t[53] = t[58] ^ t[70];
  assign t[54] = t[71] & t[65];
  assign t[55] = t[72] & t[73];
  assign t[56] = t[52] ^ t[72];
  assign t[57] = t[74] ^ t[75];
  assign t[58] = t[47] ^ t[76];
  assign t[59] = t[77] & t[78];
  assign t[5] = ~(t[9] ^ t[134]);
  assign t[60] = t[77] ^ t[79];
  assign t[61] = t[80] & t[81];
  assign t[62] = t[80] ^ t[79];
  assign t[63] = t[151] ^ t[152];
  assign t[64] = t[153] ^ t[154];
  assign t[65] = t[58] ^ t[74];
  assign t[66] = t[82] ^ t[83];
  assign t[67] = t[12] ? t[155] : t[84];
  assign t[68] = t[85] ^ t[86];
  assign t[69] = t[87] & t[77];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[66] ^ t[88];
  assign t[71] = t[72] ^ t[46];
  assign t[72] = t[89] ^ t[90];
  assign t[73] = t[12] ? t[156] : t[91];
  assign t[74] = t[92] ^ t[67];
  assign t[75] = t[82] ^ t[48];
  assign t[76] = t[12] ? t[157] : t[93];
  assign t[77] = t[94] ^ t[68];
  assign t[78] = t[94] & t[89];
  assign t[79] = t[95] & t[94];
  assign t[7] = ~(t[12]);
  assign t[80] = t[95] ^ t[89];
  assign t[81] = t[68] & t[95];
  assign t[82] = t[12] ? t[158] : t[96];
  assign t[83] = t[12] ? t[159] : t[97];
  assign t[84] = t[160] ^ t[161];
  assign t[85] = t[98] ^ t[99];
  assign t[86] = t[100] ^ t[101];
  assign t[87] = t[89] ^ t[79];
  assign t[88] = t[76] ^ t[73];
  assign t[89] = t[102] ^ t[103];
  assign t[8] = ~(t[13]);
  assign t[90] = t[104] & t[80];
  assign t[91] = t[162] ^ t[163];
  assign t[92] = t[12] ? t[164] : t[105];
  assign t[93] = t[165] ^ t[166];
  assign t[94] = t[106] ^ t[107];
  assign t[95] = t[108] ^ t[107];
  assign t[96] = t[167] ^ t[168];
  assign t[97] = t[169] ^ t[134];
  assign t[98] = t[109] ^ t[110];
  assign t[99] = t[35] ^ t[49];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = t[0] ? t[1] : t[132];
endmodule

module R1ind166(x, y);
 input [120:0] x;
 output y;

 wire [212:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[165] ^ t[166];
  assign t[101] = t[167] ^ t[168];
  assign t[102] = t[169] ^ t[170];
  assign t[103] = t[113] ^ t[114];
  assign t[104] = t[115] ^ t[114];
  assign t[105] = t[171] ^ t[172];
  assign t[106] = t[116] ^ t[117];
  assign t[107] = t[73] ^ t[118];
  assign t[108] = t[73] & t[118];
  assign t[109] = t[51] & t[119];
  assign t[10] = ~(t[16]);
  assign t[110] = t[120] ^ t[121];
  assign t[111] = t[51] ^ t[122];
  assign t[112] = t[53] ^ t[50];
  assign t[113] = t[123] ^ t[124];
  assign t[114] = t[125] ^ t[109];
  assign t[115] = t[126] ^ t[127];
  assign t[116] = t[122] & t[69];
  assign t[117] = t[76] & t[57];
  assign t[118] = t[57] ^ t[70];
  assign t[119] = t[64] ^ t[128];
  assign t[11] = t[136] & t[17];
  assign t[120] = t[111] & t[112];
  assign t[121] = t[93] & t[50];
  assign t[122] = t[70] ^ t[129];
  assign t[123] = t[130] ^ t[117];
  assign t[124] = t[55] & t[75];
  assign t[125] = t[35] & t[131];
  assign t[126] = t[132] ^ t[121];
  assign t[127] = t[74] & t[53];
  assign t[128] = t[89] ^ t[48];
  assign t[129] = t[47] ^ t[69];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[57] ^ t[128];
  assign t[131] = t[51] ^ t[65];
  assign t[132] = t[93] ^ t[50];
  assign t[133] = t[173] ^ x[2];
  assign t[134] = t[174] ^ x[6];
  assign t[135] = t[175] ^ x[9];
  assign t[136] = t[176] ^ x[12];
  assign t[137] = t[177] ^ x[15];
  assign t[138] = t[178] ^ x[18];
  assign t[139] = t[179] ^ x[21];
  assign t[13] = ~(t[136]);
  assign t[140] = t[180] ^ x[24];
  assign t[141] = t[181] ^ x[27];
  assign t[142] = t[182] ^ x[30];
  assign t[143] = t[183] ^ x[33];
  assign t[144] = t[184] ^ x[36];
  assign t[145] = t[185] ^ x[39];
  assign t[146] = t[186] ^ x[42];
  assign t[147] = t[187] ^ x[45];
  assign t[148] = t[188] ^ x[48];
  assign t[149] = t[189] ^ x[51];
  assign t[14] = t[137] & t[138];
  assign t[150] = t[190] ^ x[54];
  assign t[151] = t[191] ^ x[57];
  assign t[152] = t[192] ^ x[60];
  assign t[153] = t[193] ^ x[63];
  assign t[154] = t[194] ^ x[66];
  assign t[155] = t[195] ^ x[69];
  assign t[156] = t[196] ^ x[72];
  assign t[157] = t[197] ^ x[75];
  assign t[158] = t[198] ^ x[78];
  assign t[159] = t[199] ^ x[81];
  assign t[15] = t[20] ^ t[21];
  assign t[160] = t[200] ^ x[84];
  assign t[161] = t[201] ^ x[87];
  assign t[162] = t[202] ^ x[90];
  assign t[163] = t[203] ^ x[93];
  assign t[164] = t[204] ^ x[96];
  assign t[165] = t[205] ^ x[99];
  assign t[166] = t[206] ^ x[102];
  assign t[167] = t[207] ^ x[105];
  assign t[168] = t[208] ^ x[108];
  assign t[169] = t[209] ^ x[111];
  assign t[16] = ~(t[136] & t[22]);
  assign t[170] = t[210] ^ x[114];
  assign t[171] = t[211] ^ x[117];
  assign t[172] = t[212] ^ x[120];
  assign t[173] = (x[0] & x[1]);
  assign t[174] = (x[4] & x[5]);
  assign t[175] = (x[7] & x[8]);
  assign t[176] = (x[10] & x[11]);
  assign t[177] = (x[13] & x[14]);
  assign t[178] = (x[16] & x[17]);
  assign t[179] = (x[19] & x[20]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[22] & x[23]);
  assign t[181] = (x[25] & x[26]);
  assign t[182] = (x[28] & x[29]);
  assign t[183] = (x[31] & x[32]);
  assign t[184] = (x[34] & x[35]);
  assign t[185] = (x[37] & x[38]);
  assign t[186] = (x[40] & x[41]);
  assign t[187] = (x[43] & x[44]);
  assign t[188] = (x[46] & x[47]);
  assign t[189] = (x[49] & x[50]);
  assign t[18] = ~(t[139]);
  assign t[190] = (x[52] & x[53]);
  assign t[191] = (x[55] & x[56]);
  assign t[192] = (x[58] & x[59]);
  assign t[193] = (x[61] & x[62]);
  assign t[194] = (x[64] & x[65]);
  assign t[195] = (x[67] & x[68]);
  assign t[196] = (x[70] & x[71]);
  assign t[197] = (x[73] & x[74]);
  assign t[198] = (x[76] & x[77]);
  assign t[199] = (x[79] & x[80]);
  assign t[19] = ~(t[136]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[82] & x[83]);
  assign t[201] = (x[85] & x[86]);
  assign t[202] = (x[88] & x[89]);
  assign t[203] = (x[91] & x[92]);
  assign t[204] = (x[94] & x[95]);
  assign t[205] = (x[97] & x[98]);
  assign t[206] = (x[100] & x[101]);
  assign t[207] = (x[103] & x[104]);
  assign t[208] = (x[106] & x[107]);
  assign t[209] = (x[109] & x[110]);
  assign t[20] = t[25] ^ t[26];
  assign t[210] = (x[112] & x[113]);
  assign t[211] = (x[115] & x[116]);
  assign t[212] = (x[118] & x[119]);
  assign t[21] = t[27] ^ t[28];
  assign t[22] = ~(t[140] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = t[34] & t[35];
  assign t[26] = t[36] ^ t[37];
  assign t[27] = t[38] ^ t[39];
  assign t[28] = t[40] ^ t[41];
  assign t[29] = ~(t[42] & t[43]);
  assign t[2] = ~(t[6]);
  assign t[30] = ~(t[141] & t[142]);
  assign t[31] = ~(t[137] & t[143]);
  assign t[32] = ~(t[22]);
  assign t[33] = ~(t[144] & t[44]);
  assign t[34] = t[45] ^ t[46];
  assign t[35] = t[47] ^ t[48];
  assign t[36] = t[49] & t[50];
  assign t[37] = t[45] & t[51];
  assign t[38] = t[52] & t[53];
  assign t[39] = t[54] & t[55];
  assign t[3] = ~(t[7]);
  assign t[40] = t[56] & t[57];
  assign t[41] = t[58] ^ t[59];
  assign t[42] = ~(t[145] | t[146]);
  assign t[43] = ~(t[147] | t[148]);
  assign t[44] = ~(t[149]);
  assign t[45] = t[60] ^ t[61];
  assign t[46] = t[52] ^ t[54];
  assign t[47] = t[12] ? t[150] : t[62];
  assign t[48] = t[12] ? t[151] : t[63];
  assign t[49] = t[60] ^ t[52];
  assign t[4] = t[8] ? t[134] : x[3];
  assign t[50] = t[64] ^ t[65];
  assign t[51] = t[66] ^ t[47];
  assign t[52] = t[67] ^ t[68];
  assign t[53] = t[69] ^ t[70];
  assign t[54] = t[71] ^ t[72];
  assign t[55] = t[73] ^ t[74];
  assign t[56] = t[61] ^ t[54];
  assign t[57] = t[51] ^ t[64];
  assign t[58] = t[54] & t[75];
  assign t[59] = t[56] & t[76];
  assign t[5] = ~(t[9] ^ t[135]);
  assign t[60] = t[77] ^ t[78];
  assign t[61] = t[79] ^ t[80];
  assign t[62] = t[152] ^ t[135];
  assign t[63] = t[153] ^ t[154];
  assign t[64] = t[81] ^ t[82];
  assign t[65] = t[83] ^ t[48];
  assign t[66] = t[12] ? t[155] : t[84];
  assign t[67] = t[85] & t[86];
  assign t[68] = t[85] ^ t[87];
  assign t[69] = t[12] ? t[156] : t[88];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[89] ^ t[83];
  assign t[71] = t[90] & t[91];
  assign t[72] = t[90] ^ t[87];
  assign t[73] = t[66] ^ t[48];
  assign t[74] = t[70] ^ t[92];
  assign t[75] = t[69] ^ t[57];
  assign t[76] = t[93] ^ t[35];
  assign t[77] = t[94] ^ t[95];
  assign t[78] = t[96] & t[85];
  assign t[79] = t[97] ^ t[98];
  assign t[7] = ~(t[12]);
  assign t[80] = t[99] & t[90];
  assign t[81] = t[12] ? t[157] : t[100];
  assign t[82] = t[12] ? t[158] : t[101];
  assign t[83] = t[12] ? t[159] : t[102];
  assign t[84] = t[160] ^ t[161];
  assign t[85] = t[103] ^ t[77];
  assign t[86] = t[103] & t[79];
  assign t[87] = t[104] & t[103];
  assign t[88] = t[162] ^ t[163];
  assign t[89] = t[12] ? t[164] : t[105];
  assign t[8] = ~(t[13]);
  assign t[90] = t[104] ^ t[79];
  assign t[91] = t[77] & t[104];
  assign t[92] = t[82] ^ t[69];
  assign t[93] = t[66] ^ t[82];
  assign t[94] = t[106] ^ t[107];
  assign t[95] = t[108] ^ t[109];
  assign t[96] = t[79] ^ t[87];
  assign t[97] = t[110] ^ t[95];
  assign t[98] = t[111] ^ t[112];
  assign t[99] = t[77] ^ t[87];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = t[0] ? t[1] : t[133];
endmodule

module R1ind167(x, y);
 input [123:0] x;
 output y;

 wire [215:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[88] ^ t[65];
  assign t[101] = t[113] ^ t[114];
  assign t[102] = t[115] ^ t[114];
  assign t[103] = t[167] ^ t[168];
  assign t[104] = t[169] ^ t[170];
  assign t[105] = t[12] ? t[171] : t[116];
  assign t[106] = t[172] ^ t[173];
  assign t[107] = t[117] ^ t[118];
  assign t[108] = t[48] ^ t[119];
  assign t[109] = t[120] ^ t[121];
  assign t[10] = ~(t[16]);
  assign t[110] = t[71] ^ t[122];
  assign t[111] = t[71] & t[122];
  assign t[112] = t[48] & t[123];
  assign t[113] = t[124] ^ t[125];
  assign t[114] = t[126] ^ t[112];
  assign t[115] = t[127] ^ t[128];
  assign t[116] = t[174] ^ t[136];
  assign t[117] = t[108] & t[61];
  assign t[118] = t[74] & t[80];
  assign t[119] = t[68] ^ t[129];
  assign t[11] = t[137] & t[17];
  assign t[120] = t[119] & t[59];
  assign t[121] = t[57] & t[73];
  assign t[122] = t[73] ^ t[68];
  assign t[123] = t[92] ^ t[130];
  assign t[124] = t[131] ^ t[121];
  assign t[125] = t[54] & t[55];
  assign t[126] = t[50] & t[132];
  assign t[127] = t[133] ^ t[118];
  assign t[128] = t[72] & t[52];
  assign t[129] = t[63] ^ t[59];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[87] ^ t[65];
  assign t[131] = t[73] ^ t[130];
  assign t[132] = t[48] ^ t[100];
  assign t[133] = t[74] ^ t[80];
  assign t[134] = t[175] ^ x[2];
  assign t[135] = t[176] ^ x[6];
  assign t[136] = t[177] ^ x[9];
  assign t[137] = t[178] ^ x[12];
  assign t[138] = t[179] ^ x[15];
  assign t[139] = t[180] ^ x[18];
  assign t[13] = ~(t[137]);
  assign t[140] = t[181] ^ x[21];
  assign t[141] = t[182] ^ x[24];
  assign t[142] = t[183] ^ x[27];
  assign t[143] = t[184] ^ x[30];
  assign t[144] = t[185] ^ x[33];
  assign t[145] = t[186] ^ x[36];
  assign t[146] = t[187] ^ x[39];
  assign t[147] = t[188] ^ x[42];
  assign t[148] = t[189] ^ x[45];
  assign t[149] = t[190] ^ x[48];
  assign t[14] = ~(t[20] | t[21]);
  assign t[150] = t[191] ^ x[51];
  assign t[151] = t[192] ^ x[54];
  assign t[152] = t[193] ^ x[57];
  assign t[153] = t[194] ^ x[60];
  assign t[154] = t[195] ^ x[63];
  assign t[155] = t[196] ^ x[66];
  assign t[156] = t[197] ^ x[69];
  assign t[157] = t[198] ^ x[72];
  assign t[158] = t[199] ^ x[75];
  assign t[159] = t[200] ^ x[78];
  assign t[15] = t[22] ^ t[23];
  assign t[160] = t[201] ^ x[81];
  assign t[161] = t[202] ^ x[84];
  assign t[162] = t[203] ^ x[87];
  assign t[163] = t[204] ^ x[90];
  assign t[164] = t[205] ^ x[93];
  assign t[165] = t[206] ^ x[96];
  assign t[166] = t[207] ^ x[99];
  assign t[167] = t[208] ^ x[102];
  assign t[168] = t[209] ^ x[105];
  assign t[169] = t[210] ^ x[108];
  assign t[16] = ~(t[137] & t[24]);
  assign t[170] = t[211] ^ x[111];
  assign t[171] = t[212] ^ x[114];
  assign t[172] = t[213] ^ x[117];
  assign t[173] = t[214] ^ x[120];
  assign t[174] = t[215] ^ x[123];
  assign t[175] = (x[0] & x[1]);
  assign t[176] = (x[4] & x[5]);
  assign t[177] = (x[7] & x[8]);
  assign t[178] = (x[10] & x[11]);
  assign t[179] = (x[13] & x[14]);
  assign t[17] = t[25] & t[26];
  assign t[180] = (x[16] & x[17]);
  assign t[181] = (x[19] & x[20]);
  assign t[182] = (x[22] & x[23]);
  assign t[183] = (x[25] & x[26]);
  assign t[184] = (x[28] & x[29]);
  assign t[185] = (x[31] & x[32]);
  assign t[186] = (x[34] & x[35]);
  assign t[187] = (x[37] & x[38]);
  assign t[188] = (x[40] & x[41]);
  assign t[189] = (x[43] & x[44]);
  assign t[18] = ~(t[138]);
  assign t[190] = (x[46] & x[47]);
  assign t[191] = (x[49] & x[50]);
  assign t[192] = (x[52] & x[53]);
  assign t[193] = (x[55] & x[56]);
  assign t[194] = (x[58] & x[59]);
  assign t[195] = (x[61] & x[62]);
  assign t[196] = (x[64] & x[65]);
  assign t[197] = (x[67] & x[68]);
  assign t[198] = (x[70] & x[71]);
  assign t[199] = (x[73] & x[74]);
  assign t[19] = ~(t[137]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[76] & x[77]);
  assign t[201] = (x[79] & x[80]);
  assign t[202] = (x[82] & x[83]);
  assign t[203] = (x[85] & x[86]);
  assign t[204] = (x[88] & x[89]);
  assign t[205] = (x[91] & x[92]);
  assign t[206] = (x[94] & x[95]);
  assign t[207] = (x[97] & x[98]);
  assign t[208] = (x[100] & x[101]);
  assign t[209] = (x[103] & x[104]);
  assign t[20] = ~(t[139]);
  assign t[210] = (x[106] & x[107]);
  assign t[211] = (x[109] & x[110]);
  assign t[212] = (x[112] & x[113]);
  assign t[213] = (x[115] & x[116]);
  assign t[214] = (x[118] & x[119]);
  assign t[215] = (x[121] & x[122]);
  assign t[21] = ~(t[140]);
  assign t[22] = t[27] ^ t[28];
  assign t[23] = t[29] ^ t[30];
  assign t[24] = ~(t[141] | t[31]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[6]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = ~(t[142] & t[143]);
  assign t[33] = ~(t[144] & t[145]);
  assign t[34] = ~(t[24]);
  assign t[35] = ~(t[146] & t[46]);
  assign t[36] = t[47] & t[48];
  assign t[37] = t[49] & t[50];
  assign t[38] = t[51] & t[52];
  assign t[39] = t[53] & t[54];
  assign t[3] = ~(t[7]);
  assign t[40] = t[53] & t[55];
  assign t[41] = t[56] & t[57];
  assign t[42] = t[58] & t[59];
  assign t[43] = t[60] & t[61];
  assign t[44] = ~(t[147] | t[148]);
  assign t[45] = ~(t[149] | t[150]);
  assign t[46] = ~(t[151]);
  assign t[47] = t[60] ^ t[58];
  assign t[48] = t[62] ^ t[63];
  assign t[49] = t[47] ^ t[64];
  assign t[4] = t[8] ? t[135] : x[3];
  assign t[50] = t[63] ^ t[65];
  assign t[51] = t[66] ^ t[67];
  assign t[52] = t[59] ^ t[68];
  assign t[53] = t[69] ^ t[70];
  assign t[54] = t[71] ^ t[72];
  assign t[55] = t[59] ^ t[73];
  assign t[56] = t[58] ^ t[53];
  assign t[57] = t[74] ^ t[50];
  assign t[58] = t[75] ^ t[76];
  assign t[59] = t[12] ? t[152] : t[77];
  assign t[5] = ~(t[9] ^ t[136]);
  assign t[60] = t[78] ^ t[79];
  assign t[61] = t[52] ^ t[80];
  assign t[62] = t[12] ? t[153] : t[81];
  assign t[63] = t[12] ? t[154] : t[82];
  assign t[64] = t[51] ^ t[53];
  assign t[65] = t[12] ? t[155] : t[83];
  assign t[66] = t[84] & t[85];
  assign t[67] = t[84] ^ t[86];
  assign t[68] = t[87] ^ t[88];
  assign t[69] = t[89] & t[90];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[89] ^ t[86];
  assign t[71] = t[62] ^ t[65];
  assign t[72] = t[68] ^ t[91];
  assign t[73] = t[48] ^ t[92];
  assign t[74] = t[62] ^ t[93];
  assign t[75] = t[94] ^ t[95];
  assign t[76] = t[96] & t[89];
  assign t[77] = t[156] ^ t[157];
  assign t[78] = t[97] ^ t[98];
  assign t[79] = t[99] & t[84];
  assign t[7] = ~(t[12]);
  assign t[80] = t[92] ^ t[100];
  assign t[81] = t[158] ^ t[159];
  assign t[82] = t[160] ^ t[161];
  assign t[83] = t[162] ^ t[163];
  assign t[84] = t[101] ^ t[78];
  assign t[85] = t[101] & t[75];
  assign t[86] = t[102] & t[101];
  assign t[87] = t[12] ? t[164] : t[103];
  assign t[88] = t[12] ? t[165] : t[104];
  assign t[89] = t[102] ^ t[75];
  assign t[8] = ~(t[13]);
  assign t[90] = t[78] & t[102];
  assign t[91] = t[93] ^ t[59];
  assign t[92] = t[105] ^ t[93];
  assign t[93] = t[12] ? t[166] : t[106];
  assign t[94] = t[107] ^ t[98];
  assign t[95] = t[108] ^ t[61];
  assign t[96] = t[78] ^ t[86];
  assign t[97] = t[109] ^ t[110];
  assign t[98] = t[111] ^ t[112];
  assign t[99] = t[75] ^ t[86];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = t[0] ? t[1] : t[134];
endmodule

module R1ind168(x, y);
 input [120:0] x;
 output y;

 wire [222:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[12] ? t[171] : t[120];
  assign t[101] = t[94] & t[121];
  assign t[102] = t[94] ^ t[115];
  assign t[103] = t[99] & t[122];
  assign t[104] = t[99] ^ t[115];
  assign t[105] = t[88] ^ t[65];
  assign t[106] = t[79] ^ t[123];
  assign t[107] = t[12] ? t[172] : t[124];
  assign t[108] = t[173] ^ t[174];
  assign t[109] = t[175] ^ t[176];
  assign t[10] = ~(t[16]);
  assign t[110] = t[177] ^ t[178];
  assign t[111] = t[125] ^ t[126];
  assign t[112] = t[105] ^ t[70];
  assign t[113] = t[105] & t[70];
  assign t[114] = t[68] & t[127];
  assign t[115] = t[119] & t[116];
  assign t[116] = t[128] ^ t[129];
  assign t[117] = t[130] ^ t[131];
  assign t[118] = t[82] ^ t[67];
  assign t[119] = t[132] ^ t[129];
  assign t[11] = t[146] & t[17];
  assign t[120] = t[179] ^ t[180];
  assign t[121] = t[116] & t[77];
  assign t[122] = t[72] & t[119];
  assign t[123] = t[90] ^ t[76];
  assign t[124] = t[181] ^ t[182];
  assign t[125] = t[59] & t[76];
  assign t[126] = t[133] & t[75];
  assign t[127] = t[87] ^ t[134];
  assign t[128] = t[135] ^ t[136];
  assign t[129] = t[137] ^ t[114];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[55] & t[118];
  assign t[131] = t[71] & t[67];
  assign t[132] = t[138] ^ t[139];
  assign t[133] = t[71] ^ t[48];
  assign t[134] = t[100] ^ t[65];
  assign t[135] = t[140] ^ t[126];
  assign t[136] = t[84] & t[141];
  assign t[137] = t[48] & t[51];
  assign t[138] = t[142] ^ t[131];
  assign t[139] = t[106] & t[82];
  assign t[13] = ~(t[146]);
  assign t[140] = t[75] ^ t[134];
  assign t[141] = t[76] ^ t[75];
  assign t[142] = t[71] ^ t[67];
  assign t[143] = t[183] ^ x[2];
  assign t[144] = t[184] ^ x[6];
  assign t[145] = t[185] ^ x[9];
  assign t[146] = t[186] ^ x[12];
  assign t[147] = t[187] ^ x[15];
  assign t[148] = t[188] ^ x[18];
  assign t[149] = t[189] ^ x[21];
  assign t[14] = ~(t[20] | t[21]);
  assign t[150] = t[190] ^ x[24];
  assign t[151] = t[191] ^ x[27];
  assign t[152] = t[192] ^ x[30];
  assign t[153] = t[193] ^ x[33];
  assign t[154] = t[194] ^ x[36];
  assign t[155] = t[195] ^ x[39];
  assign t[156] = t[196] ^ x[42];
  assign t[157] = t[197] ^ x[45];
  assign t[158] = t[198] ^ x[48];
  assign t[159] = t[199] ^ x[51];
  assign t[15] = t[22] ^ t[23];
  assign t[160] = t[200] ^ x[54];
  assign t[161] = t[201] ^ x[57];
  assign t[162] = t[202] ^ x[60];
  assign t[163] = t[203] ^ x[63];
  assign t[164] = t[204] ^ x[66];
  assign t[165] = t[205] ^ x[69];
  assign t[166] = t[206] ^ x[72];
  assign t[167] = t[207] ^ x[75];
  assign t[168] = t[208] ^ x[78];
  assign t[169] = t[209] ^ x[81];
  assign t[16] = ~(t[146] & t[24]);
  assign t[170] = t[210] ^ x[84];
  assign t[171] = t[211] ^ x[87];
  assign t[172] = t[212] ^ x[90];
  assign t[173] = t[213] ^ x[93];
  assign t[174] = t[214] ^ x[96];
  assign t[175] = t[215] ^ x[99];
  assign t[176] = t[216] ^ x[102];
  assign t[177] = t[217] ^ x[105];
  assign t[178] = t[218] ^ x[108];
  assign t[179] = t[219] ^ x[111];
  assign t[17] = t[25] & t[26];
  assign t[180] = t[220] ^ x[114];
  assign t[181] = t[221] ^ x[117];
  assign t[182] = t[222] ^ x[120];
  assign t[183] = (x[0] & x[1]);
  assign t[184] = (x[4] & x[5]);
  assign t[185] = (x[7] & x[8]);
  assign t[186] = (x[10] & x[11]);
  assign t[187] = (x[13] & x[14]);
  assign t[188] = (x[16] & x[17]);
  assign t[189] = (x[19] & x[20]);
  assign t[18] = ~(t[147]);
  assign t[190] = (x[22] & x[23]);
  assign t[191] = (x[25] & x[26]);
  assign t[192] = (x[28] & x[29]);
  assign t[193] = (x[31] & x[32]);
  assign t[194] = (x[34] & x[35]);
  assign t[195] = (x[37] & x[38]);
  assign t[196] = (x[40] & x[41]);
  assign t[197] = (x[43] & x[44]);
  assign t[198] = (x[46] & x[47]);
  assign t[199] = (x[49] & x[50]);
  assign t[19] = ~(t[146]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[52] & x[53]);
  assign t[201] = (x[55] & x[56]);
  assign t[202] = (x[58] & x[59]);
  assign t[203] = (x[61] & x[62]);
  assign t[204] = (x[64] & x[65]);
  assign t[205] = (x[67] & x[68]);
  assign t[206] = (x[70] & x[71]);
  assign t[207] = (x[73] & x[74]);
  assign t[208] = (x[76] & x[77]);
  assign t[209] = (x[79] & x[80]);
  assign t[20] = ~(t[148]);
  assign t[210] = (x[82] & x[83]);
  assign t[211] = (x[85] & x[86]);
  assign t[212] = (x[88] & x[89]);
  assign t[213] = (x[91] & x[92]);
  assign t[214] = (x[94] & x[95]);
  assign t[215] = (x[97] & x[98]);
  assign t[216] = (x[100] & x[101]);
  assign t[217] = (x[103] & x[104]);
  assign t[218] = (x[106] & x[107]);
  assign t[219] = (x[109] & x[110]);
  assign t[21] = ~(t[149]);
  assign t[220] = (x[112] & x[113]);
  assign t[221] = (x[115] & x[116]);
  assign t[222] = (x[118] & x[119]);
  assign t[22] = t[27] ^ t[28];
  assign t[23] = t[29] ^ t[30];
  assign t[24] = ~(t[150] | t[31]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[6]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = ~(t[151] & t[152]);
  assign t[33] = ~(t[153] & t[148]);
  assign t[34] = ~(t[24]);
  assign t[35] = ~(t[154] & t[46]);
  assign t[36] = t[47] & t[48];
  assign t[37] = t[49] ^ t[50];
  assign t[38] = t[47] & t[51];
  assign t[39] = t[52] ^ t[53];
  assign t[3] = ~(t[7]);
  assign t[40] = t[54] & t[55];
  assign t[41] = t[56] ^ t[57];
  assign t[42] = t[58] & t[59];
  assign t[43] = t[60] ^ t[61];
  assign t[44] = ~(t[155] | t[156]);
  assign t[45] = ~(t[157] | t[158]);
  assign t[46] = ~(t[159]);
  assign t[47] = t[62] ^ t[63];
  assign t[48] = t[64] ^ t[65];
  assign t[49] = t[66] & t[67];
  assign t[4] = t[8] ? t[144] : x[3];
  assign t[50] = t[62] & t[68];
  assign t[51] = t[68] ^ t[69];
  assign t[52] = t[63] & t[70];
  assign t[53] = t[66] & t[71];
  assign t[54] = t[72] ^ t[73];
  assign t[55] = t[68] ^ t[59];
  assign t[56] = t[74] & t[75];
  assign t[57] = t[58] & t[76];
  assign t[58] = t[77] ^ t[78];
  assign t[59] = t[79] ^ t[80];
  assign t[5] = ~(t[9] ^ t[145]);
  assign t[60] = t[81] & t[82];
  assign t[61] = t[83] & t[84];
  assign t[62] = t[54] ^ t[58];
  assign t[63] = t[81] ^ t[83];
  assign t[64] = t[12] ? t[160] : t[85];
  assign t[65] = t[12] ? t[161] : t[86];
  assign t[66] = t[54] ^ t[81];
  assign t[67] = t[87] ^ t[69];
  assign t[68] = t[88] ^ t[64];
  assign t[69] = t[89] ^ t[65];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[75] ^ t[79];
  assign t[71] = t[88] ^ t[90];
  assign t[72] = t[91] ^ t[92];
  assign t[73] = t[93] & t[94];
  assign t[74] = t[58] ^ t[83];
  assign t[75] = t[68] ^ t[87];
  assign t[76] = t[12] ? t[162] : t[95];
  assign t[77] = t[96] ^ t[97];
  assign t[78] = t[98] & t[99];
  assign t[79] = t[100] ^ t[89];
  assign t[7] = ~(t[12]);
  assign t[80] = t[64] ^ t[76];
  assign t[81] = t[101] ^ t[102];
  assign t[82] = t[76] ^ t[79];
  assign t[83] = t[103] ^ t[104];
  assign t[84] = t[105] ^ t[106];
  assign t[85] = t[163] ^ t[164];
  assign t[86] = t[165] ^ t[145];
  assign t[87] = t[107] ^ t[90];
  assign t[88] = t[12] ? t[166] : t[108];
  assign t[89] = t[12] ? t[167] : t[109];
  assign t[8] = ~(t[13]);
  assign t[90] = t[12] ? t[168] : t[110];
  assign t[91] = t[111] ^ t[112];
  assign t[92] = t[113] ^ t[114];
  assign t[93] = t[77] ^ t[115];
  assign t[94] = t[116] ^ t[72];
  assign t[95] = t[169] ^ t[170];
  assign t[96] = t[117] ^ t[92];
  assign t[97] = t[55] ^ t[118];
  assign t[98] = t[72] ^ t[115];
  assign t[99] = t[119] ^ t[77];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = t[0] ? t[1] : t[143];
endmodule

module R1ind169(x, y);
 input [120:0] x;
 output y;

 wire [213:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[116] ^ t[117];
  assign t[101] = t[72] ^ t[63];
  assign t[102] = t[82] ^ t[81];
  assign t[103] = t[102] & t[118];
  assign t[104] = t[102] ^ t[63];
  assign t[105] = t[119] ^ t[120];
  assign t[106] = t[121] ^ t[77];
  assign t[107] = t[121] & t[77];
  assign t[108] = t[52] & t[122];
  assign t[109] = t[12] ? t[170] : t[123];
  assign t[10] = ~(t[16]);
  assign t[110] = t[171] ^ t[136];
  assign t[111] = t[124] ^ t[120];
  assign t[112] = t[125] & t[126];
  assign t[113] = t[54] & t[58];
  assign t[114] = t[127] ^ t[128];
  assign t[115] = t[52] ^ t[129];
  assign t[116] = t[130] ^ t[128];
  assign t[117] = t[57] & t[37];
  assign t[118] = t[72] & t[82];
  assign t[119] = t[129] & t[49];
  assign t[11] = t[137] & t[17];
  assign t[120] = t[131] & t[95];
  assign t[121] = t[68] ^ t[71];
  assign t[122] = t[93] ^ t[132];
  assign t[123] = t[172] ^ t[173];
  assign t[124] = t[95] ^ t[132];
  assign t[125] = t[121] ^ t[57];
  assign t[126] = t[49] ^ t[95];
  assign t[127] = t[115] & t[56];
  assign t[128] = t[79] & t[74];
  assign t[129] = t[50] ^ t[133];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[79] ^ t[74];
  assign t[131] = t[79] ^ t[54];
  assign t[132] = t[65] ^ t[71];
  assign t[133] = t[69] ^ t[49];
  assign t[134] = t[174] ^ x[2];
  assign t[135] = t[175] ^ x[6];
  assign t[136] = t[176] ^ x[9];
  assign t[137] = t[177] ^ x[12];
  assign t[138] = t[178] ^ x[15];
  assign t[139] = t[179] ^ x[18];
  assign t[13] = ~(t[137]);
  assign t[140] = t[180] ^ x[21];
  assign t[141] = t[181] ^ x[24];
  assign t[142] = t[182] ^ x[27];
  assign t[143] = t[183] ^ x[30];
  assign t[144] = t[184] ^ x[33];
  assign t[145] = t[185] ^ x[36];
  assign t[146] = t[186] ^ x[39];
  assign t[147] = t[187] ^ x[42];
  assign t[148] = t[188] ^ x[45];
  assign t[149] = t[189] ^ x[48];
  assign t[14] = ~(t[20] | t[21]);
  assign t[150] = t[190] ^ x[51];
  assign t[151] = t[191] ^ x[54];
  assign t[152] = t[192] ^ x[57];
  assign t[153] = t[193] ^ x[60];
  assign t[154] = t[194] ^ x[63];
  assign t[155] = t[195] ^ x[66];
  assign t[156] = t[196] ^ x[69];
  assign t[157] = t[197] ^ x[72];
  assign t[158] = t[198] ^ x[75];
  assign t[159] = t[199] ^ x[78];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[200] ^ x[81];
  assign t[161] = t[201] ^ x[84];
  assign t[162] = t[202] ^ x[87];
  assign t[163] = t[203] ^ x[90];
  assign t[164] = t[204] ^ x[93];
  assign t[165] = t[205] ^ x[96];
  assign t[166] = t[206] ^ x[99];
  assign t[167] = t[207] ^ x[102];
  assign t[168] = t[208] ^ x[105];
  assign t[169] = t[209] ^ x[108];
  assign t[16] = ~(t[137] & t[24]);
  assign t[170] = t[210] ^ x[111];
  assign t[171] = t[211] ^ x[114];
  assign t[172] = t[212] ^ x[117];
  assign t[173] = t[213] ^ x[120];
  assign t[174] = (x[0] & x[1]);
  assign t[175] = (x[4] & x[5]);
  assign t[176] = (x[7] & x[8]);
  assign t[177] = (x[10] & x[11]);
  assign t[178] = (x[13] & x[14]);
  assign t[179] = (x[16] & x[17]);
  assign t[17] = t[25] & t[26];
  assign t[180] = (x[19] & x[20]);
  assign t[181] = (x[22] & x[23]);
  assign t[182] = (x[25] & x[26]);
  assign t[183] = (x[28] & x[29]);
  assign t[184] = (x[31] & x[32]);
  assign t[185] = (x[34] & x[35]);
  assign t[186] = (x[37] & x[38]);
  assign t[187] = (x[40] & x[41]);
  assign t[188] = (x[43] & x[44]);
  assign t[189] = (x[46] & x[47]);
  assign t[18] = ~(t[138]);
  assign t[190] = (x[49] & x[50]);
  assign t[191] = (x[52] & x[53]);
  assign t[192] = (x[55] & x[56]);
  assign t[193] = (x[58] & x[59]);
  assign t[194] = (x[61] & x[62]);
  assign t[195] = (x[64] & x[65]);
  assign t[196] = (x[67] & x[68]);
  assign t[197] = (x[70] & x[71]);
  assign t[198] = (x[73] & x[74]);
  assign t[199] = (x[76] & x[77]);
  assign t[19] = ~(t[137]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[79] & x[80]);
  assign t[201] = (x[82] & x[83]);
  assign t[202] = (x[85] & x[86]);
  assign t[203] = (x[88] & x[89]);
  assign t[204] = (x[91] & x[92]);
  assign t[205] = (x[94] & x[95]);
  assign t[206] = (x[97] & x[98]);
  assign t[207] = (x[100] & x[101]);
  assign t[208] = (x[103] & x[104]);
  assign t[209] = (x[106] & x[107]);
  assign t[20] = ~(t[139]);
  assign t[210] = (x[109] & x[110]);
  assign t[211] = (x[112] & x[113]);
  assign t[212] = (x[115] & x[116]);
  assign t[213] = (x[118] & x[119]);
  assign t[21] = ~(t[140]);
  assign t[22] = t[27] ^ t[28];
  assign t[23] = t[29] ^ t[30];
  assign t[24] = ~(t[141] | t[31]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = t[36] & t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[6]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = ~(t[139] & t[142]);
  assign t[33] = ~(t[143] & t[144]);
  assign t[34] = ~(t[24]);
  assign t[35] = ~(t[145] & t[46]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = t[49] ^ t[50];
  assign t[38] = t[51] & t[52];
  assign t[39] = t[53] & t[54];
  assign t[3] = ~(t[7]);
  assign t[40] = t[55] & t[56];
  assign t[41] = t[36] & t[57];
  assign t[42] = t[53] & t[58];
  assign t[43] = t[59] ^ t[60];
  assign t[44] = ~(t[146] | t[147]);
  assign t[45] = ~(t[148] | t[149]);
  assign t[46] = ~(t[150]);
  assign t[47] = t[61] & t[62];
  assign t[48] = t[61] ^ t[63];
  assign t[49] = t[12] ? t[151] : t[64];
  assign t[4] = t[8] ? t[135] : x[3];
  assign t[50] = t[65] ^ t[66];
  assign t[51] = t[55] ^ t[67];
  assign t[52] = t[68] ^ t[69];
  assign t[53] = t[51] ^ t[70];
  assign t[54] = t[69] ^ t[71];
  assign t[55] = t[72] ^ t[73];
  assign t[56] = t[37] ^ t[74];
  assign t[57] = t[50] ^ t[75];
  assign t[58] = t[52] ^ t[76];
  assign t[59] = t[70] & t[77];
  assign t[5] = ~(t[9] ^ t[136]);
  assign t[60] = t[78] & t[79];
  assign t[61] = t[80] ^ t[72];
  assign t[62] = t[80] & t[81];
  assign t[63] = t[82] & t[80];
  assign t[64] = t[152] ^ t[153];
  assign t[65] = t[12] ? t[154] : t[83];
  assign t[66] = t[12] ? t[155] : t[84];
  assign t[67] = t[81] ^ t[85];
  assign t[68] = t[12] ? t[156] : t[86];
  assign t[69] = t[12] ? t[157] : t[87];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[36] ^ t[88];
  assign t[71] = t[12] ? t[158] : t[89];
  assign t[72] = t[90] ^ t[91];
  assign t[73] = t[92] & t[61];
  assign t[74] = t[93] ^ t[76];
  assign t[75] = t[94] ^ t[49];
  assign t[76] = t[66] ^ t[71];
  assign t[77] = t[95] ^ t[50];
  assign t[78] = t[55] ^ t[36];
  assign t[79] = t[68] ^ t[94];
  assign t[7] = ~(t[12]);
  assign t[80] = t[96] ^ t[97];
  assign t[81] = t[98] ^ t[99];
  assign t[82] = t[100] ^ t[97];
  assign t[83] = t[159] ^ t[160];
  assign t[84] = t[161] ^ t[162];
  assign t[85] = t[101] & t[102];
  assign t[86] = t[163] ^ t[164];
  assign t[87] = t[165] ^ t[166];
  assign t[88] = t[103] ^ t[104];
  assign t[89] = t[167] ^ t[168];
  assign t[8] = ~(t[13]);
  assign t[90] = t[105] ^ t[106];
  assign t[91] = t[107] ^ t[108];
  assign t[92] = t[81] ^ t[63];
  assign t[93] = t[109] ^ t[94];
  assign t[94] = t[12] ? t[169] : t[110];
  assign t[95] = t[52] ^ t[93];
  assign t[96] = t[111] ^ t[112];
  assign t[97] = t[113] ^ t[108];
  assign t[98] = t[114] ^ t[91];
  assign t[99] = t[115] ^ t[56];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = t[0] ? t[1] : t[134];
endmodule

module R1ind170(x, y);
 input [123:0] x;
 output y;

 wire [216:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[171] ^ t[172];
  assign t[101] = t[12] ? t[173] : t[110];
  assign t[102] = t[111] ^ t[112];
  assign t[103] = t[53] ^ t[113];
  assign t[104] = t[114] ^ t[115];
  assign t[105] = t[116] ^ t[117];
  assign t[106] = t[118] ^ t[119];
  assign t[107] = t[118] & t[119];
  assign t[108] = t[53] & t[120];
  assign t[109] = t[121] ^ t[115];
  assign t[10] = ~(t[16]);
  assign t[110] = t[174] ^ t[175];
  assign t[111] = t[103] & t[70];
  assign t[112] = t[54] & t[52];
  assign t[113] = t[86] ^ t[122];
  assign t[114] = t[123] ^ t[124];
  assign t[115] = t[125] ^ t[108];
  assign t[116] = t[113] & t[60];
  assign t[117] = t[126] & t[58];
  assign t[118] = t[68] ^ t[50];
  assign t[119] = t[58] ^ t[86];
  assign t[11] = t[138] & t[17];
  assign t[120] = t[66] ^ t[127];
  assign t[121] = t[128] ^ t[129];
  assign t[122] = t[49] ^ t[60];
  assign t[123] = t[130] ^ t[112];
  assign t[124] = t[71] & t[85];
  assign t[125] = t[37] & t[131];
  assign t[126] = t[54] ^ t[37];
  assign t[127] = t[101] ^ t[50];
  assign t[128] = t[132] ^ t[117];
  assign t[129] = t[133] & t[134];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[54] ^ t[52];
  assign t[131] = t[53] ^ t[67];
  assign t[132] = t[58] ^ t[127];
  assign t[133] = t[118] ^ t[71];
  assign t[134] = t[60] ^ t[58];
  assign t[135] = t[176] ^ x[2];
  assign t[136] = t[177] ^ x[6];
  assign t[137] = t[178] ^ x[9];
  assign t[138] = t[179] ^ x[12];
  assign t[139] = t[180] ^ x[15];
  assign t[13] = ~(t[138]);
  assign t[140] = t[181] ^ x[18];
  assign t[141] = t[182] ^ x[21];
  assign t[142] = t[183] ^ x[24];
  assign t[143] = t[184] ^ x[27];
  assign t[144] = t[185] ^ x[30];
  assign t[145] = t[186] ^ x[33];
  assign t[146] = t[187] ^ x[36];
  assign t[147] = t[188] ^ x[39];
  assign t[148] = t[189] ^ x[42];
  assign t[149] = t[190] ^ x[45];
  assign t[14] = ~(t[20] | t[21]);
  assign t[150] = t[191] ^ x[48];
  assign t[151] = t[192] ^ x[51];
  assign t[152] = t[193] ^ x[54];
  assign t[153] = t[194] ^ x[57];
  assign t[154] = t[195] ^ x[60];
  assign t[155] = t[196] ^ x[63];
  assign t[156] = t[197] ^ x[66];
  assign t[157] = t[198] ^ x[69];
  assign t[158] = t[199] ^ x[72];
  assign t[159] = t[200] ^ x[75];
  assign t[15] = ~(t[22] ^ t[23]);
  assign t[160] = t[201] ^ x[78];
  assign t[161] = t[202] ^ x[81];
  assign t[162] = t[203] ^ x[84];
  assign t[163] = t[204] ^ x[87];
  assign t[164] = t[205] ^ x[90];
  assign t[165] = t[206] ^ x[93];
  assign t[166] = t[207] ^ x[96];
  assign t[167] = t[208] ^ x[99];
  assign t[168] = t[209] ^ x[102];
  assign t[169] = t[210] ^ x[105];
  assign t[16] = ~(t[138] & t[24]);
  assign t[170] = t[211] ^ x[108];
  assign t[171] = t[212] ^ x[111];
  assign t[172] = t[213] ^ x[114];
  assign t[173] = t[214] ^ x[117];
  assign t[174] = t[215] ^ x[120];
  assign t[175] = t[216] ^ x[123];
  assign t[176] = (x[0] & x[1]);
  assign t[177] = (x[4] & x[5]);
  assign t[178] = (x[7] & x[8]);
  assign t[179] = (x[10] & x[11]);
  assign t[17] = t[25] & t[26];
  assign t[180] = (x[13] & x[14]);
  assign t[181] = (x[16] & x[17]);
  assign t[182] = (x[19] & x[20]);
  assign t[183] = (x[22] & x[23]);
  assign t[184] = (x[25] & x[26]);
  assign t[185] = (x[28] & x[29]);
  assign t[186] = (x[31] & x[32]);
  assign t[187] = (x[34] & x[35]);
  assign t[188] = (x[37] & x[38]);
  assign t[189] = (x[40] & x[41]);
  assign t[18] = ~(t[139]);
  assign t[190] = (x[43] & x[44]);
  assign t[191] = (x[46] & x[47]);
  assign t[192] = (x[49] & x[50]);
  assign t[193] = (x[52] & x[53]);
  assign t[194] = (x[55] & x[56]);
  assign t[195] = (x[58] & x[59]);
  assign t[196] = (x[61] & x[62]);
  assign t[197] = (x[64] & x[65]);
  assign t[198] = (x[67] & x[68]);
  assign t[199] = (x[70] & x[71]);
  assign t[19] = ~(t[138]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[200] = (x[73] & x[74]);
  assign t[201] = (x[76] & x[77]);
  assign t[202] = (x[79] & x[80]);
  assign t[203] = (x[82] & x[83]);
  assign t[204] = (x[85] & x[86]);
  assign t[205] = (x[88] & x[89]);
  assign t[206] = (x[91] & x[92]);
  assign t[207] = (x[94] & x[95]);
  assign t[208] = (x[97] & x[98]);
  assign t[209] = (x[100] & x[101]);
  assign t[20] = ~(t[140]);
  assign t[210] = (x[103] & x[104]);
  assign t[211] = (x[106] & x[107]);
  assign t[212] = (x[109] & x[110]);
  assign t[213] = (x[112] & x[113]);
  assign t[214] = (x[115] & x[116]);
  assign t[215] = (x[118] & x[119]);
  assign t[216] = (x[121] & x[122]);
  assign t[21] = ~(t[141]);
  assign t[22] = t[27] ^ t[28];
  assign t[23] = t[29] ^ t[30];
  assign t[24] = ~(t[142] | t[31]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = t[36] & t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[6]);
  assign t[30] = t[42] ^ t[43];
  assign t[31] = ~(t[44] & t[45]);
  assign t[32] = ~(t[143] & t[144]);
  assign t[33] = ~(t[145] & t[146]);
  assign t[34] = ~(t[24]);
  assign t[35] = ~(t[147] & t[46]);
  assign t[36] = t[47] ^ t[48];
  assign t[37] = t[49] ^ t[50];
  assign t[38] = t[51] & t[52];
  assign t[39] = t[47] & t[53];
  assign t[3] = ~(t[7]);
  assign t[40] = t[51] & t[54];
  assign t[41] = t[55] ^ t[56];
  assign t[42] = t[57] & t[58];
  assign t[43] = t[59] & t[60];
  assign t[44] = ~(t[148] | t[149]);
  assign t[45] = ~(t[150] | t[151]);
  assign t[46] = ~(t[152]);
  assign t[47] = t[61] ^ t[59];
  assign t[48] = t[62] ^ t[63];
  assign t[49] = t[12] ? t[153] : t[64];
  assign t[4] = t[8] ? t[136] : x[3];
  assign t[50] = t[12] ? t[154] : t[65];
  assign t[51] = t[61] ^ t[62];
  assign t[52] = t[66] ^ t[67];
  assign t[53] = t[68] ^ t[49];
  assign t[54] = t[68] ^ t[69];
  assign t[55] = t[61] & t[70];
  assign t[56] = t[62] & t[71];
  assign t[57] = t[59] ^ t[63];
  assign t[58] = t[53] ^ t[66];
  assign t[59] = t[72] ^ t[73];
  assign t[5] = ~(t[9] ^ t[137]);
  assign t[60] = t[12] ? t[155] : t[74];
  assign t[61] = t[75] ^ t[76];
  assign t[62] = t[77] ^ t[78];
  assign t[63] = t[79] ^ t[80];
  assign t[64] = t[156] ^ t[157];
  assign t[65] = t[158] ^ t[159];
  assign t[66] = t[81] ^ t[69];
  assign t[67] = t[82] ^ t[50];
  assign t[68] = t[12] ? t[160] : t[83];
  assign t[69] = t[12] ? t[161] : t[84];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[85] ^ t[52];
  assign t[71] = t[86] ^ t[87];
  assign t[72] = t[88] ^ t[89];
  assign t[73] = t[90] & t[91];
  assign t[74] = t[162] ^ t[137];
  assign t[75] = t[92] ^ t[93];
  assign t[76] = t[94] & t[95];
  assign t[77] = t[95] & t[96];
  assign t[78] = t[95] ^ t[97];
  assign t[79] = t[91] & t[98];
  assign t[7] = ~(t[12]);
  assign t[80] = t[91] ^ t[97];
  assign t[81] = t[12] ? t[163] : t[99];
  assign t[82] = t[12] ? t[164] : t[100];
  assign t[83] = t[165] ^ t[166];
  assign t[84] = t[167] ^ t[168];
  assign t[85] = t[60] ^ t[86];
  assign t[86] = t[101] ^ t[82];
  assign t[87] = t[69] ^ t[60];
  assign t[88] = t[102] ^ t[93];
  assign t[89] = t[103] ^ t[70];
  assign t[8] = ~(t[13]);
  assign t[90] = t[75] ^ t[97];
  assign t[91] = t[104] ^ t[72];
  assign t[92] = t[105] ^ t[106];
  assign t[93] = t[107] ^ t[108];
  assign t[94] = t[72] ^ t[97];
  assign t[95] = t[109] ^ t[75];
  assign t[96] = t[109] & t[72];
  assign t[97] = t[104] & t[109];
  assign t[98] = t[75] & t[104];
  assign t[99] = t[169] ^ t[170];
  assign t[9] = ~(t[14] ^ t[15]);
  assign y = t[0] ? t[1] : t[135];
endmodule

module R1ind171(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind172(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind173(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind174(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind175(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind176(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind177(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind178(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind179(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind180(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind181(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind182(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind183(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind184(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind185(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind186(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind187(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind188(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind189(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind190(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind191(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind192(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind193(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind194(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind195(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind196(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind197(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind198(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind199(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind200(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind201(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind202(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind203(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind204(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind205(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind206(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind207(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind208(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind209(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind210(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind211(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind212(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind213(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind214(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind215(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind216(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind217(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind218(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind219(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind220(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind221(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind222(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind223(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind224(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind225(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind226(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind227(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind228(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind229(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind230(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind231(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind232(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind233(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind234(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind235(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind236(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind237(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind238(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind239(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind240(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind241(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind242(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind243(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind244(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind245(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind246(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind247(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind248(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind249(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind250(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind251(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind252(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind253(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind254(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind255(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind256(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind257(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind258(x, y);
 input [48:0] x;
 output y;

 wire [58:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[30]);
  assign t[12] = ~(t[30] & t[16]);
  assign t[13] = t[17] & t[18];
  assign t[14] = ~(t[31]);
  assign t[15] = ~(t[30]);
  assign t[16] = ~(t[32] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[28] : t[4];
  assign t[20] = ~(t[33] & t[34]);
  assign t[21] = ~(t[35] & t[36]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[37] & t[26]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = ~(t[40] | t[41]);
  assign t[26] = ~(t[42]);
  assign t[27] = t[43] ^ x[2];
  assign t[28] = t[44] ^ x[5];
  assign t[29] = t[45] ^ x[9];
  assign t[2] = ~(t[5]);
  assign t[30] = t[46] ^ x[12];
  assign t[31] = t[47] ^ x[15];
  assign t[32] = t[48] ^ x[18];
  assign t[33] = t[49] ^ x[21];
  assign t[34] = t[50] ^ x[24];
  assign t[35] = t[51] ^ x[27];
  assign t[36] = t[52] ^ x[30];
  assign t[37] = t[53] ^ x[33];
  assign t[38] = t[54] ^ x[36];
  assign t[39] = t[55] ^ x[39];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ^ x[42];
  assign t[41] = t[57] ^ x[45];
  assign t[42] = t[58] ^ x[48];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[7] & x[8]);
  assign t[46] = (x[10] & x[11]);
  assign t[47] = (x[13] & x[14]);
  assign t[48] = (x[16] & x[17]);
  assign t[49] = (x[19] & x[20]);
  assign t[4] = t[7] ? t[29] : x[6];
  assign t[50] = (x[22] & x[23]);
  assign t[51] = (x[25] & x[26]);
  assign t[52] = (x[28] & x[29]);
  assign t[53] = (x[31] & x[32]);
  assign t[54] = (x[34] & x[35]);
  assign t[55] = (x[37] & x[38]);
  assign t[56] = (x[40] & x[41]);
  assign t[57] = (x[43] & x[44]);
  assign t[58] = (x[46] & x[47]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = t[30] & t[13];
  assign y = t[0] ? t[1] : t[27];
endmodule

module R1ind259(x, y);
 input [60:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[44] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = ~(t[44]);
  assign t[13] = t[19] & t[20];
  assign t[14] = t[43] ^ t[41];
  assign t[15] = ~(t[44] & t[21]);
  assign t[16] = t[22] & t[23];
  assign t[17] = ~(t[45]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[42] : t[4];
  assign t[20] = ~(t[18] | t[26]);
  assign t[21] = ~(t[46] | t[27]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[47] | t[48]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[49] | t[50]);
  assign t[27] = ~(t[34] & t[35]);
  assign t[28] = ~(t[51] & t[48]);
  assign t[29] = ~(t[47] & t[52]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[50] & t[36]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[37] & t[38]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = ~(t[49]);
  assign t[37] = ~(t[58] | t[39]);
  assign t[38] = ~(t[51] | t[40]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = t[61] ^ x[2];
  assign t[42] = t[62] ^ x[5];
  assign t[43] = t[63] ^ x[9];
  assign t[44] = t[64] ^ x[12];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[18];
  assign t[47] = t[67] ^ x[21];
  assign t[48] = t[68] ^ x[24];
  assign t[49] = t[69] ^ x[27];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[30];
  assign t[51] = t[71] ^ x[33];
  assign t[52] = t[72] ^ x[36];
  assign t[53] = t[73] ^ x[39];
  assign t[54] = t[74] ^ x[42];
  assign t[55] = t[75] ^ x[45];
  assign t[56] = t[76] ^ x[48];
  assign t[57] = t[77] ^ x[51];
  assign t[58] = t[78] ^ x[54];
  assign t[59] = t[79] ^ x[57];
  assign t[5] = ~(t[9] | t[10]);
  assign t[60] = t[80] ^ x[60];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[3] & x[4]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[11]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[12]);
  assign t[80] = (x[58] & x[59]);
  assign t[8] = t[13] ? t[14] : t[43];
  assign t[9] = ~(t[15]);
  assign y = t[0] ? t[1] : t[41];
endmodule

module R1ind260(x, y);
 input [60:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[44] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = ~(t[44]);
  assign t[13] = t[19] & t[20];
  assign t[14] = t[43] ^ t[41];
  assign t[15] = ~(t[44] & t[21]);
  assign t[16] = t[22] & t[23];
  assign t[17] = ~(t[45]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[42] : t[4];
  assign t[20] = ~(t[18] | t[26]);
  assign t[21] = ~(t[46] | t[27]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[47] | t[48]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[49] | t[50]);
  assign t[27] = ~(t[34] & t[35]);
  assign t[28] = ~(t[51] & t[48]);
  assign t[29] = ~(t[47] & t[52]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[50] & t[36]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[37] & t[38]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = ~(t[49]);
  assign t[37] = ~(t[58] | t[39]);
  assign t[38] = ~(t[51] | t[40]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = t[61] ^ x[2];
  assign t[42] = t[62] ^ x[5];
  assign t[43] = t[63] ^ x[9];
  assign t[44] = t[64] ^ x[12];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[18];
  assign t[47] = t[67] ^ x[21];
  assign t[48] = t[68] ^ x[24];
  assign t[49] = t[69] ^ x[27];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[30];
  assign t[51] = t[71] ^ x[33];
  assign t[52] = t[72] ^ x[36];
  assign t[53] = t[73] ^ x[39];
  assign t[54] = t[74] ^ x[42];
  assign t[55] = t[75] ^ x[45];
  assign t[56] = t[76] ^ x[48];
  assign t[57] = t[77] ^ x[51];
  assign t[58] = t[78] ^ x[54];
  assign t[59] = t[79] ^ x[57];
  assign t[5] = ~(t[9] | t[10]);
  assign t[60] = t[80] ^ x[60];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[3] & x[4]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[11]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[12]);
  assign t[80] = (x[58] & x[59]);
  assign t[8] = t[13] ? t[14] : t[43];
  assign t[9] = ~(t[15]);
  assign y = t[0] ? t[1] : t[41];
endmodule

module R1ind261(x, y);
 input [60:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[44] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = ~(t[44]);
  assign t[13] = t[19] & t[20];
  assign t[14] = t[43] ^ t[41];
  assign t[15] = ~(t[44] & t[21]);
  assign t[16] = t[22] & t[23];
  assign t[17] = ~(t[45]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[42] : t[4];
  assign t[20] = ~(t[18] | t[26]);
  assign t[21] = ~(t[46] | t[27]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[47] | t[48]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[49] | t[50]);
  assign t[27] = ~(t[34] & t[35]);
  assign t[28] = ~(t[51] & t[48]);
  assign t[29] = ~(t[47] & t[52]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[50] & t[36]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[37] & t[38]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = ~(t[49]);
  assign t[37] = ~(t[58] | t[39]);
  assign t[38] = ~(t[51] | t[40]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = t[61] ^ x[2];
  assign t[42] = t[62] ^ x[5];
  assign t[43] = t[63] ^ x[9];
  assign t[44] = t[64] ^ x[12];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[18];
  assign t[47] = t[67] ^ x[21];
  assign t[48] = t[68] ^ x[24];
  assign t[49] = t[69] ^ x[27];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[30];
  assign t[51] = t[71] ^ x[33];
  assign t[52] = t[72] ^ x[36];
  assign t[53] = t[73] ^ x[39];
  assign t[54] = t[74] ^ x[42];
  assign t[55] = t[75] ^ x[45];
  assign t[56] = t[76] ^ x[48];
  assign t[57] = t[77] ^ x[51];
  assign t[58] = t[78] ^ x[54];
  assign t[59] = t[79] ^ x[57];
  assign t[5] = ~(t[9] | t[10]);
  assign t[60] = t[80] ^ x[60];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[3] & x[4]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[11]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[12]);
  assign t[80] = (x[58] & x[59]);
  assign t[8] = t[13] ? t[14] : t[43];
  assign t[9] = ~(t[15]);
  assign y = t[0] ? t[1] : t[41];
endmodule

module R1ind262(x, y);
 input [60:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[44] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = ~(t[44]);
  assign t[13] = t[19] & t[20];
  assign t[14] = t[43] ^ t[41];
  assign t[15] = ~(t[44] & t[21]);
  assign t[16] = t[22] & t[23];
  assign t[17] = ~(t[45]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[42] : t[4];
  assign t[20] = ~(t[18] | t[26]);
  assign t[21] = ~(t[46] | t[27]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[47] | t[48]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[49] | t[50]);
  assign t[27] = ~(t[34] & t[35]);
  assign t[28] = ~(t[51] & t[48]);
  assign t[29] = ~(t[47] & t[52]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[50] & t[36]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[37] & t[38]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = ~(t[49]);
  assign t[37] = ~(t[58] | t[39]);
  assign t[38] = ~(t[51] | t[40]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = t[61] ^ x[2];
  assign t[42] = t[62] ^ x[5];
  assign t[43] = t[63] ^ x[9];
  assign t[44] = t[64] ^ x[12];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[18];
  assign t[47] = t[67] ^ x[21];
  assign t[48] = t[68] ^ x[24];
  assign t[49] = t[69] ^ x[27];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[30];
  assign t[51] = t[71] ^ x[33];
  assign t[52] = t[72] ^ x[36];
  assign t[53] = t[73] ^ x[39];
  assign t[54] = t[74] ^ x[42];
  assign t[55] = t[75] ^ x[45];
  assign t[56] = t[76] ^ x[48];
  assign t[57] = t[77] ^ x[51];
  assign t[58] = t[78] ^ x[54];
  assign t[59] = t[79] ^ x[57];
  assign t[5] = ~(t[9] | t[10]);
  assign t[60] = t[80] ^ x[60];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[3] & x[4]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[11]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[12]);
  assign t[80] = (x[58] & x[59]);
  assign t[8] = t[13] ? t[14] : t[43];
  assign t[9] = ~(t[15]);
  assign y = t[0] ? t[1] : t[41];
endmodule

module R1ind263(x, y);
 input [60:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[44] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = ~(t[44]);
  assign t[13] = t[19] & t[20];
  assign t[14] = t[43] ^ t[41];
  assign t[15] = ~(t[44] & t[21]);
  assign t[16] = t[22] & t[23];
  assign t[17] = ~(t[45]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[42] : t[4];
  assign t[20] = ~(t[18] | t[26]);
  assign t[21] = ~(t[46] | t[27]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[47] | t[48]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[49] | t[50]);
  assign t[27] = ~(t[34] & t[35]);
  assign t[28] = ~(t[51] & t[48]);
  assign t[29] = ~(t[47] & t[52]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[50] & t[36]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[37] & t[38]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = ~(t[49]);
  assign t[37] = ~(t[58] | t[39]);
  assign t[38] = ~(t[51] | t[40]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = t[61] ^ x[2];
  assign t[42] = t[62] ^ x[5];
  assign t[43] = t[63] ^ x[9];
  assign t[44] = t[64] ^ x[12];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[18];
  assign t[47] = t[67] ^ x[21];
  assign t[48] = t[68] ^ x[24];
  assign t[49] = t[69] ^ x[27];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[30];
  assign t[51] = t[71] ^ x[33];
  assign t[52] = t[72] ^ x[36];
  assign t[53] = t[73] ^ x[39];
  assign t[54] = t[74] ^ x[42];
  assign t[55] = t[75] ^ x[45];
  assign t[56] = t[76] ^ x[48];
  assign t[57] = t[77] ^ x[51];
  assign t[58] = t[78] ^ x[54];
  assign t[59] = t[79] ^ x[57];
  assign t[5] = ~(t[9] | t[10]);
  assign t[60] = t[80] ^ x[60];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[3] & x[4]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[11]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[12]);
  assign t[80] = (x[58] & x[59]);
  assign t[8] = t[13] ? t[14] : t[43];
  assign t[9] = ~(t[15]);
  assign y = t[0] ? t[1] : t[41];
endmodule

module R1ind264(x, y);
 input [60:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[44] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = ~(t[44]);
  assign t[13] = t[19] & t[20];
  assign t[14] = t[43] ^ t[41];
  assign t[15] = ~(t[44] & t[21]);
  assign t[16] = t[22] & t[23];
  assign t[17] = ~(t[45]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[42] : t[4];
  assign t[20] = ~(t[18] | t[26]);
  assign t[21] = ~(t[46] | t[27]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[47] | t[48]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[49] | t[50]);
  assign t[27] = ~(t[34] & t[35]);
  assign t[28] = ~(t[51] & t[48]);
  assign t[29] = ~(t[47] & t[52]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[50] & t[36]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[37] & t[38]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = ~(t[49]);
  assign t[37] = ~(t[58] | t[39]);
  assign t[38] = ~(t[51] | t[40]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = t[61] ^ x[2];
  assign t[42] = t[62] ^ x[5];
  assign t[43] = t[63] ^ x[9];
  assign t[44] = t[64] ^ x[12];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[18];
  assign t[47] = t[67] ^ x[21];
  assign t[48] = t[68] ^ x[24];
  assign t[49] = t[69] ^ x[27];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[30];
  assign t[51] = t[71] ^ x[33];
  assign t[52] = t[72] ^ x[36];
  assign t[53] = t[73] ^ x[39];
  assign t[54] = t[74] ^ x[42];
  assign t[55] = t[75] ^ x[45];
  assign t[56] = t[76] ^ x[48];
  assign t[57] = t[77] ^ x[51];
  assign t[58] = t[78] ^ x[54];
  assign t[59] = t[79] ^ x[57];
  assign t[5] = ~(t[9] | t[10]);
  assign t[60] = t[80] ^ x[60];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[3] & x[4]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[11]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[12]);
  assign t[80] = (x[58] & x[59]);
  assign t[8] = t[13] ? t[14] : t[43];
  assign t[9] = ~(t[15]);
  assign y = t[0] ? t[1] : t[41];
endmodule

module R1ind265(x, y);
 input [60:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[44] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = ~(t[44]);
  assign t[13] = t[19] & t[20];
  assign t[14] = t[43] ^ t[41];
  assign t[15] = ~(t[44] & t[21]);
  assign t[16] = t[22] & t[23];
  assign t[17] = ~(t[45]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[42] : t[4];
  assign t[20] = ~(t[18] | t[26]);
  assign t[21] = ~(t[46] | t[27]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[47] | t[48]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[49] | t[50]);
  assign t[27] = ~(t[34] & t[35]);
  assign t[28] = ~(t[51] & t[48]);
  assign t[29] = ~(t[47] & t[52]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[50] & t[36]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[37] & t[38]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = ~(t[49]);
  assign t[37] = ~(t[58] | t[39]);
  assign t[38] = ~(t[51] | t[40]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = t[61] ^ x[2];
  assign t[42] = t[62] ^ x[5];
  assign t[43] = t[63] ^ x[9];
  assign t[44] = t[64] ^ x[12];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[18];
  assign t[47] = t[67] ^ x[21];
  assign t[48] = t[68] ^ x[24];
  assign t[49] = t[69] ^ x[27];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[30];
  assign t[51] = t[71] ^ x[33];
  assign t[52] = t[72] ^ x[36];
  assign t[53] = t[73] ^ x[39];
  assign t[54] = t[74] ^ x[42];
  assign t[55] = t[75] ^ x[45];
  assign t[56] = t[76] ^ x[48];
  assign t[57] = t[77] ^ x[51];
  assign t[58] = t[78] ^ x[54];
  assign t[59] = t[79] ^ x[57];
  assign t[5] = ~(t[9] | t[10]);
  assign t[60] = t[80] ^ x[60];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[3] & x[4]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[11]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[12]);
  assign t[80] = (x[58] & x[59]);
  assign t[8] = t[13] ? t[14] : t[43];
  assign t[9] = ~(t[15]);
  assign y = t[0] ? t[1] : t[41];
endmodule

module R1ind266(x, y);
 input [60:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[44] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = ~(t[44]);
  assign t[13] = t[19] & t[20];
  assign t[14] = t[43] ^ t[41];
  assign t[15] = ~(t[44] & t[21]);
  assign t[16] = t[22] & t[23];
  assign t[17] = ~(t[45]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = t[3] ? t[42] : t[4];
  assign t[20] = ~(t[18] | t[26]);
  assign t[21] = ~(t[46] | t[27]);
  assign t[22] = ~(t[28] | t[29]);
  assign t[23] = ~(t[30] | t[31]);
  assign t[24] = ~(t[47] | t[48]);
  assign t[25] = ~(t[32] | t[33]);
  assign t[26] = ~(t[49] | t[50]);
  assign t[27] = ~(t[34] & t[35]);
  assign t[28] = ~(t[51] & t[48]);
  assign t[29] = ~(t[47] & t[52]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[21]);
  assign t[31] = ~(t[50] & t[36]);
  assign t[32] = ~(t[52] & t[53]);
  assign t[33] = ~(t[37] & t[38]);
  assign t[34] = ~(t[54] | t[55]);
  assign t[35] = ~(t[56] | t[57]);
  assign t[36] = ~(t[49]);
  assign t[37] = ~(t[58] | t[39]);
  assign t[38] = ~(t[51] | t[40]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = t[61] ^ x[2];
  assign t[42] = t[62] ^ x[5];
  assign t[43] = t[63] ^ x[9];
  assign t[44] = t[64] ^ x[12];
  assign t[45] = t[65] ^ x[15];
  assign t[46] = t[66] ^ x[18];
  assign t[47] = t[67] ^ x[21];
  assign t[48] = t[68] ^ x[24];
  assign t[49] = t[69] ^ x[27];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[30];
  assign t[51] = t[71] ^ x[33];
  assign t[52] = t[72] ^ x[36];
  assign t[53] = t[73] ^ x[39];
  assign t[54] = t[74] ^ x[42];
  assign t[55] = t[75] ^ x[45];
  assign t[56] = t[76] ^ x[48];
  assign t[57] = t[77] ^ x[51];
  assign t[58] = t[78] ^ x[54];
  assign t[59] = t[79] ^ x[57];
  assign t[5] = ~(t[9] | t[10]);
  assign t[60] = t[80] ^ x[60];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[3] & x[4]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[11]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[12]);
  assign t[80] = (x[58] & x[59]);
  assign t[8] = t[13] ? t[14] : t[43];
  assign t[9] = ~(t[15]);
  assign y = t[0] ? t[1] : t[41];
endmodule

module R1ind267(x, y);
 input [129:0] x;
 output y;

 wire [224:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[78] ^ t[103];
  assign t[101] = t[119] ^ t[80];
  assign t[102] = t[115] & t[80];
  assign t[103] = t[119] & t[115];
  assign t[104] = t[78] & t[119];
  assign t[105] = t[173] ^ t[174];
  assign t[106] = t[175] ^ t[176];
  assign t[107] = t[177] ^ t[178];
  assign t[108] = t[179] ^ t[180];
  assign t[109] = t[87] ^ t[89];
  assign t[10] = ~(t[16]);
  assign t[110] = t[155] ^ t[181];
  assign t[111] = t[120] ^ t[121];
  assign t[112] = t[91] ^ t[122];
  assign t[113] = t[91] & t[122];
  assign t[114] = t[58] & t[63];
  assign t[115] = t[123] ^ t[124];
  assign t[116] = t[125] ^ t[126];
  assign t[117] = t[58] ^ t[127];
  assign t[118] = t[75] ^ t[57];
  assign t[119] = t[128] ^ t[124];
  assign t[11] = ~(t[141]);
  assign t[120] = t[127] & t[89];
  assign t[121] = t[60] & t[129];
  assign t[122] = t[129] ^ t[90];
  assign t[123] = t[130] ^ t[131];
  assign t[124] = t[132] ^ t[114];
  assign t[125] = t[117] & t[118];
  assign t[126] = t[74] & t[57];
  assign t[127] = t[90] ^ t[133];
  assign t[128] = t[134] ^ t[135];
  assign t[129] = t[58] ^ t[71];
  assign t[12] = ~(t[17]);
  assign t[130] = t[136] ^ t[121];
  assign t[131] = t[76] & t[137];
  assign t[132] = t[45] & t[64];
  assign t[133] = t[54] ^ t[89];
  assign t[134] = t[138] ^ t[126];
  assign t[135] = t[92] & t[75];
  assign t[136] = t[129] ^ t[77];
  assign t[137] = t[89] ^ t[129];
  assign t[138] = t[74] ^ t[57];
  assign t[139] = t[182] ^ x[2];
  assign t[13] = t[18] ? t[20] : t[19];
  assign t[140] = t[183] ^ x[5];
  assign t[141] = t[184] ^ x[9];
  assign t[142] = t[185] ^ x[12];
  assign t[143] = t[186] ^ x[15];
  assign t[144] = t[187] ^ x[18];
  assign t[145] = t[188] ^ x[21];
  assign t[146] = t[189] ^ x[24];
  assign t[147] = t[190] ^ x[27];
  assign t[148] = t[191] ^ x[30];
  assign t[149] = t[192] ^ x[33];
  assign t[14] = t[18] ? t[142] : t[21];
  assign t[150] = t[193] ^ x[36];
  assign t[151] = t[194] ^ x[39];
  assign t[152] = t[195] ^ x[42];
  assign t[153] = t[196] ^ x[45];
  assign t[154] = t[197] ^ x[48];
  assign t[155] = t[198] ^ x[51];
  assign t[156] = t[199] ^ x[54];
  assign t[157] = t[200] ^ x[57];
  assign t[158] = t[201] ^ x[60];
  assign t[159] = t[202] ^ x[63];
  assign t[15] = t[18] & t[22];
  assign t[160] = t[203] ^ x[66];
  assign t[161] = t[204] ^ x[69];
  assign t[162] = t[205] ^ x[72];
  assign t[163] = t[206] ^ x[75];
  assign t[164] = t[207] ^ x[78];
  assign t[165] = t[208] ^ x[81];
  assign t[166] = t[209] ^ x[84];
  assign t[167] = t[210] ^ x[87];
  assign t[168] = t[211] ^ x[90];
  assign t[169] = t[212] ^ x[93];
  assign t[16] = ~(t[141] & t[23]);
  assign t[170] = t[213] ^ x[96];
  assign t[171] = t[214] ^ x[99];
  assign t[172] = t[215] ^ x[102];
  assign t[173] = t[216] ^ x[105];
  assign t[174] = t[217] ^ x[108];
  assign t[175] = t[218] ^ x[111];
  assign t[176] = t[219] ^ x[114];
  assign t[177] = t[220] ^ x[117];
  assign t[178] = t[221] ^ x[120];
  assign t[179] = t[222] ^ x[123];
  assign t[17] = ~(t[24]);
  assign t[180] = t[223] ^ x[126];
  assign t[181] = t[224] ^ x[129];
  assign t[182] = (x[0] & x[1]);
  assign t[183] = (x[3] & x[4]);
  assign t[184] = (x[7] & x[8]);
  assign t[185] = (x[10] & x[11]);
  assign t[186] = (x[13] & x[14]);
  assign t[187] = (x[16] & x[17]);
  assign t[188] = (x[19] & x[20]);
  assign t[189] = (x[22] & x[23]);
  assign t[18] = ~(t[25] | t[26]);
  assign t[190] = (x[25] & x[26]);
  assign t[191] = (x[28] & x[29]);
  assign t[192] = (x[31] & x[32]);
  assign t[193] = (x[34] & x[35]);
  assign t[194] = (x[37] & x[38]);
  assign t[195] = (x[40] & x[41]);
  assign t[196] = (x[43] & x[44]);
  assign t[197] = (x[46] & x[47]);
  assign t[198] = (x[49] & x[50]);
  assign t[199] = (x[52] & x[53]);
  assign t[19] = t[27] ^ t[28];
  assign t[1] = t[3] ? t[140] : t[4];
  assign t[200] = (x[55] & x[56]);
  assign t[201] = (x[58] & x[59]);
  assign t[202] = (x[61] & x[62]);
  assign t[203] = (x[64] & x[65]);
  assign t[204] = (x[67] & x[68]);
  assign t[205] = (x[70] & x[71]);
  assign t[206] = (x[73] & x[74]);
  assign t[207] = (x[76] & x[77]);
  assign t[208] = (x[79] & x[80]);
  assign t[209] = (x[82] & x[83]);
  assign t[20] = t[143] ^ t[144];
  assign t[210] = (x[85] & x[86]);
  assign t[211] = (x[88] & x[89]);
  assign t[212] = (x[91] & x[92]);
  assign t[213] = (x[94] & x[95]);
  assign t[214] = (x[97] & x[98]);
  assign t[215] = (x[100] & x[101]);
  assign t[216] = (x[103] & x[104]);
  assign t[217] = (x[106] & x[107]);
  assign t[218] = (x[109] & x[110]);
  assign t[219] = (x[112] & x[113]);
  assign t[21] = ~(t[29] ^ t[30]);
  assign t[220] = (x[115] & x[116]);
  assign t[221] = (x[118] & x[119]);
  assign t[222] = (x[121] & x[122]);
  assign t[223] = (x[124] & x[125]);
  assign t[224] = (x[127] & x[128]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[145] | t[33]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[25] = ~(t[146] & t[147]);
  assign t[26] = ~(t[148] & t[149]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[150] ^ t[40];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[151] ^ t[152]);
  assign t[31] = ~(t[23]);
  assign t[32] = ~(t[153] & t[41]);
  assign t[33] = ~(t[42] & t[43]);
  assign t[34] = ~(t[154]);
  assign t[35] = ~(t[141]);
  assign t[36] = t[44] & t[45];
  assign t[37] = t[46] ^ t[47];
  assign t[38] = t[48] ^ t[49];
  assign t[39] = t[50] ^ t[51];
  assign t[3] = ~(t[6]);
  assign t[40] = t[143] ^ t[155];
  assign t[41] = ~(t[156]);
  assign t[42] = ~(t[157] | t[158]);
  assign t[43] = ~(t[159] | t[160]);
  assign t[44] = t[52] ^ t[53];
  assign t[45] = t[54] ^ t[55];
  assign t[46] = t[56] & t[57];
  assign t[47] = t[52] & t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[61] ^ t[62];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[52] & t[63];
  assign t[51] = t[44] & t[64];
  assign t[52] = t[65] ^ t[66];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[24] ? t[161] : t[69];
  assign t[55] = t[24] ? t[162] : t[70];
  assign t[56] = t[65] ^ t[67];
  assign t[57] = t[71] ^ t[72];
  assign t[58] = t[73] ^ t[54];
  assign t[59] = t[66] ^ t[68];
  assign t[5] = ~(t[9]);
  assign t[60] = t[74] ^ t[45];
  assign t[61] = t[67] & t[75];
  assign t[62] = t[68] & t[76];
  assign t[63] = t[71] ^ t[77];
  assign t[64] = t[58] ^ t[72];
  assign t[65] = t[78] ^ t[79];
  assign t[66] = t[80] ^ t[81];
  assign t[67] = t[82] ^ t[83];
  assign t[68] = t[84] ^ t[85];
  assign t[69] = t[163] ^ t[164];
  assign t[6] = ~(t[10]);
  assign t[70] = t[165] ^ t[166];
  assign t[71] = t[86] ^ t[87];
  assign t[72] = t[88] ^ t[55];
  assign t[73] = t[24] ? t[167] : t[20];
  assign t[74] = t[73] ^ t[87];
  assign t[75] = t[89] ^ t[90];
  assign t[76] = t[91] ^ t[92];
  assign t[77] = t[93] ^ t[55];
  assign t[78] = t[94] ^ t[95];
  assign t[79] = t[96] & t[97];
  assign t[7] = ~(t[11]);
  assign t[80] = t[98] ^ t[99];
  assign t[81] = t[100] & t[101];
  assign t[82] = t[97] & t[102];
  assign t[83] = t[97] ^ t[103];
  assign t[84] = t[101] & t[104];
  assign t[85] = t[101] ^ t[103];
  assign t[86] = t[24] ? t[168] : t[105];
  assign t[87] = t[24] ? t[169] : t[106];
  assign t[88] = t[24] ? t[170] : t[107];
  assign t[89] = t[24] ? t[171] : t[108];
  assign t[8] = t[12] ? t[14] : t[13];
  assign t[90] = t[93] ^ t[88];
  assign t[91] = t[73] ^ t[55];
  assign t[92] = t[90] ^ t[109];
  assign t[93] = t[24] ? t[172] : t[110];
  assign t[94] = t[111] ^ t[112];
  assign t[95] = t[113] ^ t[114];
  assign t[96] = t[80] ^ t[103];
  assign t[97] = t[115] ^ t[78];
  assign t[98] = t[116] ^ t[95];
  assign t[99] = t[117] ^ t[118];
  assign t[9] = t[141] & t[15];
  assign y = t[0] ? t[1] : t[139];
endmodule

module R1ind268(x, y);
 input [129:0] x;
 output y;

 wire [223:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[118] ^ t[103];
  assign t[101] = t[119] ^ t[120];
  assign t[102] = t[121] ^ t[122];
  assign t[103] = t[123] ^ t[117];
  assign t[104] = t[124] ^ t[125];
  assign t[105] = t[154] ^ t[174];
  assign t[106] = t[175] ^ t[176];
  assign t[107] = t[177] ^ t[178];
  assign t[108] = t[83] ^ t[68];
  assign t[109] = t[85] ^ t[84];
  assign t[10] = ~(t[16]);
  assign t[110] = t[84] ^ t[68];
  assign t[111] = t[109] & t[126];
  assign t[112] = t[109] ^ t[68];
  assign t[113] = t[179] ^ t[180];
  assign t[114] = t[127] ^ t[128];
  assign t[115] = t[55] & t[129];
  assign t[116] = t[59] & t[65];
  assign t[117] = t[57] & t[64];
  assign t[118] = t[130] ^ t[128];
  assign t[119] = t[57] ^ t[131];
  assign t[11] = ~(t[140]);
  assign t[120] = t[129] ^ t[132];
  assign t[121] = t[133] ^ t[134];
  assign t[122] = t[54] ^ t[135];
  assign t[123] = t[54] & t[135];
  assign t[124] = t[136] ^ t[134];
  assign t[125] = t[45] & t[78];
  assign t[126] = t[85] & t[83];
  assign t[127] = t[97] ^ t[132];
  assign t[128] = t[97] & t[132];
  assign t[129] = t[91] ^ t[71];
  assign t[12] = ~(t[17]);
  assign t[130] = t[119] & t[120];
  assign t[131] = t[71] ^ t[137];
  assign t[132] = t[77] ^ t[81];
  assign t[133] = t[131] & t[91];
  assign t[134] = t[79] & t[61];
  assign t[135] = t[61] ^ t[71];
  assign t[136] = t[61] ^ t[80];
  assign t[137] = t[75] ^ t[91];
  assign t[138] = t[181] ^ x[2];
  assign t[139] = t[182] ^ x[5];
  assign t[13] = t[18] ? t[20] : t[19];
  assign t[140] = t[183] ^ x[9];
  assign t[141] = t[184] ^ x[12];
  assign t[142] = t[185] ^ x[15];
  assign t[143] = t[186] ^ x[18];
  assign t[144] = t[187] ^ x[21];
  assign t[145] = t[188] ^ x[24];
  assign t[146] = t[189] ^ x[27];
  assign t[147] = t[190] ^ x[30];
  assign t[148] = t[191] ^ x[33];
  assign t[149] = t[192] ^ x[36];
  assign t[14] = t[18] ? t[141] : t[21];
  assign t[150] = t[193] ^ x[39];
  assign t[151] = t[194] ^ x[42];
  assign t[152] = t[195] ^ x[45];
  assign t[153] = t[196] ^ x[48];
  assign t[154] = t[197] ^ x[51];
  assign t[155] = t[198] ^ x[54];
  assign t[156] = t[199] ^ x[57];
  assign t[157] = t[200] ^ x[60];
  assign t[158] = t[201] ^ x[63];
  assign t[159] = t[202] ^ x[66];
  assign t[15] = t[18] & t[22];
  assign t[160] = t[203] ^ x[69];
  assign t[161] = t[204] ^ x[72];
  assign t[162] = t[205] ^ x[75];
  assign t[163] = t[206] ^ x[78];
  assign t[164] = t[207] ^ x[81];
  assign t[165] = t[208] ^ x[84];
  assign t[166] = t[209] ^ x[87];
  assign t[167] = t[210] ^ x[90];
  assign t[168] = t[211] ^ x[93];
  assign t[169] = t[212] ^ x[96];
  assign t[16] = ~(t[140] & t[23]);
  assign t[170] = t[213] ^ x[99];
  assign t[171] = t[214] ^ x[102];
  assign t[172] = t[215] ^ x[105];
  assign t[173] = t[216] ^ x[108];
  assign t[174] = t[217] ^ x[111];
  assign t[175] = t[218] ^ x[114];
  assign t[176] = t[219] ^ x[117];
  assign t[177] = t[220] ^ x[120];
  assign t[178] = t[221] ^ x[123];
  assign t[179] = t[222] ^ x[126];
  assign t[17] = ~(t[24]);
  assign t[180] = t[223] ^ x[129];
  assign t[181] = (x[0] & x[1]);
  assign t[182] = (x[3] & x[4]);
  assign t[183] = (x[7] & x[8]);
  assign t[184] = (x[10] & x[11]);
  assign t[185] = (x[13] & x[14]);
  assign t[186] = (x[16] & x[17]);
  assign t[187] = (x[19] & x[20]);
  assign t[188] = (x[22] & x[23]);
  assign t[189] = (x[25] & x[26]);
  assign t[18] = ~(t[25] | t[26]);
  assign t[190] = (x[28] & x[29]);
  assign t[191] = (x[31] & x[32]);
  assign t[192] = (x[34] & x[35]);
  assign t[193] = (x[37] & x[38]);
  assign t[194] = (x[40] & x[41]);
  assign t[195] = (x[43] & x[44]);
  assign t[196] = (x[46] & x[47]);
  assign t[197] = (x[49] & x[50]);
  assign t[198] = (x[52] & x[53]);
  assign t[199] = (x[55] & x[56]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = t[3] ? t[139] : t[4];
  assign t[200] = (x[58] & x[59]);
  assign t[201] = (x[61] & x[62]);
  assign t[202] = (x[64] & x[65]);
  assign t[203] = (x[67] & x[68]);
  assign t[204] = (x[70] & x[71]);
  assign t[205] = (x[73] & x[74]);
  assign t[206] = (x[76] & x[77]);
  assign t[207] = (x[79] & x[80]);
  assign t[208] = (x[82] & x[83]);
  assign t[209] = (x[85] & x[86]);
  assign t[20] = t[142] ^ t[143];
  assign t[210] = (x[88] & x[89]);
  assign t[211] = (x[91] & x[92]);
  assign t[212] = (x[94] & x[95]);
  assign t[213] = (x[97] & x[98]);
  assign t[214] = (x[100] & x[101]);
  assign t[215] = (x[103] & x[104]);
  assign t[216] = (x[106] & x[107]);
  assign t[217] = (x[109] & x[110]);
  assign t[218] = (x[112] & x[113]);
  assign t[219] = (x[115] & x[116]);
  assign t[21] = ~(t[29] ^ t[30]);
  assign t[220] = (x[118] & x[119]);
  assign t[221] = (x[121] & x[122]);
  assign t[222] = (x[124] & x[125]);
  assign t[223] = (x[127] & x[128]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[144] | t[33]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[25] = ~(t[145] & t[146]);
  assign t[26] = ~(t[147] & t[148]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[149] ^ t[40];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[150] ^ t[151]);
  assign t[31] = ~(t[23]);
  assign t[32] = ~(t[152] & t[41]);
  assign t[33] = ~(t[42] & t[43]);
  assign t[34] = ~(t[153]);
  assign t[35] = ~(t[140]);
  assign t[36] = t[44] & t[45];
  assign t[37] = t[46] ^ t[47];
  assign t[38] = t[48] ^ t[49];
  assign t[39] = t[50] ^ t[51];
  assign t[3] = ~(t[6]);
  assign t[40] = t[142] ^ t[154];
  assign t[41] = ~(t[155]);
  assign t[42] = ~(t[156] | t[157]);
  assign t[43] = ~(t[158] | t[159]);
  assign t[44] = t[52] ^ t[53];
  assign t[45] = t[54] ^ t[55];
  assign t[46] = t[56] & t[57];
  assign t[47] = t[58] & t[59];
  assign t[48] = t[60] & t[61];
  assign t[49] = t[62] ^ t[63];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[56] & t[64];
  assign t[51] = t[58] & t[65];
  assign t[52] = t[66] & t[67];
  assign t[53] = t[66] ^ t[68];
  assign t[54] = t[69] ^ t[70];
  assign t[55] = t[71] ^ t[72];
  assign t[56] = t[73] ^ t[74];
  assign t[57] = t[69] ^ t[75];
  assign t[58] = t[56] ^ t[76];
  assign t[59] = t[75] ^ t[70];
  assign t[5] = ~(t[9]);
  assign t[60] = t[74] ^ t[44];
  assign t[61] = t[57] ^ t[77];
  assign t[62] = t[44] & t[78];
  assign t[63] = t[60] & t[79];
  assign t[64] = t[77] ^ t[80];
  assign t[65] = t[57] ^ t[81];
  assign t[66] = t[82] ^ t[83];
  assign t[67] = t[84] & t[82];
  assign t[68] = t[82] & t[85];
  assign t[69] = t[24] ? t[160] : t[86];
  assign t[6] = ~(t[10]);
  assign t[70] = t[24] ? t[161] : t[87];
  assign t[71] = t[88] ^ t[89];
  assign t[72] = t[90] ^ t[91];
  assign t[73] = t[84] ^ t[92];
  assign t[74] = t[83] ^ t[93];
  assign t[75] = t[24] ? t[162] : t[94];
  assign t[76] = t[95] ^ t[44];
  assign t[77] = t[96] ^ t[90];
  assign t[78] = t[91] ^ t[61];
  assign t[79] = t[97] ^ t[59];
  assign t[7] = ~(t[11]);
  assign t[80] = t[88] ^ t[70];
  assign t[81] = t[89] ^ t[70];
  assign t[82] = t[98] ^ t[99];
  assign t[83] = t[100] ^ t[101];
  assign t[84] = t[102] ^ t[103];
  assign t[85] = t[104] ^ t[99];
  assign t[86] = t[163] ^ t[164];
  assign t[87] = t[165] ^ t[166];
  assign t[88] = t[24] ? t[167] : t[20];
  assign t[89] = t[24] ? t[168] : t[105];
  assign t[8] = t[12] ? t[14] : t[13];
  assign t[90] = t[24] ? t[169] : t[106];
  assign t[91] = t[24] ? t[170] : t[107];
  assign t[92] = t[108] & t[109];
  assign t[93] = t[110] & t[66];
  assign t[94] = t[171] ^ t[172];
  assign t[95] = t[111] ^ t[112];
  assign t[96] = t[24] ? t[173] : t[113];
  assign t[97] = t[69] ^ t[90];
  assign t[98] = t[114] ^ t[115];
  assign t[99] = t[116] ^ t[117];
  assign t[9] = t[140] & t[15];
  assign y = t[0] ? t[1] : t[138];
endmodule

module R1ind269(x, y);
 input [129:0] x;
 output y;

 wire [223:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[154] ^ t[176];
  assign t[101] = t[112] ^ t[113];
  assign t[102] = t[114] ^ t[113];
  assign t[103] = t[177] ^ t[178];
  assign t[104] = t[115] ^ t[116];
  assign t[105] = t[45] ^ t[56];
  assign t[106] = t[45] & t[56];
  assign t[107] = t[65] & t[64];
  assign t[108] = t[117] ^ t[93];
  assign t[109] = t[60] ^ t[118];
  assign t[10] = ~(t[16]);
  assign t[110] = t[75] ^ t[86];
  assign t[111] = t[179] ^ t[180];
  assign t[112] = t[119] ^ t[120];
  assign t[113] = t[121] ^ t[107];
  assign t[114] = t[122] ^ t[123];
  assign t[115] = t[77] & t[80];
  assign t[116] = t[124] & t[72];
  assign t[117] = t[125] ^ t[126];
  assign t[118] = t[127] ^ t[128];
  assign t[119] = t[129] ^ t[116];
  assign t[11] = ~(t[140]);
  assign t[120] = t[130] & t[131];
  assign t[121] = t[132] & t[133];
  assign t[122] = t[134] ^ t[126];
  assign t[123] = t[135] & t[127];
  assign t[124] = t[58] ^ t[132];
  assign t[125] = t[60] & t[118];
  assign t[126] = t[58] & t[128];
  assign t[127] = t[80] ^ t[73];
  assign t[128] = t[81] ^ t[136];
  assign t[129] = t[72] ^ t[82];
  assign t[12] = ~(t[17]);
  assign t[130] = t[45] ^ t[135];
  assign t[131] = t[80] ^ t[72];
  assign t[132] = t[83] ^ t[55];
  assign t[133] = t[65] ^ t[136];
  assign t[134] = t[58] ^ t[128];
  assign t[135] = t[73] ^ t[137];
  assign t[136] = t[90] ^ t[55];
  assign t[137] = t[74] ^ t[80];
  assign t[138] = t[181] ^ x[2];
  assign t[139] = t[182] ^ x[5];
  assign t[13] = t[18] ? t[20] : t[19];
  assign t[140] = t[183] ^ x[9];
  assign t[141] = t[184] ^ x[12];
  assign t[142] = t[185] ^ x[15];
  assign t[143] = t[186] ^ x[18];
  assign t[144] = t[187] ^ x[21];
  assign t[145] = t[188] ^ x[24];
  assign t[146] = t[189] ^ x[27];
  assign t[147] = t[190] ^ x[30];
  assign t[148] = t[191] ^ x[33];
  assign t[149] = t[192] ^ x[36];
  assign t[14] = t[18] ? t[141] : t[21];
  assign t[150] = t[193] ^ x[39];
  assign t[151] = t[194] ^ x[42];
  assign t[152] = t[195] ^ x[45];
  assign t[153] = t[196] ^ x[48];
  assign t[154] = t[197] ^ x[51];
  assign t[155] = t[198] ^ x[54];
  assign t[156] = t[199] ^ x[57];
  assign t[157] = t[200] ^ x[60];
  assign t[158] = t[201] ^ x[63];
  assign t[159] = t[202] ^ x[66];
  assign t[15] = t[18] & t[22];
  assign t[160] = t[203] ^ x[69];
  assign t[161] = t[204] ^ x[72];
  assign t[162] = t[205] ^ x[75];
  assign t[163] = t[206] ^ x[78];
  assign t[164] = t[207] ^ x[81];
  assign t[165] = t[208] ^ x[84];
  assign t[166] = t[209] ^ x[87];
  assign t[167] = t[210] ^ x[90];
  assign t[168] = t[211] ^ x[93];
  assign t[169] = t[212] ^ x[96];
  assign t[16] = ~(t[140] & t[23]);
  assign t[170] = t[213] ^ x[99];
  assign t[171] = t[214] ^ x[102];
  assign t[172] = t[215] ^ x[105];
  assign t[173] = t[216] ^ x[108];
  assign t[174] = t[217] ^ x[111];
  assign t[175] = t[218] ^ x[114];
  assign t[176] = t[219] ^ x[117];
  assign t[177] = t[220] ^ x[120];
  assign t[178] = t[221] ^ x[123];
  assign t[179] = t[222] ^ x[126];
  assign t[17] = ~(t[24]);
  assign t[180] = t[223] ^ x[129];
  assign t[181] = (x[0] & x[1]);
  assign t[182] = (x[3] & x[4]);
  assign t[183] = (x[7] & x[8]);
  assign t[184] = (x[10] & x[11]);
  assign t[185] = (x[13] & x[14]);
  assign t[186] = (x[16] & x[17]);
  assign t[187] = (x[19] & x[20]);
  assign t[188] = (x[22] & x[23]);
  assign t[189] = (x[25] & x[26]);
  assign t[18] = ~(t[25] | t[26]);
  assign t[190] = (x[28] & x[29]);
  assign t[191] = (x[31] & x[32]);
  assign t[192] = (x[34] & x[35]);
  assign t[193] = (x[37] & x[38]);
  assign t[194] = (x[40] & x[41]);
  assign t[195] = (x[43] & x[44]);
  assign t[196] = (x[46] & x[47]);
  assign t[197] = (x[49] & x[50]);
  assign t[198] = (x[52] & x[53]);
  assign t[199] = (x[55] & x[56]);
  assign t[19] = ~(t[27] ^ t[28]);
  assign t[1] = t[3] ? t[139] : t[4];
  assign t[200] = (x[58] & x[59]);
  assign t[201] = (x[61] & x[62]);
  assign t[202] = (x[64] & x[65]);
  assign t[203] = (x[67] & x[68]);
  assign t[204] = (x[70] & x[71]);
  assign t[205] = (x[73] & x[74]);
  assign t[206] = (x[76] & x[77]);
  assign t[207] = (x[79] & x[80]);
  assign t[208] = (x[82] & x[83]);
  assign t[209] = (x[85] & x[86]);
  assign t[20] = t[142] ^ t[143];
  assign t[210] = (x[88] & x[89]);
  assign t[211] = (x[91] & x[92]);
  assign t[212] = (x[94] & x[95]);
  assign t[213] = (x[97] & x[98]);
  assign t[214] = (x[100] & x[101]);
  assign t[215] = (x[103] & x[104]);
  assign t[216] = (x[106] & x[107]);
  assign t[217] = (x[109] & x[110]);
  assign t[218] = (x[112] & x[113]);
  assign t[219] = (x[115] & x[116]);
  assign t[21] = ~(t[29] ^ t[30]);
  assign t[220] = (x[118] & x[119]);
  assign t[221] = (x[121] & x[122]);
  assign t[222] = (x[124] & x[125]);
  assign t[223] = (x[127] & x[128]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[144] | t[33]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[25] = ~(t[145] & t[146]);
  assign t[26] = ~(t[147] & t[148]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[149] ^ t[40];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[150] ^ t[151]);
  assign t[31] = ~(t[23]);
  assign t[32] = ~(t[152] & t[41]);
  assign t[33] = ~(t[42] & t[43]);
  assign t[34] = ~(t[153]);
  assign t[35] = ~(t[140]);
  assign t[36] = t[44] & t[45];
  assign t[37] = t[46] ^ t[47];
  assign t[38] = t[48] ^ t[49];
  assign t[39] = t[50] ^ t[51];
  assign t[3] = ~(t[6]);
  assign t[40] = t[142] ^ t[154];
  assign t[41] = ~(t[155]);
  assign t[42] = ~(t[156] | t[157]);
  assign t[43] = ~(t[158] | t[159]);
  assign t[44] = t[52] ^ t[53];
  assign t[45] = t[54] ^ t[55];
  assign t[46] = t[44] & t[56];
  assign t[47] = t[57] & t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[61] ^ t[62];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[63] & t[64];
  assign t[51] = t[63] & t[65];
  assign t[52] = t[66] ^ t[67];
  assign t[53] = t[68] ^ t[69];
  assign t[54] = t[24] ? t[160] : t[70];
  assign t[55] = t[24] ? t[161] : t[71];
  assign t[56] = t[72] ^ t[73];
  assign t[57] = t[59] ^ t[52];
  assign t[58] = t[54] ^ t[74];
  assign t[59] = t[75] ^ t[76];
  assign t[5] = ~(t[9]);
  assign t[60] = t[65] ^ t[77];
  assign t[61] = t[78] & t[72];
  assign t[62] = t[79] & t[80];
  assign t[63] = t[59] ^ t[79];
  assign t[64] = t[81] ^ t[82];
  assign t[65] = t[54] ^ t[83];
  assign t[66] = t[84] & t[85];
  assign t[67] = t[84] ^ t[86];
  assign t[68] = t[87] & t[88];
  assign t[69] = t[87] ^ t[86];
  assign t[6] = ~(t[10]);
  assign t[70] = t[162] ^ t[163];
  assign t[71] = t[164] ^ t[165];
  assign t[72] = t[65] ^ t[81];
  assign t[73] = t[89] ^ t[90];
  assign t[74] = t[24] ? t[166] : t[91];
  assign t[75] = t[92] ^ t[93];
  assign t[76] = t[94] & t[84];
  assign t[77] = t[73] ^ t[95];
  assign t[78] = t[79] ^ t[53];
  assign t[79] = t[96] ^ t[97];
  assign t[7] = ~(t[11]);
  assign t[80] = t[24] ? t[167] : t[98];
  assign t[81] = t[99] ^ t[74];
  assign t[82] = t[89] ^ t[55];
  assign t[83] = t[24] ? t[168] : t[100];
  assign t[84] = t[101] ^ t[75];
  assign t[85] = t[101] & t[96];
  assign t[86] = t[102] & t[101];
  assign t[87] = t[102] ^ t[96];
  assign t[88] = t[75] & t[102];
  assign t[89] = t[24] ? t[169] : t[103];
  assign t[8] = t[12] ? t[14] : t[13];
  assign t[90] = t[24] ? t[170] : t[20];
  assign t[91] = t[171] ^ t[172];
  assign t[92] = t[104] ^ t[105];
  assign t[93] = t[106] ^ t[107];
  assign t[94] = t[96] ^ t[86];
  assign t[95] = t[83] ^ t[80];
  assign t[96] = t[108] ^ t[109];
  assign t[97] = t[110] & t[87];
  assign t[98] = t[173] ^ t[174];
  assign t[99] = t[24] ? t[175] : t[111];
  assign t[9] = t[140] & t[15];
  assign y = t[0] ? t[1] : t[138];
endmodule

module R1ind270(x, y);
 input [132:0] x;
 output y;

 wire [228:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[90] ^ t[77];
  assign t[101] = t[74] ^ t[90];
  assign t[102] = t[114] ^ t[115];
  assign t[103] = t[116] ^ t[117];
  assign t[104] = t[87] ^ t[95];
  assign t[105] = t[118] ^ t[103];
  assign t[106] = t[119] ^ t[120];
  assign t[107] = t[85] ^ t[95];
  assign t[108] = t[164] ^ t[178];
  assign t[109] = t[179] ^ t[180];
  assign t[10] = ~(t[16]);
  assign t[110] = t[181] ^ t[182];
  assign t[111] = t[121] ^ t[122];
  assign t[112] = t[123] ^ t[122];
  assign t[113] = t[183] ^ t[184];
  assign t[114] = t[124] ^ t[125];
  assign t[115] = t[81] ^ t[126];
  assign t[116] = t[81] & t[126];
  assign t[117] = t[60] & t[127];
  assign t[118] = t[128] ^ t[129];
  assign t[119] = t[60] ^ t[130];
  assign t[11] = ~(t[143]);
  assign t[120] = t[62] ^ t[59];
  assign t[121] = t[131] ^ t[132];
  assign t[122] = t[133] ^ t[117];
  assign t[123] = t[134] ^ t[135];
  assign t[124] = t[130] & t[77];
  assign t[125] = t[84] & t[66];
  assign t[126] = t[66] ^ t[78];
  assign t[127] = t[72] ^ t[136];
  assign t[128] = t[119] & t[120];
  assign t[129] = t[101] & t[59];
  assign t[12] = ~(t[17]);
  assign t[130] = t[78] ^ t[137];
  assign t[131] = t[138] ^ t[125];
  assign t[132] = t[64] & t[83];
  assign t[133] = t[46] & t[139];
  assign t[134] = t[140] ^ t[129];
  assign t[135] = t[82] & t[62];
  assign t[136] = t[97] ^ t[57];
  assign t[137] = t[56] ^ t[77];
  assign t[138] = t[66] ^ t[136];
  assign t[139] = t[60] ^ t[73];
  assign t[13] = t[18] ? t[20] : t[19];
  assign t[140] = t[101] ^ t[59];
  assign t[141] = t[185] ^ x[2];
  assign t[142] = t[186] ^ x[5];
  assign t[143] = t[187] ^ x[9];
  assign t[144] = t[188] ^ x[12];
  assign t[145] = t[189] ^ x[15];
  assign t[146] = t[190] ^ x[18];
  assign t[147] = t[191] ^ x[21];
  assign t[148] = t[192] ^ x[24];
  assign t[149] = t[193] ^ x[27];
  assign t[14] = t[18] ? t[144] : t[21];
  assign t[150] = t[194] ^ x[30];
  assign t[151] = t[195] ^ x[33];
  assign t[152] = t[196] ^ x[36];
  assign t[153] = t[197] ^ x[39];
  assign t[154] = t[198] ^ x[42];
  assign t[155] = t[199] ^ x[45];
  assign t[156] = t[200] ^ x[48];
  assign t[157] = t[201] ^ x[51];
  assign t[158] = t[202] ^ x[54];
  assign t[159] = t[203] ^ x[57];
  assign t[15] = t[18] & t[22];
  assign t[160] = t[204] ^ x[60];
  assign t[161] = t[205] ^ x[63];
  assign t[162] = t[206] ^ x[66];
  assign t[163] = t[207] ^ x[69];
  assign t[164] = t[208] ^ x[72];
  assign t[165] = t[209] ^ x[75];
  assign t[166] = t[210] ^ x[78];
  assign t[167] = t[211] ^ x[81];
  assign t[168] = t[212] ^ x[84];
  assign t[169] = t[213] ^ x[87];
  assign t[16] = ~(t[143] & t[23]);
  assign t[170] = t[214] ^ x[90];
  assign t[171] = t[215] ^ x[93];
  assign t[172] = t[216] ^ x[96];
  assign t[173] = t[217] ^ x[99];
  assign t[174] = t[218] ^ x[102];
  assign t[175] = t[219] ^ x[105];
  assign t[176] = t[220] ^ x[108];
  assign t[177] = t[221] ^ x[111];
  assign t[178] = t[222] ^ x[114];
  assign t[179] = t[223] ^ x[117];
  assign t[17] = ~(t[24]);
  assign t[180] = t[224] ^ x[120];
  assign t[181] = t[225] ^ x[123];
  assign t[182] = t[226] ^ x[126];
  assign t[183] = t[227] ^ x[129];
  assign t[184] = t[228] ^ x[132];
  assign t[185] = (x[0] & x[1]);
  assign t[186] = (x[3] & x[4]);
  assign t[187] = (x[7] & x[8]);
  assign t[188] = (x[10] & x[11]);
  assign t[189] = (x[13] & x[14]);
  assign t[18] = ~(t[25] | t[26]);
  assign t[190] = (x[16] & x[17]);
  assign t[191] = (x[19] & x[20]);
  assign t[192] = (x[22] & x[23]);
  assign t[193] = (x[25] & x[26]);
  assign t[194] = (x[28] & x[29]);
  assign t[195] = (x[31] & x[32]);
  assign t[196] = (x[34] & x[35]);
  assign t[197] = (x[37] & x[38]);
  assign t[198] = (x[40] & x[41]);
  assign t[199] = (x[43] & x[44]);
  assign t[19] = t[27] ^ t[28];
  assign t[1] = t[3] ? t[142] : t[4];
  assign t[200] = (x[46] & x[47]);
  assign t[201] = (x[49] & x[50]);
  assign t[202] = (x[52] & x[53]);
  assign t[203] = (x[55] & x[56]);
  assign t[204] = (x[58] & x[59]);
  assign t[205] = (x[61] & x[62]);
  assign t[206] = (x[64] & x[65]);
  assign t[207] = (x[67] & x[68]);
  assign t[208] = (x[70] & x[71]);
  assign t[209] = (x[73] & x[74]);
  assign t[20] = t[145] ^ t[146];
  assign t[210] = (x[76] & x[77]);
  assign t[211] = (x[79] & x[80]);
  assign t[212] = (x[82] & x[83]);
  assign t[213] = (x[85] & x[86]);
  assign t[214] = (x[88] & x[89]);
  assign t[215] = (x[91] & x[92]);
  assign t[216] = (x[94] & x[95]);
  assign t[217] = (x[97] & x[98]);
  assign t[218] = (x[100] & x[101]);
  assign t[219] = (x[103] & x[104]);
  assign t[21] = ~(t[29] ^ t[30]);
  assign t[220] = (x[106] & x[107]);
  assign t[221] = (x[109] & x[110]);
  assign t[222] = (x[112] & x[113]);
  assign t[223] = (x[115] & x[116]);
  assign t[224] = (x[118] & x[119]);
  assign t[225] = (x[121] & x[122]);
  assign t[226] = (x[124] & x[125]);
  assign t[227] = (x[127] & x[128]);
  assign t[228] = (x[130] & x[131]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[147] | t[33]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[25] = ~(t[148] & t[149]);
  assign t[26] = ~(t[150] & t[151]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[152] ^ t[153]);
  assign t[31] = ~(t[23]);
  assign t[32] = ~(t[154] & t[42]);
  assign t[33] = ~(t[43] & t[44]);
  assign t[34] = ~(t[155]);
  assign t[35] = ~(t[143]);
  assign t[36] = t[45] & t[46];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[49] ^ t[50];
  assign t[39] = t[51] ^ t[52];
  assign t[3] = ~(t[6]);
  assign t[40] = t[156] ^ t[157];
  assign t[41] = t[145] ^ t[53];
  assign t[42] = ~(t[158]);
  assign t[43] = ~(t[159] | t[160]);
  assign t[44] = ~(t[161] | t[162]);
  assign t[45] = t[54] ^ t[55];
  assign t[46] = t[56] ^ t[57];
  assign t[47] = t[58] & t[59];
  assign t[48] = t[54] & t[60];
  assign t[49] = t[61] & t[62];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[63] & t[64];
  assign t[51] = t[65] & t[66];
  assign t[52] = t[67] ^ t[68];
  assign t[53] = t[163] ^ t[164];
  assign t[54] = t[69] ^ t[70];
  assign t[55] = t[61] ^ t[63];
  assign t[56] = t[24] ? t[165] : t[20];
  assign t[57] = t[24] ? t[166] : t[71];
  assign t[58] = t[69] ^ t[61];
  assign t[59] = t[72] ^ t[73];
  assign t[5] = ~(t[9]);
  assign t[60] = t[74] ^ t[56];
  assign t[61] = t[75] ^ t[76];
  assign t[62] = t[77] ^ t[78];
  assign t[63] = t[79] ^ t[80];
  assign t[64] = t[81] ^ t[82];
  assign t[65] = t[70] ^ t[63];
  assign t[66] = t[60] ^ t[72];
  assign t[67] = t[63] & t[83];
  assign t[68] = t[65] & t[84];
  assign t[69] = t[85] ^ t[86];
  assign t[6] = ~(t[10]);
  assign t[70] = t[87] ^ t[88];
  assign t[71] = t[167] ^ t[168];
  assign t[72] = t[89] ^ t[90];
  assign t[73] = t[91] ^ t[57];
  assign t[74] = t[24] ? t[169] : t[92];
  assign t[75] = t[93] & t[94];
  assign t[76] = t[93] ^ t[95];
  assign t[77] = t[24] ? t[170] : t[96];
  assign t[78] = t[97] ^ t[91];
  assign t[79] = t[98] & t[99];
  assign t[7] = ~(t[11]);
  assign t[80] = t[98] ^ t[95];
  assign t[81] = t[74] ^ t[57];
  assign t[82] = t[78] ^ t[100];
  assign t[83] = t[77] ^ t[66];
  assign t[84] = t[101] ^ t[46];
  assign t[85] = t[102] ^ t[103];
  assign t[86] = t[104] & t[93];
  assign t[87] = t[105] ^ t[106];
  assign t[88] = t[107] & t[98];
  assign t[89] = t[24] ? t[171] : t[108];
  assign t[8] = t[12] ? t[14] : t[13];
  assign t[90] = t[24] ? t[172] : t[109];
  assign t[91] = t[24] ? t[173] : t[110];
  assign t[92] = t[163] ^ t[174];
  assign t[93] = t[111] ^ t[85];
  assign t[94] = t[111] & t[87];
  assign t[95] = t[112] & t[111];
  assign t[96] = t[175] ^ t[176];
  assign t[97] = t[24] ? t[177] : t[113];
  assign t[98] = t[112] ^ t[87];
  assign t[99] = t[85] & t[112];
  assign t[9] = t[143] & t[15];
  assign y = t[0] ? t[1] : t[141];
endmodule

module R1ind271(x, y);
 input [132:0] x;
 output y;

 wire [227:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[24] ? t[176] : t[113];
  assign t[101] = t[114] ^ t[105];
  assign t[102] = t[115] ^ t[68];
  assign t[103] = t[85] ^ t[93];
  assign t[104] = t[116] ^ t[117];
  assign t[105] = t[118] ^ t[119];
  assign t[106] = t[82] ^ t[93];
  assign t[107] = t[95] ^ t[72];
  assign t[108] = t[120] ^ t[121];
  assign t[109] = t[122] ^ t[121];
  assign t[10] = ~(t[16]);
  assign t[110] = t[177] ^ t[178];
  assign t[111] = t[179] ^ t[180];
  assign t[112] = t[24] ? t[181] : t[20];
  assign t[113] = t[182] ^ t[183];
  assign t[114] = t[123] ^ t[124];
  assign t[115] = t[55] ^ t[125];
  assign t[116] = t[126] ^ t[127];
  assign t[117] = t[78] ^ t[128];
  assign t[118] = t[78] & t[128];
  assign t[119] = t[55] & t[129];
  assign t[11] = ~(t[142]);
  assign t[120] = t[130] ^ t[131];
  assign t[121] = t[132] ^ t[119];
  assign t[122] = t[133] ^ t[134];
  assign t[123] = t[115] & t[68];
  assign t[124] = t[81] & t[87];
  assign t[125] = t[75] ^ t[135];
  assign t[126] = t[125] & t[66];
  assign t[127] = t[64] & t[80];
  assign t[128] = t[80] ^ t[75];
  assign t[129] = t[99] ^ t[136];
  assign t[12] = ~(t[17]);
  assign t[130] = t[137] ^ t[127];
  assign t[131] = t[61] & t[62];
  assign t[132] = t[57] & t[138];
  assign t[133] = t[139] ^ t[124];
  assign t[134] = t[79] & t[59];
  assign t[135] = t[70] ^ t[66];
  assign t[136] = t[94] ^ t[72];
  assign t[137] = t[80] ^ t[136];
  assign t[138] = t[55] ^ t[107];
  assign t[139] = t[81] ^ t[87];
  assign t[13] = t[18] ? t[20] : t[19];
  assign t[140] = t[184] ^ x[2];
  assign t[141] = t[185] ^ x[5];
  assign t[142] = t[186] ^ x[9];
  assign t[143] = t[187] ^ x[12];
  assign t[144] = t[188] ^ x[15];
  assign t[145] = t[189] ^ x[18];
  assign t[146] = t[190] ^ x[21];
  assign t[147] = t[191] ^ x[24];
  assign t[148] = t[192] ^ x[27];
  assign t[149] = t[193] ^ x[30];
  assign t[14] = t[18] ? t[143] : t[21];
  assign t[150] = t[194] ^ x[33];
  assign t[151] = t[195] ^ x[36];
  assign t[152] = t[196] ^ x[39];
  assign t[153] = t[197] ^ x[42];
  assign t[154] = t[198] ^ x[45];
  assign t[155] = t[199] ^ x[48];
  assign t[156] = t[200] ^ x[51];
  assign t[157] = t[201] ^ x[54];
  assign t[158] = t[202] ^ x[57];
  assign t[159] = t[203] ^ x[60];
  assign t[15] = t[18] & t[22];
  assign t[160] = t[204] ^ x[63];
  assign t[161] = t[205] ^ x[66];
  assign t[162] = t[206] ^ x[69];
  assign t[163] = t[207] ^ x[72];
  assign t[164] = t[208] ^ x[75];
  assign t[165] = t[209] ^ x[78];
  assign t[166] = t[210] ^ x[81];
  assign t[167] = t[211] ^ x[84];
  assign t[168] = t[212] ^ x[87];
  assign t[169] = t[213] ^ x[90];
  assign t[16] = ~(t[142] & t[23]);
  assign t[170] = t[214] ^ x[93];
  assign t[171] = t[215] ^ x[96];
  assign t[172] = t[216] ^ x[99];
  assign t[173] = t[217] ^ x[102];
  assign t[174] = t[218] ^ x[105];
  assign t[175] = t[219] ^ x[108];
  assign t[176] = t[220] ^ x[111];
  assign t[177] = t[221] ^ x[114];
  assign t[178] = t[222] ^ x[117];
  assign t[179] = t[223] ^ x[120];
  assign t[17] = ~(t[24]);
  assign t[180] = t[224] ^ x[123];
  assign t[181] = t[225] ^ x[126];
  assign t[182] = t[226] ^ x[129];
  assign t[183] = t[227] ^ x[132];
  assign t[184] = (x[0] & x[1]);
  assign t[185] = (x[3] & x[4]);
  assign t[186] = (x[7] & x[8]);
  assign t[187] = (x[10] & x[11]);
  assign t[188] = (x[13] & x[14]);
  assign t[189] = (x[16] & x[17]);
  assign t[18] = ~(t[25] | t[26]);
  assign t[190] = (x[19] & x[20]);
  assign t[191] = (x[22] & x[23]);
  assign t[192] = (x[25] & x[26]);
  assign t[193] = (x[28] & x[29]);
  assign t[194] = (x[31] & x[32]);
  assign t[195] = (x[34] & x[35]);
  assign t[196] = (x[37] & x[38]);
  assign t[197] = (x[40] & x[41]);
  assign t[198] = (x[43] & x[44]);
  assign t[199] = (x[46] & x[47]);
  assign t[19] = t[27] ^ t[28];
  assign t[1] = t[3] ? t[141] : t[4];
  assign t[200] = (x[49] & x[50]);
  assign t[201] = (x[52] & x[53]);
  assign t[202] = (x[55] & x[56]);
  assign t[203] = (x[58] & x[59]);
  assign t[204] = (x[61] & x[62]);
  assign t[205] = (x[64] & x[65]);
  assign t[206] = (x[67] & x[68]);
  assign t[207] = (x[70] & x[71]);
  assign t[208] = (x[73] & x[74]);
  assign t[209] = (x[76] & x[77]);
  assign t[20] = t[144] ^ t[145];
  assign t[210] = (x[79] & x[80]);
  assign t[211] = (x[82] & x[83]);
  assign t[212] = (x[85] & x[86]);
  assign t[213] = (x[88] & x[89]);
  assign t[214] = (x[91] & x[92]);
  assign t[215] = (x[94] & x[95]);
  assign t[216] = (x[97] & x[98]);
  assign t[217] = (x[100] & x[101]);
  assign t[218] = (x[103] & x[104]);
  assign t[219] = (x[106] & x[107]);
  assign t[21] = ~(t[29] ^ t[30]);
  assign t[220] = (x[109] & x[110]);
  assign t[221] = (x[112] & x[113]);
  assign t[222] = (x[115] & x[116]);
  assign t[223] = (x[118] & x[119]);
  assign t[224] = (x[121] & x[122]);
  assign t[225] = (x[124] & x[125]);
  assign t[226] = (x[127] & x[128]);
  assign t[227] = (x[130] & x[131]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[146] | t[33]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[25] = ~(t[147] & t[148]);
  assign t[26] = ~(t[149] & t[150]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[151] ^ t[152]);
  assign t[31] = ~(t[23]);
  assign t[32] = ~(t[153] & t[42]);
  assign t[33] = ~(t[43] & t[44]);
  assign t[34] = ~(t[154]);
  assign t[35] = ~(t[142]);
  assign t[36] = t[45] ^ t[46];
  assign t[37] = t[47] ^ t[48];
  assign t[38] = t[49] ^ t[50];
  assign t[39] = t[51] ^ t[52];
  assign t[3] = ~(t[6]);
  assign t[40] = t[155] ^ t[156];
  assign t[41] = t[144] ^ t[53];
  assign t[42] = ~(t[157]);
  assign t[43] = ~(t[158] | t[159]);
  assign t[44] = ~(t[160] | t[161]);
  assign t[45] = t[54] & t[55];
  assign t[46] = t[56] & t[57];
  assign t[47] = t[58] & t[59];
  assign t[48] = t[60] & t[61];
  assign t[49] = t[60] & t[62];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[63] & t[64];
  assign t[51] = t[65] & t[66];
  assign t[52] = t[67] & t[68];
  assign t[53] = t[162] ^ t[163];
  assign t[54] = t[67] ^ t[65];
  assign t[55] = t[69] ^ t[70];
  assign t[56] = t[54] ^ t[71];
  assign t[57] = t[70] ^ t[72];
  assign t[58] = t[73] ^ t[74];
  assign t[59] = t[66] ^ t[75];
  assign t[5] = ~(t[9]);
  assign t[60] = t[76] ^ t[77];
  assign t[61] = t[78] ^ t[79];
  assign t[62] = t[66] ^ t[80];
  assign t[63] = t[65] ^ t[60];
  assign t[64] = t[81] ^ t[57];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[24] ? t[164] : t[84];
  assign t[67] = t[85] ^ t[86];
  assign t[68] = t[59] ^ t[87];
  assign t[69] = t[24] ? t[165] : t[88];
  assign t[6] = ~(t[10]);
  assign t[70] = t[24] ? t[166] : t[89];
  assign t[71] = t[58] ^ t[60];
  assign t[72] = t[24] ? t[167] : t[90];
  assign t[73] = t[91] & t[92];
  assign t[74] = t[91] ^ t[93];
  assign t[75] = t[94] ^ t[95];
  assign t[76] = t[96] & t[97];
  assign t[77] = t[96] ^ t[93];
  assign t[78] = t[69] ^ t[72];
  assign t[79] = t[75] ^ t[98];
  assign t[7] = ~(t[11]);
  assign t[80] = t[55] ^ t[99];
  assign t[81] = t[69] ^ t[100];
  assign t[82] = t[101] ^ t[102];
  assign t[83] = t[103] & t[96];
  assign t[84] = t[168] ^ t[169];
  assign t[85] = t[104] ^ t[105];
  assign t[86] = t[106] & t[91];
  assign t[87] = t[99] ^ t[107];
  assign t[88] = t[162] ^ t[170];
  assign t[89] = t[171] ^ t[172];
  assign t[8] = t[12] ? t[14] : t[13];
  assign t[90] = t[163] ^ t[173];
  assign t[91] = t[108] ^ t[85];
  assign t[92] = t[108] & t[82];
  assign t[93] = t[109] & t[108];
  assign t[94] = t[24] ? t[174] : t[110];
  assign t[95] = t[24] ? t[175] : t[111];
  assign t[96] = t[109] ^ t[82];
  assign t[97] = t[85] & t[109];
  assign t[98] = t[100] ^ t[66];
  assign t[99] = t[112] ^ t[100];
  assign t[9] = t[142] & t[15];
  assign y = t[0] ? t[1] : t[140];
endmodule

module R1ind272(x, y);
 input [129:0] x;
 output y;

 wire [232:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[121] ^ t[96];
  assign t[101] = t[60] ^ t[122];
  assign t[102] = t[77] ^ t[119];
  assign t[103] = t[123] ^ t[82];
  assign t[104] = t[24] ? t[179] : t[124];
  assign t[105] = t[98] & t[125];
  assign t[106] = t[98] ^ t[119];
  assign t[107] = t[103] & t[126];
  assign t[108] = t[103] ^ t[119];
  assign t[109] = t[92] ^ t[70];
  assign t[10] = ~(t[16]);
  assign t[110] = t[84] ^ t[127];
  assign t[111] = t[24] ? t[180] : t[128];
  assign t[112] = t[181] ^ t[182];
  assign t[113] = t[183] ^ t[184];
  assign t[114] = t[163] ^ t[185];
  assign t[115] = t[129] ^ t[130];
  assign t[116] = t[109] ^ t[75];
  assign t[117] = t[109] & t[75];
  assign t[118] = t[73] & t[131];
  assign t[119] = t[123] & t[120];
  assign t[11] = ~(t[149]);
  assign t[120] = t[132] ^ t[133];
  assign t[121] = t[134] ^ t[135];
  assign t[122] = t[87] ^ t[72];
  assign t[123] = t[136] ^ t[133];
  assign t[124] = t[186] ^ t[187];
  assign t[125] = t[120] & t[82];
  assign t[126] = t[77] & t[123];
  assign t[127] = t[94] ^ t[81];
  assign t[128] = t[188] ^ t[189];
  assign t[129] = t[64] & t[81];
  assign t[12] = ~(t[17]);
  assign t[130] = t[137] & t[80];
  assign t[131] = t[91] ^ t[138];
  assign t[132] = t[139] ^ t[140];
  assign t[133] = t[141] ^ t[118];
  assign t[134] = t[60] & t[122];
  assign t[135] = t[76] & t[72];
  assign t[136] = t[142] ^ t[143];
  assign t[137] = t[76] ^ t[53];
  assign t[138] = t[104] ^ t[70];
  assign t[139] = t[144] ^ t[130];
  assign t[13] = t[18] ? t[20] : t[19];
  assign t[140] = t[89] & t[145];
  assign t[141] = t[53] & t[56];
  assign t[142] = t[146] ^ t[135];
  assign t[143] = t[110] & t[87];
  assign t[144] = t[80] ^ t[138];
  assign t[145] = t[81] ^ t[80];
  assign t[146] = t[76] ^ t[72];
  assign t[147] = t[190] ^ x[2];
  assign t[148] = t[191] ^ x[5];
  assign t[149] = t[192] ^ x[9];
  assign t[14] = t[18] ? t[150] : t[21];
  assign t[150] = t[193] ^ x[12];
  assign t[151] = t[194] ^ x[15];
  assign t[152] = t[195] ^ x[18];
  assign t[153] = t[196] ^ x[21];
  assign t[154] = t[197] ^ x[24];
  assign t[155] = t[198] ^ x[27];
  assign t[156] = t[199] ^ x[30];
  assign t[157] = t[200] ^ x[33];
  assign t[158] = t[201] ^ x[36];
  assign t[159] = t[202] ^ x[39];
  assign t[15] = t[18] & t[22];
  assign t[160] = t[203] ^ x[42];
  assign t[161] = t[204] ^ x[45];
  assign t[162] = t[205] ^ x[48];
  assign t[163] = t[206] ^ x[51];
  assign t[164] = t[207] ^ x[54];
  assign t[165] = t[208] ^ x[57];
  assign t[166] = t[209] ^ x[60];
  assign t[167] = t[210] ^ x[63];
  assign t[168] = t[211] ^ x[66];
  assign t[169] = t[212] ^ x[69];
  assign t[16] = ~(t[149] & t[23]);
  assign t[170] = t[213] ^ x[72];
  assign t[171] = t[214] ^ x[75];
  assign t[172] = t[215] ^ x[78];
  assign t[173] = t[216] ^ x[81];
  assign t[174] = t[217] ^ x[84];
  assign t[175] = t[218] ^ x[87];
  assign t[176] = t[219] ^ x[90];
  assign t[177] = t[220] ^ x[93];
  assign t[178] = t[221] ^ x[96];
  assign t[179] = t[222] ^ x[99];
  assign t[17] = ~(t[24]);
  assign t[180] = t[223] ^ x[102];
  assign t[181] = t[224] ^ x[105];
  assign t[182] = t[225] ^ x[108];
  assign t[183] = t[226] ^ x[111];
  assign t[184] = t[227] ^ x[114];
  assign t[185] = t[228] ^ x[117];
  assign t[186] = t[229] ^ x[120];
  assign t[187] = t[230] ^ x[123];
  assign t[188] = t[231] ^ x[126];
  assign t[189] = t[232] ^ x[129];
  assign t[18] = ~(t[25] | t[26]);
  assign t[190] = (x[0] & x[1]);
  assign t[191] = (x[3] & x[4]);
  assign t[192] = (x[7] & x[8]);
  assign t[193] = (x[10] & x[11]);
  assign t[194] = (x[13] & x[14]);
  assign t[195] = (x[16] & x[17]);
  assign t[196] = (x[19] & x[20]);
  assign t[197] = (x[22] & x[23]);
  assign t[198] = (x[25] & x[26]);
  assign t[199] = (x[28] & x[29]);
  assign t[19] = t[27] ^ t[28];
  assign t[1] = t[3] ? t[148] : t[4];
  assign t[200] = (x[31] & x[32]);
  assign t[201] = (x[34] & x[35]);
  assign t[202] = (x[37] & x[38]);
  assign t[203] = (x[40] & x[41]);
  assign t[204] = (x[43] & x[44]);
  assign t[205] = (x[46] & x[47]);
  assign t[206] = (x[49] & x[50]);
  assign t[207] = (x[52] & x[53]);
  assign t[208] = (x[55] & x[56]);
  assign t[209] = (x[58] & x[59]);
  assign t[20] = t[151] ^ t[152];
  assign t[210] = (x[61] & x[62]);
  assign t[211] = (x[64] & x[65]);
  assign t[212] = (x[67] & x[68]);
  assign t[213] = (x[70] & x[71]);
  assign t[214] = (x[73] & x[74]);
  assign t[215] = (x[76] & x[77]);
  assign t[216] = (x[79] & x[80]);
  assign t[217] = (x[82] & x[83]);
  assign t[218] = (x[85] & x[86]);
  assign t[219] = (x[88] & x[89]);
  assign t[21] = ~(t[29] ^ t[30]);
  assign t[220] = (x[91] & x[92]);
  assign t[221] = (x[94] & x[95]);
  assign t[222] = (x[97] & x[98]);
  assign t[223] = (x[100] & x[101]);
  assign t[224] = (x[103] & x[104]);
  assign t[225] = (x[106] & x[107]);
  assign t[226] = (x[109] & x[110]);
  assign t[227] = (x[112] & x[113]);
  assign t[228] = (x[115] & x[116]);
  assign t[229] = (x[118] & x[119]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[230] = (x[121] & x[122]);
  assign t[231] = (x[124] & x[125]);
  assign t[232] = (x[127] & x[128]);
  assign t[23] = ~(t[153] | t[33]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[25] = ~(t[154] & t[155]);
  assign t[26] = ~(t[156] & t[157]);
  assign t[27] = t[36] ^ t[37];
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[158] ^ t[40];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[159] ^ t[160]);
  assign t[31] = ~(t[23]);
  assign t[32] = ~(t[161] & t[41]);
  assign t[33] = ~(t[42] & t[43]);
  assign t[34] = ~(t[162]);
  assign t[35] = ~(t[149]);
  assign t[36] = t[44] ^ t[45];
  assign t[37] = t[46] ^ t[47];
  assign t[38] = t[48] ^ t[49];
  assign t[39] = t[50] ^ t[51];
  assign t[3] = ~(t[6]);
  assign t[40] = t[151] ^ t[163];
  assign t[41] = ~(t[164]);
  assign t[42] = ~(t[165] | t[166]);
  assign t[43] = ~(t[167] | t[168]);
  assign t[44] = t[52] & t[53];
  assign t[45] = t[54] ^ t[55];
  assign t[46] = t[52] & t[56];
  assign t[47] = t[57] ^ t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[61] ^ t[62];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[63] & t[64];
  assign t[51] = t[65] ^ t[66];
  assign t[52] = t[67] ^ t[68];
  assign t[53] = t[69] ^ t[70];
  assign t[54] = t[71] & t[72];
  assign t[55] = t[67] & t[73];
  assign t[56] = t[73] ^ t[74];
  assign t[57] = t[68] & t[75];
  assign t[58] = t[71] & t[76];
  assign t[59] = t[77] ^ t[78];
  assign t[5] = ~(t[9]);
  assign t[60] = t[73] ^ t[64];
  assign t[61] = t[79] & t[80];
  assign t[62] = t[63] & t[81];
  assign t[63] = t[82] ^ t[83];
  assign t[64] = t[84] ^ t[85];
  assign t[65] = t[86] & t[87];
  assign t[66] = t[88] & t[89];
  assign t[67] = t[59] ^ t[63];
  assign t[68] = t[86] ^ t[88];
  assign t[69] = t[24] ? t[169] : t[90];
  assign t[6] = ~(t[10]);
  assign t[70] = t[24] ? t[170] : t[20];
  assign t[71] = t[59] ^ t[86];
  assign t[72] = t[91] ^ t[74];
  assign t[73] = t[92] ^ t[69];
  assign t[74] = t[93] ^ t[70];
  assign t[75] = t[80] ^ t[84];
  assign t[76] = t[92] ^ t[94];
  assign t[77] = t[95] ^ t[96];
  assign t[78] = t[97] & t[98];
  assign t[79] = t[63] ^ t[88];
  assign t[7] = ~(t[11]);
  assign t[80] = t[73] ^ t[91];
  assign t[81] = t[24] ? t[171] : t[99];
  assign t[82] = t[100] ^ t[101];
  assign t[83] = t[102] & t[103];
  assign t[84] = t[104] ^ t[93];
  assign t[85] = t[69] ^ t[81];
  assign t[86] = t[105] ^ t[106];
  assign t[87] = t[81] ^ t[84];
  assign t[88] = t[107] ^ t[108];
  assign t[89] = t[109] ^ t[110];
  assign t[8] = t[12] ? t[14] : t[13];
  assign t[90] = t[172] ^ t[173];
  assign t[91] = t[111] ^ t[94];
  assign t[92] = t[24] ? t[174] : t[112];
  assign t[93] = t[24] ? t[175] : t[113];
  assign t[94] = t[24] ? t[176] : t[114];
  assign t[95] = t[115] ^ t[116];
  assign t[96] = t[117] ^ t[118];
  assign t[97] = t[82] ^ t[119];
  assign t[98] = t[120] ^ t[77];
  assign t[99] = t[177] ^ t[178];
  assign t[9] = t[149] & t[15];
  assign y = t[0] ? t[1] : t[147];
endmodule

module R1ind273(x, y);
 input [132:0] x;
 output y;

 wire [229:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[116] ^ t[117];
  assign t[101] = t[90] ^ t[72];
  assign t[102] = t[118] ^ t[103];
  assign t[103] = t[25] ? t[182] : t[20];
  assign t[104] = t[61] ^ t[102];
  assign t[105] = t[119] ^ t[120];
  assign t[106] = t[121] ^ t[117];
  assign t[107] = t[122] ^ t[100];
  assign t[108] = t[123] ^ t[65];
  assign t[109] = t[124] ^ t[125];
  assign t[10] = ~(t[16]);
  assign t[110] = t[81] ^ t[72];
  assign t[111] = t[91] ^ t[90];
  assign t[112] = t[111] & t[126];
  assign t[113] = t[111] ^ t[72];
  assign t[114] = t[127] ^ t[128];
  assign t[115] = t[129] ^ t[86];
  assign t[116] = t[129] & t[86];
  assign t[117] = t[61] & t[130];
  assign t[118] = t[25] ? t[183] : t[131];
  assign t[119] = t[132] ^ t[128];
  assign t[11] = ~(t[144]);
  assign t[120] = t[133] & t[134];
  assign t[121] = t[63] & t[67];
  assign t[122] = t[135] ^ t[136];
  assign t[123] = t[61] ^ t[137];
  assign t[124] = t[138] ^ t[136];
  assign t[125] = t[66] & t[48];
  assign t[126] = t[81] & t[91];
  assign t[127] = t[137] & t[58];
  assign t[128] = t[139] & t[104];
  assign t[129] = t[77] ^ t[80];
  assign t[12] = ~(t[17]);
  assign t[130] = t[102] ^ t[140];
  assign t[131] = t[184] ^ t[185];
  assign t[132] = t[104] ^ t[140];
  assign t[133] = t[129] ^ t[66];
  assign t[134] = t[58] ^ t[104];
  assign t[135] = t[123] & t[65];
  assign t[136] = t[88] & t[83];
  assign t[137] = t[59] ^ t[141];
  assign t[138] = t[88] ^ t[83];
  assign t[139] = t[88] ^ t[63];
  assign t[13] = t[18] ? t[20] : t[19];
  assign t[140] = t[74] ^ t[80];
  assign t[141] = t[78] ^ t[58];
  assign t[142] = t[186] ^ x[2];
  assign t[143] = t[187] ^ x[5];
  assign t[144] = t[188] ^ x[9];
  assign t[145] = t[189] ^ x[12];
  assign t[146] = t[190] ^ x[15];
  assign t[147] = t[191] ^ x[18];
  assign t[148] = t[192] ^ x[21];
  assign t[149] = t[193] ^ x[24];
  assign t[14] = t[21] ? t[145] : t[22];
  assign t[150] = t[194] ^ x[27];
  assign t[151] = t[195] ^ x[30];
  assign t[152] = t[196] ^ x[33];
  assign t[153] = t[197] ^ x[36];
  assign t[154] = t[198] ^ x[39];
  assign t[155] = t[199] ^ x[42];
  assign t[156] = t[200] ^ x[45];
  assign t[157] = t[201] ^ x[48];
  assign t[158] = t[202] ^ x[51];
  assign t[159] = t[203] ^ x[54];
  assign t[15] = t[18] & t[23];
  assign t[160] = t[204] ^ x[57];
  assign t[161] = t[205] ^ x[60];
  assign t[162] = t[206] ^ x[63];
  assign t[163] = t[207] ^ x[66];
  assign t[164] = t[208] ^ x[69];
  assign t[165] = t[209] ^ x[72];
  assign t[166] = t[210] ^ x[75];
  assign t[167] = t[211] ^ x[78];
  assign t[168] = t[212] ^ x[81];
  assign t[169] = t[213] ^ x[84];
  assign t[16] = ~(t[144] & t[24]);
  assign t[170] = t[214] ^ x[87];
  assign t[171] = t[215] ^ x[90];
  assign t[172] = t[216] ^ x[93];
  assign t[173] = t[217] ^ x[96];
  assign t[174] = t[218] ^ x[99];
  assign t[175] = t[219] ^ x[102];
  assign t[176] = t[220] ^ x[105];
  assign t[177] = t[221] ^ x[108];
  assign t[178] = t[222] ^ x[111];
  assign t[179] = t[223] ^ x[114];
  assign t[17] = ~(t[25]);
  assign t[180] = t[224] ^ x[117];
  assign t[181] = t[225] ^ x[120];
  assign t[182] = t[226] ^ x[123];
  assign t[183] = t[227] ^ x[126];
  assign t[184] = t[228] ^ x[129];
  assign t[185] = t[229] ^ x[132];
  assign t[186] = (x[0] & x[1]);
  assign t[187] = (x[3] & x[4]);
  assign t[188] = (x[7] & x[8]);
  assign t[189] = (x[10] & x[11]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[190] = (x[13] & x[14]);
  assign t[191] = (x[16] & x[17]);
  assign t[192] = (x[19] & x[20]);
  assign t[193] = (x[22] & x[23]);
  assign t[194] = (x[25] & x[26]);
  assign t[195] = (x[28] & x[29]);
  assign t[196] = (x[31] & x[32]);
  assign t[197] = (x[34] & x[35]);
  assign t[198] = (x[37] & x[38]);
  assign t[199] = (x[40] & x[41]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = t[3] ? t[143] : t[4];
  assign t[200] = (x[43] & x[44]);
  assign t[201] = (x[46] & x[47]);
  assign t[202] = (x[49] & x[50]);
  assign t[203] = (x[52] & x[53]);
  assign t[204] = (x[55] & x[56]);
  assign t[205] = (x[58] & x[59]);
  assign t[206] = (x[61] & x[62]);
  assign t[207] = (x[64] & x[65]);
  assign t[208] = (x[67] & x[68]);
  assign t[209] = (x[70] & x[71]);
  assign t[20] = t[146] ^ t[147];
  assign t[210] = (x[73] & x[74]);
  assign t[211] = (x[76] & x[77]);
  assign t[212] = (x[79] & x[80]);
  assign t[213] = (x[82] & x[83]);
  assign t[214] = (x[85] & x[86]);
  assign t[215] = (x[88] & x[89]);
  assign t[216] = (x[91] & x[92]);
  assign t[217] = (x[94] & x[95]);
  assign t[218] = (x[97] & x[98]);
  assign t[219] = (x[100] & x[101]);
  assign t[21] = ~(t[30]);
  assign t[220] = (x[103] & x[104]);
  assign t[221] = (x[106] & x[107]);
  assign t[222] = (x[109] & x[110]);
  assign t[223] = (x[112] & x[113]);
  assign t[224] = (x[115] & x[116]);
  assign t[225] = (x[118] & x[119]);
  assign t[226] = (x[121] & x[122]);
  assign t[227] = (x[124] & x[125]);
  assign t[228] = (x[127] & x[128]);
  assign t[229] = (x[130] & x[131]);
  assign t[22] = ~(t[31] ^ t[32]);
  assign t[23] = ~(t[33] | t[34]);
  assign t[24] = ~(t[148] | t[35]);
  assign t[25] = ~(t[36] | t[37]);
  assign t[26] = ~(t[149] & t[150]);
  assign t[27] = ~(t[151] & t[152]);
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[18]);
  assign t[31] = t[42] ^ t[43];
  assign t[32] = ~(t[153] ^ t[154]);
  assign t[33] = ~(t[24]);
  assign t[34] = ~(t[155] & t[44]);
  assign t[35] = ~(t[45] & t[46]);
  assign t[36] = ~(t[156]);
  assign t[37] = ~(t[144]);
  assign t[38] = t[47] & t[48];
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ t[52];
  assign t[41] = t[53] ^ t[54];
  assign t[42] = t[157] ^ t[158];
  assign t[43] = t[146] ^ t[55];
  assign t[44] = ~(t[159]);
  assign t[45] = ~(t[160] | t[161]);
  assign t[46] = ~(t[162] | t[163]);
  assign t[47] = t[56] ^ t[57];
  assign t[48] = t[58] ^ t[59];
  assign t[49] = t[60] & t[61];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[62] & t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[47] & t[66];
  assign t[53] = t[62] & t[67];
  assign t[54] = t[68] ^ t[69];
  assign t[55] = t[164] ^ t[165];
  assign t[56] = t[70] & t[71];
  assign t[57] = t[70] ^ t[72];
  assign t[58] = t[25] ? t[166] : t[73];
  assign t[59] = t[74] ^ t[75];
  assign t[5] = ~(t[9]);
  assign t[60] = t[64] ^ t[76];
  assign t[61] = t[77] ^ t[78];
  assign t[62] = t[60] ^ t[79];
  assign t[63] = t[78] ^ t[80];
  assign t[64] = t[81] ^ t[82];
  assign t[65] = t[48] ^ t[83];
  assign t[66] = t[59] ^ t[84];
  assign t[67] = t[61] ^ t[85];
  assign t[68] = t[79] & t[86];
  assign t[69] = t[87] & t[88];
  assign t[6] = ~(t[10]);
  assign t[70] = t[89] ^ t[81];
  assign t[71] = t[89] & t[90];
  assign t[72] = t[91] & t[89];
  assign t[73] = t[165] ^ t[167];
  assign t[74] = t[25] ? t[168] : t[92];
  assign t[75] = t[25] ? t[169] : t[93];
  assign t[76] = t[90] ^ t[94];
  assign t[77] = t[25] ? t[170] : t[95];
  assign t[78] = t[25] ? t[171] : t[96];
  assign t[79] = t[47] ^ t[97];
  assign t[7] = ~(t[11]);
  assign t[80] = t[25] ? t[172] : t[98];
  assign t[81] = t[99] ^ t[100];
  assign t[82] = t[101] & t[70];
  assign t[83] = t[102] ^ t[85];
  assign t[84] = t[103] ^ t[58];
  assign t[85] = t[75] ^ t[80];
  assign t[86] = t[104] ^ t[59];
  assign t[87] = t[64] ^ t[47];
  assign t[88] = t[77] ^ t[103];
  assign t[89] = t[105] ^ t[106];
  assign t[8] = t[12] ? t[14] : t[13];
  assign t[90] = t[107] ^ t[108];
  assign t[91] = t[109] ^ t[106];
  assign t[92] = t[173] ^ t[174];
  assign t[93] = t[175] ^ t[176];
  assign t[94] = t[110] & t[111];
  assign t[95] = t[164] ^ t[177];
  assign t[96] = t[178] ^ t[179];
  assign t[97] = t[112] ^ t[113];
  assign t[98] = t[180] ^ t[181];
  assign t[99] = t[114] ^ t[115];
  assign t[9] = t[144] & t[15];
  assign y = t[0] ? t[1] : t[142];
endmodule

module R1ind274(x, y);
 input [129:0] x;
 output y;

 wire [226:0] t;
  assign t[0] = ~(t[2]);
  assign t[100] = t[79] ^ t[103];
  assign t[101] = t[115] ^ t[81];
  assign t[102] = t[115] & t[79];
  assign t[103] = t[110] & t[115];
  assign t[104] = t[81] & t[110];
  assign t[105] = t[177] ^ t[178];
  assign t[106] = t[179] ^ t[180];
  assign t[107] = t[25] ? t[181] : t[116];
  assign t[108] = t[117] ^ t[118];
  assign t[109] = t[60] ^ t[119];
  assign t[10] = ~(t[16]);
  assign t[110] = t[120] ^ t[121];
  assign t[111] = t[122] ^ t[123];
  assign t[112] = t[124] ^ t[125];
  assign t[113] = t[124] & t[125];
  assign t[114] = t[60] & t[126];
  assign t[115] = t[127] ^ t[121];
  assign t[116] = t[182] ^ t[183];
  assign t[117] = t[109] & t[77];
  assign t[118] = t[61] & t[59];
  assign t[119] = t[92] ^ t[128];
  assign t[11] = ~(t[143]);
  assign t[120] = t[129] ^ t[130];
  assign t[121] = t[131] ^ t[114];
  assign t[122] = t[119] & t[67];
  assign t[123] = t[132] & t[65];
  assign t[124] = t[75] ^ t[57];
  assign t[125] = t[65] ^ t[92];
  assign t[126] = t[73] ^ t[133];
  assign t[127] = t[134] ^ t[135];
  assign t[128] = t[56] ^ t[67];
  assign t[129] = t[136] ^ t[118];
  assign t[12] = ~(t[17]);
  assign t[130] = t[78] & t[91];
  assign t[131] = t[47] & t[137];
  assign t[132] = t[61] ^ t[47];
  assign t[133] = t[107] ^ t[57];
  assign t[134] = t[138] ^ t[123];
  assign t[135] = t[139] & t[140];
  assign t[136] = t[61] ^ t[59];
  assign t[137] = t[60] ^ t[74];
  assign t[138] = t[65] ^ t[133];
  assign t[139] = t[124] ^ t[78];
  assign t[13] = t[18] ? t[20] : t[19];
  assign t[140] = t[67] ^ t[65];
  assign t[141] = t[184] ^ x[2];
  assign t[142] = t[185] ^ x[5];
  assign t[143] = t[186] ^ x[9];
  assign t[144] = t[187] ^ x[12];
  assign t[145] = t[188] ^ x[15];
  assign t[146] = t[189] ^ x[18];
  assign t[147] = t[190] ^ x[21];
  assign t[148] = t[191] ^ x[24];
  assign t[149] = t[192] ^ x[27];
  assign t[14] = t[21] ? t[144] : t[22];
  assign t[150] = t[193] ^ x[30];
  assign t[151] = t[194] ^ x[33];
  assign t[152] = t[195] ^ x[36];
  assign t[153] = t[196] ^ x[39];
  assign t[154] = t[197] ^ x[42];
  assign t[155] = t[198] ^ x[45];
  assign t[156] = t[199] ^ x[48];
  assign t[157] = t[200] ^ x[51];
  assign t[158] = t[201] ^ x[54];
  assign t[159] = t[202] ^ x[57];
  assign t[15] = t[18] & t[23];
  assign t[160] = t[203] ^ x[60];
  assign t[161] = t[204] ^ x[63];
  assign t[162] = t[205] ^ x[66];
  assign t[163] = t[206] ^ x[69];
  assign t[164] = t[207] ^ x[72];
  assign t[165] = t[208] ^ x[75];
  assign t[166] = t[209] ^ x[78];
  assign t[167] = t[210] ^ x[81];
  assign t[168] = t[211] ^ x[84];
  assign t[169] = t[212] ^ x[87];
  assign t[16] = ~(t[143] & t[24]);
  assign t[170] = t[213] ^ x[90];
  assign t[171] = t[214] ^ x[93];
  assign t[172] = t[215] ^ x[96];
  assign t[173] = t[216] ^ x[99];
  assign t[174] = t[217] ^ x[102];
  assign t[175] = t[218] ^ x[105];
  assign t[176] = t[219] ^ x[108];
  assign t[177] = t[220] ^ x[111];
  assign t[178] = t[221] ^ x[114];
  assign t[179] = t[222] ^ x[117];
  assign t[17] = ~(t[25]);
  assign t[180] = t[223] ^ x[120];
  assign t[181] = t[224] ^ x[123];
  assign t[182] = t[225] ^ x[126];
  assign t[183] = t[226] ^ x[129];
  assign t[184] = (x[0] & x[1]);
  assign t[185] = (x[3] & x[4]);
  assign t[186] = (x[7] & x[8]);
  assign t[187] = (x[10] & x[11]);
  assign t[188] = (x[13] & x[14]);
  assign t[189] = (x[16] & x[17]);
  assign t[18] = ~(t[26] | t[27]);
  assign t[190] = (x[19] & x[20]);
  assign t[191] = (x[22] & x[23]);
  assign t[192] = (x[25] & x[26]);
  assign t[193] = (x[28] & x[29]);
  assign t[194] = (x[31] & x[32]);
  assign t[195] = (x[34] & x[35]);
  assign t[196] = (x[37] & x[38]);
  assign t[197] = (x[40] & x[41]);
  assign t[198] = (x[43] & x[44]);
  assign t[199] = (x[46] & x[47]);
  assign t[19] = ~(t[28] ^ t[29]);
  assign t[1] = t[3] ? t[142] : t[4];
  assign t[200] = (x[49] & x[50]);
  assign t[201] = (x[52] & x[53]);
  assign t[202] = (x[55] & x[56]);
  assign t[203] = (x[58] & x[59]);
  assign t[204] = (x[61] & x[62]);
  assign t[205] = (x[64] & x[65]);
  assign t[206] = (x[67] & x[68]);
  assign t[207] = (x[70] & x[71]);
  assign t[208] = (x[73] & x[74]);
  assign t[209] = (x[76] & x[77]);
  assign t[20] = t[145] ^ t[146];
  assign t[210] = (x[79] & x[80]);
  assign t[211] = (x[82] & x[83]);
  assign t[212] = (x[85] & x[86]);
  assign t[213] = (x[88] & x[89]);
  assign t[214] = (x[91] & x[92]);
  assign t[215] = (x[94] & x[95]);
  assign t[216] = (x[97] & x[98]);
  assign t[217] = (x[100] & x[101]);
  assign t[218] = (x[103] & x[104]);
  assign t[219] = (x[106] & x[107]);
  assign t[21] = ~(t[30]);
  assign t[220] = (x[109] & x[110]);
  assign t[221] = (x[112] & x[113]);
  assign t[222] = (x[115] & x[116]);
  assign t[223] = (x[118] & x[119]);
  assign t[224] = (x[121] & x[122]);
  assign t[225] = (x[124] & x[125]);
  assign t[226] = (x[127] & x[128]);
  assign t[22] = ~(t[31] ^ t[32]);
  assign t[23] = ~(t[33] | t[34]);
  assign t[24] = ~(t[147] | t[35]);
  assign t[25] = ~(t[36] | t[37]);
  assign t[26] = ~(t[148] & t[149]);
  assign t[27] = ~(t[150] & t[151]);
  assign t[28] = t[38] ^ t[39];
  assign t[29] = t[40] ^ t[41];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[18]);
  assign t[31] = t[152] ^ t[42];
  assign t[32] = ~(t[153] ^ t[154]);
  assign t[33] = ~(t[24]);
  assign t[34] = ~(t[155] & t[43]);
  assign t[35] = ~(t[44] & t[45]);
  assign t[36] = ~(t[156]);
  assign t[37] = ~(t[143]);
  assign t[38] = t[46] & t[47];
  assign t[39] = t[48] ^ t[49];
  assign t[3] = ~(t[6]);
  assign t[40] = t[50] ^ t[51];
  assign t[41] = t[52] ^ t[53];
  assign t[42] = t[145] ^ t[157];
  assign t[43] = ~(t[158]);
  assign t[44] = ~(t[159] | t[160]);
  assign t[45] = ~(t[161] | t[162]);
  assign t[46] = t[54] ^ t[55];
  assign t[47] = t[56] ^ t[57];
  assign t[48] = t[58] & t[59];
  assign t[49] = t[54] & t[60];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[58] & t[61];
  assign t[51] = t[62] ^ t[63];
  assign t[52] = t[64] & t[65];
  assign t[53] = t[66] & t[67];
  assign t[54] = t[68] ^ t[66];
  assign t[55] = t[69] ^ t[70];
  assign t[56] = t[25] ? t[163] : t[71];
  assign t[57] = t[25] ? t[164] : t[72];
  assign t[58] = t[68] ^ t[69];
  assign t[59] = t[73] ^ t[74];
  assign t[5] = ~(t[9]);
  assign t[60] = t[75] ^ t[56];
  assign t[61] = t[75] ^ t[76];
  assign t[62] = t[68] & t[77];
  assign t[63] = t[69] & t[78];
  assign t[64] = t[66] ^ t[70];
  assign t[65] = t[60] ^ t[73];
  assign t[66] = t[79] ^ t[80];
  assign t[67] = t[25] ? t[165] : t[20];
  assign t[68] = t[81] ^ t[82];
  assign t[69] = t[83] ^ t[84];
  assign t[6] = ~(t[10]);
  assign t[70] = t[85] ^ t[86];
  assign t[71] = t[166] ^ t[167];
  assign t[72] = t[168] ^ t[169];
  assign t[73] = t[87] ^ t[76];
  assign t[74] = t[88] ^ t[57];
  assign t[75] = t[25] ? t[170] : t[89];
  assign t[76] = t[25] ? t[171] : t[90];
  assign t[77] = t[91] ^ t[59];
  assign t[78] = t[92] ^ t[93];
  assign t[79] = t[94] ^ t[95];
  assign t[7] = ~(t[11]);
  assign t[80] = t[96] & t[97];
  assign t[81] = t[98] ^ t[99];
  assign t[82] = t[100] & t[101];
  assign t[83] = t[101] & t[102];
  assign t[84] = t[101] ^ t[103];
  assign t[85] = t[97] & t[104];
  assign t[86] = t[97] ^ t[103];
  assign t[87] = t[25] ? t[172] : t[105];
  assign t[88] = t[25] ? t[173] : t[106];
  assign t[89] = t[157] ^ t[174];
  assign t[8] = t[12] ? t[14] : t[13];
  assign t[90] = t[175] ^ t[176];
  assign t[91] = t[67] ^ t[92];
  assign t[92] = t[107] ^ t[88];
  assign t[93] = t[76] ^ t[67];
  assign t[94] = t[108] ^ t[99];
  assign t[95] = t[109] ^ t[77];
  assign t[96] = t[81] ^ t[103];
  assign t[97] = t[110] ^ t[79];
  assign t[98] = t[111] ^ t[112];
  assign t[99] = t[113] ^ t[114];
  assign t[9] = t[143] & t[15];
  assign y = t[0] ? t[1] : t[141];
endmodule

module R1ind275(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind276(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind277(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind278(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind279(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind280(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind281(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind282(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind283(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind284(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind285(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind286(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind287(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind288(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind289(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind290(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind291(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind292(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind293(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind294(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind295(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind296(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind297(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind298(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind299(x, y);
 input [63:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[40]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[41] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[40] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[38] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[42] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[43] ^ t[33];
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[50] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[40]);
  assign t[33] = t[39] ^ t[52];
  assign t[34] = ~(t[53]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = t[58] ^ x[2];
  assign t[38] = t[59] ^ x[5];
  assign t[39] = t[60] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[61] ^ x[12];
  assign t[41] = t[62] ^ x[15];
  assign t[42] = t[63] ^ x[18];
  assign t[43] = t[64] ^ x[21];
  assign t[44] = t[65] ^ x[24];
  assign t[45] = t[66] ^ x[27];
  assign t[46] = t[67] ^ x[30];
  assign t[47] = t[68] ^ x[33];
  assign t[48] = t[69] ^ x[36];
  assign t[49] = t[70] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[71] ^ x[42];
  assign t[51] = t[72] ^ x[45];
  assign t[52] = t[73] ^ x[48];
  assign t[53] = t[74] ^ x[51];
  assign t[54] = t[75] ^ x[54];
  assign t[55] = t[76] ^ x[57];
  assign t[56] = t[77] ^ x[60];
  assign t[57] = t[78] ^ x[63];
  assign t[58] = (x[0] & x[1]);
  assign t[59] = (x[3] & x[4]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[7] & x[8]);
  assign t[61] = (x[10] & x[11]);
  assign t[62] = (x[13] & x[14]);
  assign t[63] = (x[16] & x[17]);
  assign t[64] = (x[19] & x[20]);
  assign t[65] = (x[22] & x[23]);
  assign t[66] = (x[25] & x[26]);
  assign t[67] = (x[28] & x[29]);
  assign t[68] = (x[31] & x[32]);
  assign t[69] = (x[34] & x[35]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[37] & x[38]);
  assign t[71] = (x[40] & x[41]);
  assign t[72] = (x[43] & x[44]);
  assign t[73] = (x[46] & x[47]);
  assign t[74] = (x[49] & x[50]);
  assign t[75] = (x[52] & x[53]);
  assign t[76] = (x[55] & x[56]);
  assign t[77] = (x[58] & x[59]);
  assign t[78] = (x[61] & x[62]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[39];
  assign t[9] = t[40] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind300(x, y);
 input [63:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[40]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[41] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[40] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[38] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[42] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[43] ^ t[33];
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[50] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[40]);
  assign t[33] = t[39] ^ t[52];
  assign t[34] = ~(t[53]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = t[58] ^ x[2];
  assign t[38] = t[59] ^ x[5];
  assign t[39] = t[60] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[61] ^ x[12];
  assign t[41] = t[62] ^ x[15];
  assign t[42] = t[63] ^ x[18];
  assign t[43] = t[64] ^ x[21];
  assign t[44] = t[65] ^ x[24];
  assign t[45] = t[66] ^ x[27];
  assign t[46] = t[67] ^ x[30];
  assign t[47] = t[68] ^ x[33];
  assign t[48] = t[69] ^ x[36];
  assign t[49] = t[70] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[71] ^ x[42];
  assign t[51] = t[72] ^ x[45];
  assign t[52] = t[73] ^ x[48];
  assign t[53] = t[74] ^ x[51];
  assign t[54] = t[75] ^ x[54];
  assign t[55] = t[76] ^ x[57];
  assign t[56] = t[77] ^ x[60];
  assign t[57] = t[78] ^ x[63];
  assign t[58] = (x[0] & x[1]);
  assign t[59] = (x[3] & x[4]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[7] & x[8]);
  assign t[61] = (x[10] & x[11]);
  assign t[62] = (x[13] & x[14]);
  assign t[63] = (x[16] & x[17]);
  assign t[64] = (x[19] & x[20]);
  assign t[65] = (x[22] & x[23]);
  assign t[66] = (x[25] & x[26]);
  assign t[67] = (x[28] & x[29]);
  assign t[68] = (x[31] & x[32]);
  assign t[69] = (x[34] & x[35]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[37] & x[38]);
  assign t[71] = (x[40] & x[41]);
  assign t[72] = (x[43] & x[44]);
  assign t[73] = (x[46] & x[47]);
  assign t[74] = (x[49] & x[50]);
  assign t[75] = (x[52] & x[53]);
  assign t[76] = (x[55] & x[56]);
  assign t[77] = (x[58] & x[59]);
  assign t[78] = (x[61] & x[62]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[39];
  assign t[9] = t[40] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind301(x, y);
 input [63:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[40]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[41] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[40] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[38] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[42] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[43] ^ t[33];
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[50] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[40]);
  assign t[33] = t[39] ^ t[52];
  assign t[34] = ~(t[53]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = t[58] ^ x[2];
  assign t[38] = t[59] ^ x[5];
  assign t[39] = t[60] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[61] ^ x[12];
  assign t[41] = t[62] ^ x[15];
  assign t[42] = t[63] ^ x[18];
  assign t[43] = t[64] ^ x[21];
  assign t[44] = t[65] ^ x[24];
  assign t[45] = t[66] ^ x[27];
  assign t[46] = t[67] ^ x[30];
  assign t[47] = t[68] ^ x[33];
  assign t[48] = t[69] ^ x[36];
  assign t[49] = t[70] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[71] ^ x[42];
  assign t[51] = t[72] ^ x[45];
  assign t[52] = t[73] ^ x[48];
  assign t[53] = t[74] ^ x[51];
  assign t[54] = t[75] ^ x[54];
  assign t[55] = t[76] ^ x[57];
  assign t[56] = t[77] ^ x[60];
  assign t[57] = t[78] ^ x[63];
  assign t[58] = (x[0] & x[1]);
  assign t[59] = (x[3] & x[4]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[7] & x[8]);
  assign t[61] = (x[10] & x[11]);
  assign t[62] = (x[13] & x[14]);
  assign t[63] = (x[16] & x[17]);
  assign t[64] = (x[19] & x[20]);
  assign t[65] = (x[22] & x[23]);
  assign t[66] = (x[25] & x[26]);
  assign t[67] = (x[28] & x[29]);
  assign t[68] = (x[31] & x[32]);
  assign t[69] = (x[34] & x[35]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[37] & x[38]);
  assign t[71] = (x[40] & x[41]);
  assign t[72] = (x[43] & x[44]);
  assign t[73] = (x[46] & x[47]);
  assign t[74] = (x[49] & x[50]);
  assign t[75] = (x[52] & x[53]);
  assign t[76] = (x[55] & x[56]);
  assign t[77] = (x[58] & x[59]);
  assign t[78] = (x[61] & x[62]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[39];
  assign t[9] = t[40] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind302(x, y);
 input [69:0] x;
 output y;

 wire [84:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[42]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[43] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[42] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[40] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[44] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49] & t[50]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[51] & t[35]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[36] & t[37]);
  assign t[31] = ~(t[52]);
  assign t[32] = ~(t[42]);
  assign t[33] = t[53] ^ t[54];
  assign t[34] = t[41] ^ t[38];
  assign t[35] = ~(t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[62] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[63] ^ x[5];
  assign t[41] = t[64] ^ x[9];
  assign t[42] = t[65] ^ x[12];
  assign t[43] = t[66] ^ x[15];
  assign t[44] = t[67] ^ x[18];
  assign t[45] = t[68] ^ x[21];
  assign t[46] = t[69] ^ x[24];
  assign t[47] = t[70] ^ x[27];
  assign t[48] = t[71] ^ x[30];
  assign t[49] = t[72] ^ x[33];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[73] ^ x[36];
  assign t[51] = t[74] ^ x[39];
  assign t[52] = t[75] ^ x[42];
  assign t[53] = t[76] ^ x[45];
  assign t[54] = t[77] ^ x[48];
  assign t[55] = t[78] ^ x[51];
  assign t[56] = t[79] ^ x[54];
  assign t[57] = t[80] ^ x[57];
  assign t[58] = t[81] ^ x[60];
  assign t[59] = t[82] ^ x[63];
  assign t[5] = ~(t[9]);
  assign t[60] = t[83] ^ x[66];
  assign t[61] = t[84] ^ x[69];
  assign t[62] = (x[0] & x[1]);
  assign t[63] = (x[3] & x[4]);
  assign t[64] = (x[7] & x[8]);
  assign t[65] = (x[10] & x[11]);
  assign t[66] = (x[13] & x[14]);
  assign t[67] = (x[16] & x[17]);
  assign t[68] = (x[19] & x[20]);
  assign t[69] = (x[22] & x[23]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[25] & x[26]);
  assign t[71] = (x[28] & x[29]);
  assign t[72] = (x[31] & x[32]);
  assign t[73] = (x[34] & x[35]);
  assign t[74] = (x[37] & x[38]);
  assign t[75] = (x[40] & x[41]);
  assign t[76] = (x[43] & x[44]);
  assign t[77] = (x[46] & x[47]);
  assign t[78] = (x[49] & x[50]);
  assign t[79] = (x[52] & x[53]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[55] & x[56]);
  assign t[81] = (x[58] & x[59]);
  assign t[82] = (x[61] & x[62]);
  assign t[83] = (x[64] & x[65]);
  assign t[84] = (x[67] & x[68]);
  assign t[8] = t[12] ? t[13] : t[41];
  assign t[9] = t[42] & t[14];
  assign y = t[0] ? t[1] : t[39];
endmodule

module R1ind303(x, y);
 input [69:0] x;
 output y;

 wire [84:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[42]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[43] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[42] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[40] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[44] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49] & t[50]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[51] & t[35]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[36] & t[37]);
  assign t[31] = ~(t[52]);
  assign t[32] = ~(t[42]);
  assign t[33] = t[53] ^ t[54];
  assign t[34] = t[41] ^ t[38];
  assign t[35] = ~(t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[62] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[63] ^ x[5];
  assign t[41] = t[64] ^ x[9];
  assign t[42] = t[65] ^ x[12];
  assign t[43] = t[66] ^ x[15];
  assign t[44] = t[67] ^ x[18];
  assign t[45] = t[68] ^ x[21];
  assign t[46] = t[69] ^ x[24];
  assign t[47] = t[70] ^ x[27];
  assign t[48] = t[71] ^ x[30];
  assign t[49] = t[72] ^ x[33];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[73] ^ x[36];
  assign t[51] = t[74] ^ x[39];
  assign t[52] = t[75] ^ x[42];
  assign t[53] = t[76] ^ x[45];
  assign t[54] = t[77] ^ x[48];
  assign t[55] = t[78] ^ x[51];
  assign t[56] = t[79] ^ x[54];
  assign t[57] = t[80] ^ x[57];
  assign t[58] = t[81] ^ x[60];
  assign t[59] = t[82] ^ x[63];
  assign t[5] = ~(t[9]);
  assign t[60] = t[83] ^ x[66];
  assign t[61] = t[84] ^ x[69];
  assign t[62] = (x[0] & x[1]);
  assign t[63] = (x[3] & x[4]);
  assign t[64] = (x[7] & x[8]);
  assign t[65] = (x[10] & x[11]);
  assign t[66] = (x[13] & x[14]);
  assign t[67] = (x[16] & x[17]);
  assign t[68] = (x[19] & x[20]);
  assign t[69] = (x[22] & x[23]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[25] & x[26]);
  assign t[71] = (x[28] & x[29]);
  assign t[72] = (x[31] & x[32]);
  assign t[73] = (x[34] & x[35]);
  assign t[74] = (x[37] & x[38]);
  assign t[75] = (x[40] & x[41]);
  assign t[76] = (x[43] & x[44]);
  assign t[77] = (x[46] & x[47]);
  assign t[78] = (x[49] & x[50]);
  assign t[79] = (x[52] & x[53]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[55] & x[56]);
  assign t[81] = (x[58] & x[59]);
  assign t[82] = (x[61] & x[62]);
  assign t[83] = (x[64] & x[65]);
  assign t[84] = (x[67] & x[68]);
  assign t[8] = t[12] ? t[13] : t[41];
  assign t[9] = t[42] & t[14];
  assign y = t[0] ? t[1] : t[39];
endmodule

module R1ind304(x, y);
 input [63:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[40]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[41] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[40] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[38] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[42] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[43] ^ t[33];
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[50] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[40]);
  assign t[33] = t[39] ^ t[52];
  assign t[34] = ~(t[53]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = t[58] ^ x[2];
  assign t[38] = t[59] ^ x[5];
  assign t[39] = t[60] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[61] ^ x[12];
  assign t[41] = t[62] ^ x[15];
  assign t[42] = t[63] ^ x[18];
  assign t[43] = t[64] ^ x[21];
  assign t[44] = t[65] ^ x[24];
  assign t[45] = t[66] ^ x[27];
  assign t[46] = t[67] ^ x[30];
  assign t[47] = t[68] ^ x[33];
  assign t[48] = t[69] ^ x[36];
  assign t[49] = t[70] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[71] ^ x[42];
  assign t[51] = t[72] ^ x[45];
  assign t[52] = t[73] ^ x[48];
  assign t[53] = t[74] ^ x[51];
  assign t[54] = t[75] ^ x[54];
  assign t[55] = t[76] ^ x[57];
  assign t[56] = t[77] ^ x[60];
  assign t[57] = t[78] ^ x[63];
  assign t[58] = (x[0] & x[1]);
  assign t[59] = (x[3] & x[4]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[7] & x[8]);
  assign t[61] = (x[10] & x[11]);
  assign t[62] = (x[13] & x[14]);
  assign t[63] = (x[16] & x[17]);
  assign t[64] = (x[19] & x[20]);
  assign t[65] = (x[22] & x[23]);
  assign t[66] = (x[25] & x[26]);
  assign t[67] = (x[28] & x[29]);
  assign t[68] = (x[31] & x[32]);
  assign t[69] = (x[34] & x[35]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[37] & x[38]);
  assign t[71] = (x[40] & x[41]);
  assign t[72] = (x[43] & x[44]);
  assign t[73] = (x[46] & x[47]);
  assign t[74] = (x[49] & x[50]);
  assign t[75] = (x[52] & x[53]);
  assign t[76] = (x[55] & x[56]);
  assign t[77] = (x[58] & x[59]);
  assign t[78] = (x[61] & x[62]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[39];
  assign t[9] = t[40] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind305(x, y);
 input [69:0] x;
 output y;

 wire [84:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[42]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[43] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[42] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[40] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[44] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[45] ^ t[46]);
  assign t[26] = ~(t[47] & t[48]);
  assign t[27] = ~(t[49] & t[50]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[51] & t[35]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[36] & t[37]);
  assign t[31] = ~(t[52]);
  assign t[32] = ~(t[42]);
  assign t[33] = t[53] ^ t[54];
  assign t[34] = t[41] ^ t[38];
  assign t[35] = ~(t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = ~(t[58] | t[59]);
  assign t[38] = t[60] ^ t[61];
  assign t[39] = t[62] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[63] ^ x[5];
  assign t[41] = t[64] ^ x[9];
  assign t[42] = t[65] ^ x[12];
  assign t[43] = t[66] ^ x[15];
  assign t[44] = t[67] ^ x[18];
  assign t[45] = t[68] ^ x[21];
  assign t[46] = t[69] ^ x[24];
  assign t[47] = t[70] ^ x[27];
  assign t[48] = t[71] ^ x[30];
  assign t[49] = t[72] ^ x[33];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[73] ^ x[36];
  assign t[51] = t[74] ^ x[39];
  assign t[52] = t[75] ^ x[42];
  assign t[53] = t[76] ^ x[45];
  assign t[54] = t[77] ^ x[48];
  assign t[55] = t[78] ^ x[51];
  assign t[56] = t[79] ^ x[54];
  assign t[57] = t[80] ^ x[57];
  assign t[58] = t[81] ^ x[60];
  assign t[59] = t[82] ^ x[63];
  assign t[5] = ~(t[9]);
  assign t[60] = t[83] ^ x[66];
  assign t[61] = t[84] ^ x[69];
  assign t[62] = (x[0] & x[1]);
  assign t[63] = (x[3] & x[4]);
  assign t[64] = (x[7] & x[8]);
  assign t[65] = (x[10] & x[11]);
  assign t[66] = (x[13] & x[14]);
  assign t[67] = (x[16] & x[17]);
  assign t[68] = (x[19] & x[20]);
  assign t[69] = (x[22] & x[23]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[25] & x[26]);
  assign t[71] = (x[28] & x[29]);
  assign t[72] = (x[31] & x[32]);
  assign t[73] = (x[34] & x[35]);
  assign t[74] = (x[37] & x[38]);
  assign t[75] = (x[40] & x[41]);
  assign t[76] = (x[43] & x[44]);
  assign t[77] = (x[46] & x[47]);
  assign t[78] = (x[49] & x[50]);
  assign t[79] = (x[52] & x[53]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[55] & x[56]);
  assign t[81] = (x[58] & x[59]);
  assign t[82] = (x[61] & x[62]);
  assign t[83] = (x[64] & x[65]);
  assign t[84] = (x[67] & x[68]);
  assign t[8] = t[12] ? t[13] : t[41];
  assign t[9] = t[42] & t[14];
  assign y = t[0] ? t[1] : t[39];
endmodule

module R1ind306(x, y);
 input [63:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[40]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[41] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[40] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[38] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[42] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[43] ^ t[33];
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[50] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[40]);
  assign t[33] = t[39] ^ t[52];
  assign t[34] = ~(t[53]);
  assign t[35] = ~(t[54] | t[55]);
  assign t[36] = ~(t[56] | t[57]);
  assign t[37] = t[58] ^ x[2];
  assign t[38] = t[59] ^ x[5];
  assign t[39] = t[60] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[61] ^ x[12];
  assign t[41] = t[62] ^ x[15];
  assign t[42] = t[63] ^ x[18];
  assign t[43] = t[64] ^ x[21];
  assign t[44] = t[65] ^ x[24];
  assign t[45] = t[66] ^ x[27];
  assign t[46] = t[67] ^ x[30];
  assign t[47] = t[68] ^ x[33];
  assign t[48] = t[69] ^ x[36];
  assign t[49] = t[70] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[71] ^ x[42];
  assign t[51] = t[72] ^ x[45];
  assign t[52] = t[73] ^ x[48];
  assign t[53] = t[74] ^ x[51];
  assign t[54] = t[75] ^ x[54];
  assign t[55] = t[76] ^ x[57];
  assign t[56] = t[77] ^ x[60];
  assign t[57] = t[78] ^ x[63];
  assign t[58] = (x[0] & x[1]);
  assign t[59] = (x[3] & x[4]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[7] & x[8]);
  assign t[61] = (x[10] & x[11]);
  assign t[62] = (x[13] & x[14]);
  assign t[63] = (x[16] & x[17]);
  assign t[64] = (x[19] & x[20]);
  assign t[65] = (x[22] & x[23]);
  assign t[66] = (x[25] & x[26]);
  assign t[67] = (x[28] & x[29]);
  assign t[68] = (x[31] & x[32]);
  assign t[69] = (x[34] & x[35]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[37] & x[38]);
  assign t[71] = (x[40] & x[41]);
  assign t[72] = (x[43] & x[44]);
  assign t[73] = (x[46] & x[47]);
  assign t[74] = (x[49] & x[50]);
  assign t[75] = (x[52] & x[53]);
  assign t[76] = (x[55] & x[56]);
  assign t[77] = (x[58] & x[59]);
  assign t[78] = (x[61] & x[62]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[39];
  assign t[9] = t[40] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind307(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind308(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind309(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind310(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind311(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind312(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind313(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind314(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind315(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind316(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind317(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind318(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind319(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind320(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind321(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind322(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind323(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind324(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind325(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind326(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind327(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind328(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind329(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind330(x, y);
 input [45:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[27]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[27] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[28] | t[20]);
  assign t[16] = ~(t[29] & t[30]);
  assign t[17] = ~(t[31] & t[32]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[33] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[35] | t[36]);
  assign t[23] = ~(t[37] | t[38]);
  assign t[24] = t[39] ^ x[2];
  assign t[25] = t[40] ^ x[5];
  assign t[26] = t[41] ^ x[9];
  assign t[27] = t[42] ^ x[12];
  assign t[28] = t[43] ^ x[15];
  assign t[29] = t[44] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[45] ^ x[21];
  assign t[31] = t[46] ^ x[24];
  assign t[32] = t[47] ^ x[27];
  assign t[33] = t[48] ^ x[30];
  assign t[34] = t[49] ^ x[33];
  assign t[35] = t[50] ^ x[36];
  assign t[36] = t[51] ^ x[39];
  assign t[37] = t[52] ^ x[42];
  assign t[38] = t[53] ^ x[45];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[3] & x[4]);
  assign t[41] = (x[7] & x[8]);
  assign t[42] = (x[10] & x[11]);
  assign t[43] = (x[13] & x[14]);
  assign t[44] = (x[16] & x[17]);
  assign t[45] = (x[19] & x[20]);
  assign t[46] = (x[22] & x[23]);
  assign t[47] = (x[25] & x[26]);
  assign t[48] = (x[28] & x[29]);
  assign t[49] = (x[31] & x[32]);
  assign t[4] = t[7] ? t[26] : x[6];
  assign t[50] = (x[34] & x[35]);
  assign t[51] = (x[37] & x[38]);
  assign t[52] = (x[40] & x[41]);
  assign t[53] = (x[43] & x[44]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[27] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind331(x, y);
 input [60:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[39] | t[15]);
  assign t[11] = ~(t[37]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[36] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = t[3] ? t[36] : t[4];
  assign t[20] = ~(t[29] | t[30]);
  assign t[21] = ~(t[40] | t[41]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[31] | t[32]);
  assign t[24] = ~(t[19]);
  assign t[25] = t[44] ^ t[33];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[51] & t[34]);
  assign t[31] = ~(t[52]);
  assign t[32] = ~(t[37]);
  assign t[33] = t[38] ^ t[53];
  assign t[34] = ~(t[54]);
  assign t[35] = t[55] ^ x[2];
  assign t[36] = t[56] ^ x[5];
  assign t[37] = t[57] ^ x[9];
  assign t[38] = t[58] ^ x[12];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[18];
  assign t[41] = t[61] ^ x[21];
  assign t[42] = t[62] ^ x[24];
  assign t[43] = t[63] ^ x[27];
  assign t[44] = t[64] ^ x[30];
  assign t[45] = t[65] ^ x[33];
  assign t[46] = t[66] ^ x[36];
  assign t[47] = t[67] ^ x[39];
  assign t[48] = t[68] ^ x[42];
  assign t[49] = t[69] ^ x[45];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[48];
  assign t[51] = t[71] ^ x[51];
  assign t[52] = t[72] ^ x[54];
  assign t[53] = t[73] ^ x[57];
  assign t[54] = t[74] ^ x[60];
  assign t[55] = (x[0] & x[1]);
  assign t[56] = (x[3] & x[4]);
  assign t[57] = (x[7] & x[8]);
  assign t[58] = (x[10] & x[11]);
  assign t[59] = (x[13] & x[14]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[16] & x[17]);
  assign t[61] = (x[19] & x[20]);
  assign t[62] = (x[22] & x[23]);
  assign t[63] = (x[25] & x[26]);
  assign t[64] = (x[28] & x[29]);
  assign t[65] = (x[31] & x[32]);
  assign t[66] = (x[34] & x[35]);
  assign t[67] = (x[37] & x[38]);
  assign t[68] = (x[40] & x[41]);
  assign t[69] = (x[43] & x[44]);
  assign t[6] = ~(t[37] & t[10]);
  assign t[70] = (x[46] & x[47]);
  assign t[71] = (x[49] & x[50]);
  assign t[72] = (x[52] & x[53]);
  assign t[73] = (x[55] & x[56]);
  assign t[74] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[37] & t[14];
  assign y = t[0] ? t[1] : t[35];
endmodule

module R1ind332(x, y);
 input [60:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[39] | t[15]);
  assign t[11] = ~(t[37]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[36] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = t[3] ? t[36] : t[4];
  assign t[20] = ~(t[29] | t[30]);
  assign t[21] = ~(t[40] | t[41]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[31] | t[32]);
  assign t[24] = ~(t[19]);
  assign t[25] = t[44] ^ t[33];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[51] & t[34]);
  assign t[31] = ~(t[52]);
  assign t[32] = ~(t[37]);
  assign t[33] = t[38] ^ t[53];
  assign t[34] = ~(t[54]);
  assign t[35] = t[55] ^ x[2];
  assign t[36] = t[56] ^ x[5];
  assign t[37] = t[57] ^ x[9];
  assign t[38] = t[58] ^ x[12];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[18];
  assign t[41] = t[61] ^ x[21];
  assign t[42] = t[62] ^ x[24];
  assign t[43] = t[63] ^ x[27];
  assign t[44] = t[64] ^ x[30];
  assign t[45] = t[65] ^ x[33];
  assign t[46] = t[66] ^ x[36];
  assign t[47] = t[67] ^ x[39];
  assign t[48] = t[68] ^ x[42];
  assign t[49] = t[69] ^ x[45];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[48];
  assign t[51] = t[71] ^ x[51];
  assign t[52] = t[72] ^ x[54];
  assign t[53] = t[73] ^ x[57];
  assign t[54] = t[74] ^ x[60];
  assign t[55] = (x[0] & x[1]);
  assign t[56] = (x[3] & x[4]);
  assign t[57] = (x[7] & x[8]);
  assign t[58] = (x[10] & x[11]);
  assign t[59] = (x[13] & x[14]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[16] & x[17]);
  assign t[61] = (x[19] & x[20]);
  assign t[62] = (x[22] & x[23]);
  assign t[63] = (x[25] & x[26]);
  assign t[64] = (x[28] & x[29]);
  assign t[65] = (x[31] & x[32]);
  assign t[66] = (x[34] & x[35]);
  assign t[67] = (x[37] & x[38]);
  assign t[68] = (x[40] & x[41]);
  assign t[69] = (x[43] & x[44]);
  assign t[6] = ~(t[37] & t[10]);
  assign t[70] = (x[46] & x[47]);
  assign t[71] = (x[49] & x[50]);
  assign t[72] = (x[52] & x[53]);
  assign t[73] = (x[55] & x[56]);
  assign t[74] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[37] & t[14];
  assign y = t[0] ? t[1] : t[35];
endmodule

module R1ind333(x, y);
 input [60:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[39] | t[15]);
  assign t[11] = ~(t[37]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[36] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = t[3] ? t[36] : t[4];
  assign t[20] = ~(t[29] | t[30]);
  assign t[21] = ~(t[40] | t[41]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[31] | t[32]);
  assign t[24] = ~(t[19]);
  assign t[25] = t[44] ^ t[33];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[51] & t[34]);
  assign t[31] = ~(t[52]);
  assign t[32] = ~(t[37]);
  assign t[33] = t[38] ^ t[53];
  assign t[34] = ~(t[54]);
  assign t[35] = t[55] ^ x[2];
  assign t[36] = t[56] ^ x[5];
  assign t[37] = t[57] ^ x[9];
  assign t[38] = t[58] ^ x[12];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[18];
  assign t[41] = t[61] ^ x[21];
  assign t[42] = t[62] ^ x[24];
  assign t[43] = t[63] ^ x[27];
  assign t[44] = t[64] ^ x[30];
  assign t[45] = t[65] ^ x[33];
  assign t[46] = t[66] ^ x[36];
  assign t[47] = t[67] ^ x[39];
  assign t[48] = t[68] ^ x[42];
  assign t[49] = t[69] ^ x[45];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[48];
  assign t[51] = t[71] ^ x[51];
  assign t[52] = t[72] ^ x[54];
  assign t[53] = t[73] ^ x[57];
  assign t[54] = t[74] ^ x[60];
  assign t[55] = (x[0] & x[1]);
  assign t[56] = (x[3] & x[4]);
  assign t[57] = (x[7] & x[8]);
  assign t[58] = (x[10] & x[11]);
  assign t[59] = (x[13] & x[14]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[16] & x[17]);
  assign t[61] = (x[19] & x[20]);
  assign t[62] = (x[22] & x[23]);
  assign t[63] = (x[25] & x[26]);
  assign t[64] = (x[28] & x[29]);
  assign t[65] = (x[31] & x[32]);
  assign t[66] = (x[34] & x[35]);
  assign t[67] = (x[37] & x[38]);
  assign t[68] = (x[40] & x[41]);
  assign t[69] = (x[43] & x[44]);
  assign t[6] = ~(t[37] & t[10]);
  assign t[70] = (x[46] & x[47]);
  assign t[71] = (x[49] & x[50]);
  assign t[72] = (x[52] & x[53]);
  assign t[73] = (x[55] & x[56]);
  assign t[74] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[37] & t[14];
  assign y = t[0] ? t[1] : t[35];
endmodule

module R1ind334(x, y);
 input [66:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[41] | t[15]);
  assign t[11] = ~(t[39]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[38] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = t[3] ? t[38] : t[4];
  assign t[20] = ~(t[29] | t[30]);
  assign t[21] = ~(t[42] | t[43]);
  assign t[22] = ~(t[44] | t[45]);
  assign t[23] = ~(t[31] | t[32]);
  assign t[24] = ~(t[19]);
  assign t[25] = t[33] ^ t[34];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[52] & t[35]);
  assign t[31] = ~(t[53]);
  assign t[32] = ~(t[39]);
  assign t[33] = t[54] ^ t[55];
  assign t[34] = t[40] ^ t[36];
  assign t[35] = ~(t[56]);
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ x[2];
  assign t[38] = t[60] ^ x[5];
  assign t[39] = t[61] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ x[12];
  assign t[41] = t[63] ^ x[15];
  assign t[42] = t[64] ^ x[18];
  assign t[43] = t[65] ^ x[21];
  assign t[44] = t[66] ^ x[24];
  assign t[45] = t[67] ^ x[27];
  assign t[46] = t[68] ^ x[30];
  assign t[47] = t[69] ^ x[33];
  assign t[48] = t[70] ^ x[36];
  assign t[49] = t[71] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[72] ^ x[42];
  assign t[51] = t[73] ^ x[45];
  assign t[52] = t[74] ^ x[48];
  assign t[53] = t[75] ^ x[51];
  assign t[54] = t[76] ^ x[54];
  assign t[55] = t[77] ^ x[57];
  assign t[56] = t[78] ^ x[60];
  assign t[57] = t[79] ^ x[63];
  assign t[58] = t[80] ^ x[66];
  assign t[59] = (x[0] & x[1]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[3] & x[4]);
  assign t[61] = (x[7] & x[8]);
  assign t[62] = (x[10] & x[11]);
  assign t[63] = (x[13] & x[14]);
  assign t[64] = (x[16] & x[17]);
  assign t[65] = (x[19] & x[20]);
  assign t[66] = (x[22] & x[23]);
  assign t[67] = (x[25] & x[26]);
  assign t[68] = (x[28] & x[29]);
  assign t[69] = (x[31] & x[32]);
  assign t[6] = ~(t[39] & t[10]);
  assign t[70] = (x[34] & x[35]);
  assign t[71] = (x[37] & x[38]);
  assign t[72] = (x[40] & x[41]);
  assign t[73] = (x[43] & x[44]);
  assign t[74] = (x[46] & x[47]);
  assign t[75] = (x[49] & x[50]);
  assign t[76] = (x[52] & x[53]);
  assign t[77] = (x[55] & x[56]);
  assign t[78] = (x[58] & x[59]);
  assign t[79] = (x[61] & x[62]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[64] & x[65]);
  assign t[8] = t[12] ? t[13] : t[40];
  assign t[9] = t[39] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind335(x, y);
 input [66:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[41] | t[15]);
  assign t[11] = ~(t[39]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[38] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = t[3] ? t[38] : t[4];
  assign t[20] = ~(t[29] | t[30]);
  assign t[21] = ~(t[42] | t[43]);
  assign t[22] = ~(t[44] | t[45]);
  assign t[23] = ~(t[31] | t[32]);
  assign t[24] = ~(t[19]);
  assign t[25] = t[33] ^ t[34];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[52] & t[35]);
  assign t[31] = ~(t[53]);
  assign t[32] = ~(t[39]);
  assign t[33] = t[54] ^ t[55];
  assign t[34] = t[40] ^ t[36];
  assign t[35] = ~(t[56]);
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ x[2];
  assign t[38] = t[60] ^ x[5];
  assign t[39] = t[61] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ x[12];
  assign t[41] = t[63] ^ x[15];
  assign t[42] = t[64] ^ x[18];
  assign t[43] = t[65] ^ x[21];
  assign t[44] = t[66] ^ x[24];
  assign t[45] = t[67] ^ x[27];
  assign t[46] = t[68] ^ x[30];
  assign t[47] = t[69] ^ x[33];
  assign t[48] = t[70] ^ x[36];
  assign t[49] = t[71] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[72] ^ x[42];
  assign t[51] = t[73] ^ x[45];
  assign t[52] = t[74] ^ x[48];
  assign t[53] = t[75] ^ x[51];
  assign t[54] = t[76] ^ x[54];
  assign t[55] = t[77] ^ x[57];
  assign t[56] = t[78] ^ x[60];
  assign t[57] = t[79] ^ x[63];
  assign t[58] = t[80] ^ x[66];
  assign t[59] = (x[0] & x[1]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[3] & x[4]);
  assign t[61] = (x[7] & x[8]);
  assign t[62] = (x[10] & x[11]);
  assign t[63] = (x[13] & x[14]);
  assign t[64] = (x[16] & x[17]);
  assign t[65] = (x[19] & x[20]);
  assign t[66] = (x[22] & x[23]);
  assign t[67] = (x[25] & x[26]);
  assign t[68] = (x[28] & x[29]);
  assign t[69] = (x[31] & x[32]);
  assign t[6] = ~(t[39] & t[10]);
  assign t[70] = (x[34] & x[35]);
  assign t[71] = (x[37] & x[38]);
  assign t[72] = (x[40] & x[41]);
  assign t[73] = (x[43] & x[44]);
  assign t[74] = (x[46] & x[47]);
  assign t[75] = (x[49] & x[50]);
  assign t[76] = (x[52] & x[53]);
  assign t[77] = (x[55] & x[56]);
  assign t[78] = (x[58] & x[59]);
  assign t[79] = (x[61] & x[62]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[64] & x[65]);
  assign t[8] = t[12] ? t[13] : t[40];
  assign t[9] = t[39] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind336(x, y);
 input [60:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[39] | t[15]);
  assign t[11] = ~(t[37]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[36] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = t[3] ? t[36] : t[4];
  assign t[20] = ~(t[29] | t[30]);
  assign t[21] = ~(t[40] | t[41]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[31] | t[32]);
  assign t[24] = ~(t[19]);
  assign t[25] = t[44] ^ t[33];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[51] & t[34]);
  assign t[31] = ~(t[52]);
  assign t[32] = ~(t[37]);
  assign t[33] = t[38] ^ t[53];
  assign t[34] = ~(t[54]);
  assign t[35] = t[55] ^ x[2];
  assign t[36] = t[56] ^ x[5];
  assign t[37] = t[57] ^ x[9];
  assign t[38] = t[58] ^ x[12];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[18];
  assign t[41] = t[61] ^ x[21];
  assign t[42] = t[62] ^ x[24];
  assign t[43] = t[63] ^ x[27];
  assign t[44] = t[64] ^ x[30];
  assign t[45] = t[65] ^ x[33];
  assign t[46] = t[66] ^ x[36];
  assign t[47] = t[67] ^ x[39];
  assign t[48] = t[68] ^ x[42];
  assign t[49] = t[69] ^ x[45];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[48];
  assign t[51] = t[71] ^ x[51];
  assign t[52] = t[72] ^ x[54];
  assign t[53] = t[73] ^ x[57];
  assign t[54] = t[74] ^ x[60];
  assign t[55] = (x[0] & x[1]);
  assign t[56] = (x[3] & x[4]);
  assign t[57] = (x[7] & x[8]);
  assign t[58] = (x[10] & x[11]);
  assign t[59] = (x[13] & x[14]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[16] & x[17]);
  assign t[61] = (x[19] & x[20]);
  assign t[62] = (x[22] & x[23]);
  assign t[63] = (x[25] & x[26]);
  assign t[64] = (x[28] & x[29]);
  assign t[65] = (x[31] & x[32]);
  assign t[66] = (x[34] & x[35]);
  assign t[67] = (x[37] & x[38]);
  assign t[68] = (x[40] & x[41]);
  assign t[69] = (x[43] & x[44]);
  assign t[6] = ~(t[37] & t[10]);
  assign t[70] = (x[46] & x[47]);
  assign t[71] = (x[49] & x[50]);
  assign t[72] = (x[52] & x[53]);
  assign t[73] = (x[55] & x[56]);
  assign t[74] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[37] & t[14];
  assign y = t[0] ? t[1] : t[35];
endmodule

module R1ind337(x, y);
 input [66:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[41] | t[15]);
  assign t[11] = ~(t[39]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[38] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = t[3] ? t[38] : t[4];
  assign t[20] = ~(t[29] | t[30]);
  assign t[21] = ~(t[42] | t[43]);
  assign t[22] = ~(t[44] | t[45]);
  assign t[23] = ~(t[31] | t[32]);
  assign t[24] = ~(t[19]);
  assign t[25] = t[33] ^ t[34];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[52] & t[35]);
  assign t[31] = ~(t[53]);
  assign t[32] = ~(t[39]);
  assign t[33] = t[54] ^ t[55];
  assign t[34] = t[40] ^ t[36];
  assign t[35] = ~(t[56]);
  assign t[36] = t[57] ^ t[58];
  assign t[37] = t[59] ^ x[2];
  assign t[38] = t[60] ^ x[5];
  assign t[39] = t[61] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ x[12];
  assign t[41] = t[63] ^ x[15];
  assign t[42] = t[64] ^ x[18];
  assign t[43] = t[65] ^ x[21];
  assign t[44] = t[66] ^ x[24];
  assign t[45] = t[67] ^ x[27];
  assign t[46] = t[68] ^ x[30];
  assign t[47] = t[69] ^ x[33];
  assign t[48] = t[70] ^ x[36];
  assign t[49] = t[71] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[72] ^ x[42];
  assign t[51] = t[73] ^ x[45];
  assign t[52] = t[74] ^ x[48];
  assign t[53] = t[75] ^ x[51];
  assign t[54] = t[76] ^ x[54];
  assign t[55] = t[77] ^ x[57];
  assign t[56] = t[78] ^ x[60];
  assign t[57] = t[79] ^ x[63];
  assign t[58] = t[80] ^ x[66];
  assign t[59] = (x[0] & x[1]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[3] & x[4]);
  assign t[61] = (x[7] & x[8]);
  assign t[62] = (x[10] & x[11]);
  assign t[63] = (x[13] & x[14]);
  assign t[64] = (x[16] & x[17]);
  assign t[65] = (x[19] & x[20]);
  assign t[66] = (x[22] & x[23]);
  assign t[67] = (x[25] & x[26]);
  assign t[68] = (x[28] & x[29]);
  assign t[69] = (x[31] & x[32]);
  assign t[6] = ~(t[39] & t[10]);
  assign t[70] = (x[34] & x[35]);
  assign t[71] = (x[37] & x[38]);
  assign t[72] = (x[40] & x[41]);
  assign t[73] = (x[43] & x[44]);
  assign t[74] = (x[46] & x[47]);
  assign t[75] = (x[49] & x[50]);
  assign t[76] = (x[52] & x[53]);
  assign t[77] = (x[55] & x[56]);
  assign t[78] = (x[58] & x[59]);
  assign t[79] = (x[61] & x[62]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[64] & x[65]);
  assign t[8] = t[12] ? t[13] : t[40];
  assign t[9] = t[39] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind338(x, y);
 input [60:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[39] | t[15]);
  assign t[11] = ~(t[37]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[36] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25] ^ t[26]);
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = t[3] ? t[36] : t[4];
  assign t[20] = ~(t[29] | t[30]);
  assign t[21] = ~(t[40] | t[41]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[31] | t[32]);
  assign t[24] = ~(t[19]);
  assign t[25] = t[44] ^ t[33];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[10]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[51] & t[34]);
  assign t[31] = ~(t[52]);
  assign t[32] = ~(t[37]);
  assign t[33] = t[38] ^ t[53];
  assign t[34] = ~(t[54]);
  assign t[35] = t[55] ^ x[2];
  assign t[36] = t[56] ^ x[5];
  assign t[37] = t[57] ^ x[9];
  assign t[38] = t[58] ^ x[12];
  assign t[39] = t[59] ^ x[15];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[18];
  assign t[41] = t[61] ^ x[21];
  assign t[42] = t[62] ^ x[24];
  assign t[43] = t[63] ^ x[27];
  assign t[44] = t[64] ^ x[30];
  assign t[45] = t[65] ^ x[33];
  assign t[46] = t[66] ^ x[36];
  assign t[47] = t[67] ^ x[39];
  assign t[48] = t[68] ^ x[42];
  assign t[49] = t[69] ^ x[45];
  assign t[4] = t[7] ? t[8] : x[6];
  assign t[50] = t[70] ^ x[48];
  assign t[51] = t[71] ^ x[51];
  assign t[52] = t[72] ^ x[54];
  assign t[53] = t[73] ^ x[57];
  assign t[54] = t[74] ^ x[60];
  assign t[55] = (x[0] & x[1]);
  assign t[56] = (x[3] & x[4]);
  assign t[57] = (x[7] & x[8]);
  assign t[58] = (x[10] & x[11]);
  assign t[59] = (x[13] & x[14]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[16] & x[17]);
  assign t[61] = (x[19] & x[20]);
  assign t[62] = (x[22] & x[23]);
  assign t[63] = (x[25] & x[26]);
  assign t[64] = (x[28] & x[29]);
  assign t[65] = (x[31] & x[32]);
  assign t[66] = (x[34] & x[35]);
  assign t[67] = (x[37] & x[38]);
  assign t[68] = (x[40] & x[41]);
  assign t[69] = (x[43] & x[44]);
  assign t[6] = ~(t[37] & t[10]);
  assign t[70] = (x[46] & x[47]);
  assign t[71] = (x[49] & x[50]);
  assign t[72] = (x[52] & x[53]);
  assign t[73] = (x[55] & x[56]);
  assign t[74] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[37] & t[14];
  assign y = t[0] ? t[1] : t[35];
endmodule

module R1ind339(x, y);
 input [42:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[9]);
  assign t[1] = t[3] ? t[23] : t[4];
  assign t[20] = ~(t[34] & t[21]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[36] ^ x[2];
  assign t[23] = t[37] ^ x[5];
  assign t[24] = t[38] ^ x[9];
  assign t[25] = t[39] ^ x[12];
  assign t[26] = t[40] ^ x[15];
  assign t[27] = t[41] ^ x[18];
  assign t[28] = t[42] ^ x[21];
  assign t[29] = t[43] ^ x[24];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[27];
  assign t[31] = t[45] ^ x[30];
  assign t[32] = t[46] ^ x[33];
  assign t[33] = t[47] ^ x[36];
  assign t[34] = t[48] ^ x[39];
  assign t[35] = t[49] ^ x[42];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[25] & x[26]);
  assign t[45] = (x[28] & x[29]);
  assign t[46] = (x[31] & x[32]);
  assign t[47] = (x[34] & x[35]);
  assign t[48] = (x[37] & x[38]);
  assign t[49] = (x[40] & x[41]);
  assign t[4] = t[7] ? t[23] : x[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[24] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[24] & t[11];
  assign t[9] = ~(t[25] | t[12]);
  assign y = t[0] ? t[1] : t[22];
endmodule

module R1ind340(x, y);
 input [42:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[9]);
  assign t[1] = t[3] ? t[23] : t[4];
  assign t[20] = ~(t[34] & t[21]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[36] ^ x[2];
  assign t[23] = t[37] ^ x[5];
  assign t[24] = t[38] ^ x[9];
  assign t[25] = t[39] ^ x[12];
  assign t[26] = t[40] ^ x[15];
  assign t[27] = t[41] ^ x[18];
  assign t[28] = t[42] ^ x[21];
  assign t[29] = t[43] ^ x[24];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[27];
  assign t[31] = t[45] ^ x[30];
  assign t[32] = t[46] ^ x[33];
  assign t[33] = t[47] ^ x[36];
  assign t[34] = t[48] ^ x[39];
  assign t[35] = t[49] ^ x[42];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[25] & x[26]);
  assign t[45] = (x[28] & x[29]);
  assign t[46] = (x[31] & x[32]);
  assign t[47] = (x[34] & x[35]);
  assign t[48] = (x[37] & x[38]);
  assign t[49] = (x[40] & x[41]);
  assign t[4] = t[7] ? t[23] : x[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[24] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[24] & t[11];
  assign t[9] = ~(t[25] | t[12]);
  assign y = t[0] ? t[1] : t[22];
endmodule

module R1ind341(x, y);
 input [42:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[9]);
  assign t[1] = t[3] ? t[23] : t[4];
  assign t[20] = ~(t[34] & t[21]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[36] ^ x[2];
  assign t[23] = t[37] ^ x[5];
  assign t[24] = t[38] ^ x[9];
  assign t[25] = t[39] ^ x[12];
  assign t[26] = t[40] ^ x[15];
  assign t[27] = t[41] ^ x[18];
  assign t[28] = t[42] ^ x[21];
  assign t[29] = t[43] ^ x[24];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[27];
  assign t[31] = t[45] ^ x[30];
  assign t[32] = t[46] ^ x[33];
  assign t[33] = t[47] ^ x[36];
  assign t[34] = t[48] ^ x[39];
  assign t[35] = t[49] ^ x[42];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[25] & x[26]);
  assign t[45] = (x[28] & x[29]);
  assign t[46] = (x[31] & x[32]);
  assign t[47] = (x[34] & x[35]);
  assign t[48] = (x[37] & x[38]);
  assign t[49] = (x[40] & x[41]);
  assign t[4] = t[7] ? t[23] : x[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[24] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[24] & t[11];
  assign t[9] = ~(t[25] | t[12]);
  assign y = t[0] ? t[1] : t[22];
endmodule

module R1ind342(x, y);
 input [42:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[9]);
  assign t[1] = t[3] ? t[23] : t[4];
  assign t[20] = ~(t[34] & t[21]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[36] ^ x[2];
  assign t[23] = t[37] ^ x[5];
  assign t[24] = t[38] ^ x[9];
  assign t[25] = t[39] ^ x[12];
  assign t[26] = t[40] ^ x[15];
  assign t[27] = t[41] ^ x[18];
  assign t[28] = t[42] ^ x[21];
  assign t[29] = t[43] ^ x[24];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[27];
  assign t[31] = t[45] ^ x[30];
  assign t[32] = t[46] ^ x[33];
  assign t[33] = t[47] ^ x[36];
  assign t[34] = t[48] ^ x[39];
  assign t[35] = t[49] ^ x[42];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[25] & x[26]);
  assign t[45] = (x[28] & x[29]);
  assign t[46] = (x[31] & x[32]);
  assign t[47] = (x[34] & x[35]);
  assign t[48] = (x[37] & x[38]);
  assign t[49] = (x[40] & x[41]);
  assign t[4] = t[7] ? t[23] : x[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[24] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[24] & t[11];
  assign t[9] = ~(t[25] | t[12]);
  assign y = t[0] ? t[1] : t[22];
endmodule

module R1ind343(x, y);
 input [42:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[9]);
  assign t[1] = t[3] ? t[23] : t[4];
  assign t[20] = ~(t[34] & t[21]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[36] ^ x[2];
  assign t[23] = t[37] ^ x[5];
  assign t[24] = t[38] ^ x[9];
  assign t[25] = t[39] ^ x[12];
  assign t[26] = t[40] ^ x[15];
  assign t[27] = t[41] ^ x[18];
  assign t[28] = t[42] ^ x[21];
  assign t[29] = t[43] ^ x[24];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[27];
  assign t[31] = t[45] ^ x[30];
  assign t[32] = t[46] ^ x[33];
  assign t[33] = t[47] ^ x[36];
  assign t[34] = t[48] ^ x[39];
  assign t[35] = t[49] ^ x[42];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[25] & x[26]);
  assign t[45] = (x[28] & x[29]);
  assign t[46] = (x[31] & x[32]);
  assign t[47] = (x[34] & x[35]);
  assign t[48] = (x[37] & x[38]);
  assign t[49] = (x[40] & x[41]);
  assign t[4] = t[7] ? t[23] : x[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[24] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[24] & t[11];
  assign t[9] = ~(t[25] | t[12]);
  assign y = t[0] ? t[1] : t[22];
endmodule

module R1ind344(x, y);
 input [42:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[9]);
  assign t[1] = t[3] ? t[23] : t[4];
  assign t[20] = ~(t[34] & t[21]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[36] ^ x[2];
  assign t[23] = t[37] ^ x[5];
  assign t[24] = t[38] ^ x[9];
  assign t[25] = t[39] ^ x[12];
  assign t[26] = t[40] ^ x[15];
  assign t[27] = t[41] ^ x[18];
  assign t[28] = t[42] ^ x[21];
  assign t[29] = t[43] ^ x[24];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[27];
  assign t[31] = t[45] ^ x[30];
  assign t[32] = t[46] ^ x[33];
  assign t[33] = t[47] ^ x[36];
  assign t[34] = t[48] ^ x[39];
  assign t[35] = t[49] ^ x[42];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[25] & x[26]);
  assign t[45] = (x[28] & x[29]);
  assign t[46] = (x[31] & x[32]);
  assign t[47] = (x[34] & x[35]);
  assign t[48] = (x[37] & x[38]);
  assign t[49] = (x[40] & x[41]);
  assign t[4] = t[7] ? t[23] : x[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[24] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[24] & t[11];
  assign t[9] = ~(t[25] | t[12]);
  assign y = t[0] ? t[1] : t[22];
endmodule

module R1ind345(x, y);
 input [42:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[9]);
  assign t[1] = t[3] ? t[23] : t[4];
  assign t[20] = ~(t[34] & t[21]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[36] ^ x[2];
  assign t[23] = t[37] ^ x[5];
  assign t[24] = t[38] ^ x[9];
  assign t[25] = t[39] ^ x[12];
  assign t[26] = t[40] ^ x[15];
  assign t[27] = t[41] ^ x[18];
  assign t[28] = t[42] ^ x[21];
  assign t[29] = t[43] ^ x[24];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[27];
  assign t[31] = t[45] ^ x[30];
  assign t[32] = t[46] ^ x[33];
  assign t[33] = t[47] ^ x[36];
  assign t[34] = t[48] ^ x[39];
  assign t[35] = t[49] ^ x[42];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[25] & x[26]);
  assign t[45] = (x[28] & x[29]);
  assign t[46] = (x[31] & x[32]);
  assign t[47] = (x[34] & x[35]);
  assign t[48] = (x[37] & x[38]);
  assign t[49] = (x[40] & x[41]);
  assign t[4] = t[7] ? t[23] : x[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[24] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[24] & t[11];
  assign t[9] = ~(t[25] | t[12]);
  assign y = t[0] ? t[1] : t[22];
endmodule

module R1ind346(x, y);
 input [42:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[24]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] | t[20]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[9]);
  assign t[1] = t[3] ? t[23] : t[4];
  assign t[20] = ~(t[34] & t[21]);
  assign t[21] = ~(t[35]);
  assign t[22] = t[36] ^ x[2];
  assign t[23] = t[37] ^ x[5];
  assign t[24] = t[38] ^ x[9];
  assign t[25] = t[39] ^ x[12];
  assign t[26] = t[40] ^ x[15];
  assign t[27] = t[41] ^ x[18];
  assign t[28] = t[42] ^ x[21];
  assign t[29] = t[43] ^ x[24];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[27];
  assign t[31] = t[45] ^ x[30];
  assign t[32] = t[46] ^ x[33];
  assign t[33] = t[47] ^ x[36];
  assign t[34] = t[48] ^ x[39];
  assign t[35] = t[49] ^ x[42];
  assign t[36] = (x[0] & x[1]);
  assign t[37] = (x[3] & x[4]);
  assign t[38] = (x[7] & x[8]);
  assign t[39] = (x[10] & x[11]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[13] & x[14]);
  assign t[41] = (x[16] & x[17]);
  assign t[42] = (x[19] & x[20]);
  assign t[43] = (x[22] & x[23]);
  assign t[44] = (x[25] & x[26]);
  assign t[45] = (x[28] & x[29]);
  assign t[46] = (x[31] & x[32]);
  assign t[47] = (x[34] & x[35]);
  assign t[48] = (x[37] & x[38]);
  assign t[49] = (x[40] & x[41]);
  assign t[4] = t[7] ? t[23] : x[6];
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[24] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[24] & t[11];
  assign t[9] = ~(t[25] | t[12]);
  assign y = t[0] ? t[1] : t[22];
endmodule

module R1ind347(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind348(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind349(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind350(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind351(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind352(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind353(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind354(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind355(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind356(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind357(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind358(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind359(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind360(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind361(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind362(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[25] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[5];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[3] & x[4]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[6];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind363(x, y);
 input [60:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[39]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[40] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[39] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[37] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[41] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[42] ^ t[33];
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[49] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[50]);
  assign t[32] = ~(t[39]);
  assign t[33] = t[38] ^ t[51];
  assign t[34] = ~(t[52]);
  assign t[35] = ~(t[53] | t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = t[57] ^ x[2];
  assign t[38] = t[58] ^ x[6];
  assign t[39] = t[59] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[12];
  assign t[41] = t[61] ^ x[15];
  assign t[42] = t[62] ^ x[18];
  assign t[43] = t[63] ^ x[21];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[27];
  assign t[46] = t[66] ^ x[30];
  assign t[47] = t[67] ^ x[33];
  assign t[48] = t[68] ^ x[36];
  assign t[49] = t[69] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[3];
  assign t[50] = t[70] ^ x[42];
  assign t[51] = t[71] ^ x[45];
  assign t[52] = t[72] ^ x[48];
  assign t[53] = t[73] ^ x[51];
  assign t[54] = t[74] ^ x[54];
  assign t[55] = t[75] ^ x[57];
  assign t[56] = t[76] ^ x[60];
  assign t[57] = (x[0] & x[1]);
  assign t[58] = (x[4] & x[5]);
  assign t[59] = (x[7] & x[8]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[10] & x[11]);
  assign t[61] = (x[13] & x[14]);
  assign t[62] = (x[16] & x[17]);
  assign t[63] = (x[19] & x[20]);
  assign t[64] = (x[22] & x[23]);
  assign t[65] = (x[25] & x[26]);
  assign t[66] = (x[28] & x[29]);
  assign t[67] = (x[31] & x[32]);
  assign t[68] = (x[34] & x[35]);
  assign t[69] = (x[37] & x[38]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[40] & x[41]);
  assign t[71] = (x[43] & x[44]);
  assign t[72] = (x[46] & x[47]);
  assign t[73] = (x[49] & x[50]);
  assign t[74] = (x[52] & x[53]);
  assign t[75] = (x[55] & x[56]);
  assign t[76] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[39] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind364(x, y);
 input [60:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[39]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[40] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[39] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[37] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[41] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[42] ^ t[33];
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[49] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[50]);
  assign t[32] = ~(t[39]);
  assign t[33] = t[38] ^ t[51];
  assign t[34] = ~(t[52]);
  assign t[35] = ~(t[53] | t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = t[57] ^ x[2];
  assign t[38] = t[58] ^ x[6];
  assign t[39] = t[59] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[12];
  assign t[41] = t[61] ^ x[15];
  assign t[42] = t[62] ^ x[18];
  assign t[43] = t[63] ^ x[21];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[27];
  assign t[46] = t[66] ^ x[30];
  assign t[47] = t[67] ^ x[33];
  assign t[48] = t[68] ^ x[36];
  assign t[49] = t[69] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[3];
  assign t[50] = t[70] ^ x[42];
  assign t[51] = t[71] ^ x[45];
  assign t[52] = t[72] ^ x[48];
  assign t[53] = t[73] ^ x[51];
  assign t[54] = t[74] ^ x[54];
  assign t[55] = t[75] ^ x[57];
  assign t[56] = t[76] ^ x[60];
  assign t[57] = (x[0] & x[1]);
  assign t[58] = (x[4] & x[5]);
  assign t[59] = (x[7] & x[8]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[10] & x[11]);
  assign t[61] = (x[13] & x[14]);
  assign t[62] = (x[16] & x[17]);
  assign t[63] = (x[19] & x[20]);
  assign t[64] = (x[22] & x[23]);
  assign t[65] = (x[25] & x[26]);
  assign t[66] = (x[28] & x[29]);
  assign t[67] = (x[31] & x[32]);
  assign t[68] = (x[34] & x[35]);
  assign t[69] = (x[37] & x[38]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[40] & x[41]);
  assign t[71] = (x[43] & x[44]);
  assign t[72] = (x[46] & x[47]);
  assign t[73] = (x[49] & x[50]);
  assign t[74] = (x[52] & x[53]);
  assign t[75] = (x[55] & x[56]);
  assign t[76] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[39] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind365(x, y);
 input [60:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[39]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[40] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[39] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[37] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[41] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[42] ^ t[33];
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[49] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[50]);
  assign t[32] = ~(t[39]);
  assign t[33] = t[38] ^ t[51];
  assign t[34] = ~(t[52]);
  assign t[35] = ~(t[53] | t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = t[57] ^ x[2];
  assign t[38] = t[58] ^ x[6];
  assign t[39] = t[59] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[12];
  assign t[41] = t[61] ^ x[15];
  assign t[42] = t[62] ^ x[18];
  assign t[43] = t[63] ^ x[21];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[27];
  assign t[46] = t[66] ^ x[30];
  assign t[47] = t[67] ^ x[33];
  assign t[48] = t[68] ^ x[36];
  assign t[49] = t[69] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[3];
  assign t[50] = t[70] ^ x[42];
  assign t[51] = t[71] ^ x[45];
  assign t[52] = t[72] ^ x[48];
  assign t[53] = t[73] ^ x[51];
  assign t[54] = t[74] ^ x[54];
  assign t[55] = t[75] ^ x[57];
  assign t[56] = t[76] ^ x[60];
  assign t[57] = (x[0] & x[1]);
  assign t[58] = (x[4] & x[5]);
  assign t[59] = (x[7] & x[8]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[10] & x[11]);
  assign t[61] = (x[13] & x[14]);
  assign t[62] = (x[16] & x[17]);
  assign t[63] = (x[19] & x[20]);
  assign t[64] = (x[22] & x[23]);
  assign t[65] = (x[25] & x[26]);
  assign t[66] = (x[28] & x[29]);
  assign t[67] = (x[31] & x[32]);
  assign t[68] = (x[34] & x[35]);
  assign t[69] = (x[37] & x[38]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[40] & x[41]);
  assign t[71] = (x[43] & x[44]);
  assign t[72] = (x[46] & x[47]);
  assign t[73] = (x[49] & x[50]);
  assign t[74] = (x[52] & x[53]);
  assign t[75] = (x[55] & x[56]);
  assign t[76] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[39] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind366(x, y);
 input [66:0] x;
 output y;

 wire [82:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[42] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[41] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[39] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[43] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[50] & t[35]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[36] & t[37]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[41]);
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[40] ^ t[38];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[61] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ x[6];
  assign t[41] = t[63] ^ x[9];
  assign t[42] = t[64] ^ x[12];
  assign t[43] = t[65] ^ x[15];
  assign t[44] = t[66] ^ x[18];
  assign t[45] = t[67] ^ x[21];
  assign t[46] = t[68] ^ x[24];
  assign t[47] = t[69] ^ x[27];
  assign t[48] = t[70] ^ x[30];
  assign t[49] = t[71] ^ x[33];
  assign t[4] = t[7] ? t[8] : x[3];
  assign t[50] = t[72] ^ x[36];
  assign t[51] = t[73] ^ x[39];
  assign t[52] = t[74] ^ x[42];
  assign t[53] = t[75] ^ x[45];
  assign t[54] = t[76] ^ x[48];
  assign t[55] = t[77] ^ x[51];
  assign t[56] = t[78] ^ x[54];
  assign t[57] = t[79] ^ x[57];
  assign t[58] = t[80] ^ x[60];
  assign t[59] = t[81] ^ x[63];
  assign t[5] = ~(t[9]);
  assign t[60] = t[82] ^ x[66];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[4] & x[5]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[58] & x[59]);
  assign t[81] = (x[61] & x[62]);
  assign t[82] = (x[64] & x[65]);
  assign t[8] = t[12] ? t[13] : t[40];
  assign t[9] = t[41] & t[14];
  assign y = t[0] ? t[1] : t[39];
endmodule

module R1ind367(x, y);
 input [66:0] x;
 output y;

 wire [82:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[42] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[41] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[39] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[43] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[50] & t[35]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[36] & t[37]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[41]);
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[40] ^ t[38];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[61] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ x[6];
  assign t[41] = t[63] ^ x[9];
  assign t[42] = t[64] ^ x[12];
  assign t[43] = t[65] ^ x[15];
  assign t[44] = t[66] ^ x[18];
  assign t[45] = t[67] ^ x[21];
  assign t[46] = t[68] ^ x[24];
  assign t[47] = t[69] ^ x[27];
  assign t[48] = t[70] ^ x[30];
  assign t[49] = t[71] ^ x[33];
  assign t[4] = t[7] ? t[8] : x[3];
  assign t[50] = t[72] ^ x[36];
  assign t[51] = t[73] ^ x[39];
  assign t[52] = t[74] ^ x[42];
  assign t[53] = t[75] ^ x[45];
  assign t[54] = t[76] ^ x[48];
  assign t[55] = t[77] ^ x[51];
  assign t[56] = t[78] ^ x[54];
  assign t[57] = t[79] ^ x[57];
  assign t[58] = t[80] ^ x[60];
  assign t[59] = t[81] ^ x[63];
  assign t[5] = ~(t[9]);
  assign t[60] = t[82] ^ x[66];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[4] & x[5]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[58] & x[59]);
  assign t[81] = (x[61] & x[62]);
  assign t[82] = (x[64] & x[65]);
  assign t[8] = t[12] ? t[13] : t[40];
  assign t[9] = t[41] & t[14];
  assign y = t[0] ? t[1] : t[39];
endmodule

module R1ind368(x, y);
 input [60:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[39]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[40] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[39] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[37] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[41] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[42] ^ t[33];
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[49] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[50]);
  assign t[32] = ~(t[39]);
  assign t[33] = t[38] ^ t[51];
  assign t[34] = ~(t[52]);
  assign t[35] = ~(t[53] | t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = t[57] ^ x[2];
  assign t[38] = t[58] ^ x[6];
  assign t[39] = t[59] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[12];
  assign t[41] = t[61] ^ x[15];
  assign t[42] = t[62] ^ x[18];
  assign t[43] = t[63] ^ x[21];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[27];
  assign t[46] = t[66] ^ x[30];
  assign t[47] = t[67] ^ x[33];
  assign t[48] = t[68] ^ x[36];
  assign t[49] = t[69] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[3];
  assign t[50] = t[70] ^ x[42];
  assign t[51] = t[71] ^ x[45];
  assign t[52] = t[72] ^ x[48];
  assign t[53] = t[73] ^ x[51];
  assign t[54] = t[74] ^ x[54];
  assign t[55] = t[75] ^ x[57];
  assign t[56] = t[76] ^ x[60];
  assign t[57] = (x[0] & x[1]);
  assign t[58] = (x[4] & x[5]);
  assign t[59] = (x[7] & x[8]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[10] & x[11]);
  assign t[61] = (x[13] & x[14]);
  assign t[62] = (x[16] & x[17]);
  assign t[63] = (x[19] & x[20]);
  assign t[64] = (x[22] & x[23]);
  assign t[65] = (x[25] & x[26]);
  assign t[66] = (x[28] & x[29]);
  assign t[67] = (x[31] & x[32]);
  assign t[68] = (x[34] & x[35]);
  assign t[69] = (x[37] & x[38]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[40] & x[41]);
  assign t[71] = (x[43] & x[44]);
  assign t[72] = (x[46] & x[47]);
  assign t[73] = (x[49] & x[50]);
  assign t[74] = (x[52] & x[53]);
  assign t[75] = (x[55] & x[56]);
  assign t[76] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[39] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind369(x, y);
 input [66:0] x;
 output y;

 wire [82:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[41]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[42] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[41] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[39] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[43] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[33] ^ t[34];
  assign t[25] = ~(t[44] ^ t[45]);
  assign t[26] = ~(t[46] & t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[50] & t[35]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[36] & t[37]);
  assign t[31] = ~(t[51]);
  assign t[32] = ~(t[41]);
  assign t[33] = t[52] ^ t[53];
  assign t[34] = t[40] ^ t[38];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = t[59] ^ t[60];
  assign t[39] = t[61] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[62] ^ x[6];
  assign t[41] = t[63] ^ x[9];
  assign t[42] = t[64] ^ x[12];
  assign t[43] = t[65] ^ x[15];
  assign t[44] = t[66] ^ x[18];
  assign t[45] = t[67] ^ x[21];
  assign t[46] = t[68] ^ x[24];
  assign t[47] = t[69] ^ x[27];
  assign t[48] = t[70] ^ x[30];
  assign t[49] = t[71] ^ x[33];
  assign t[4] = t[7] ? t[8] : x[3];
  assign t[50] = t[72] ^ x[36];
  assign t[51] = t[73] ^ x[39];
  assign t[52] = t[74] ^ x[42];
  assign t[53] = t[75] ^ x[45];
  assign t[54] = t[76] ^ x[48];
  assign t[55] = t[77] ^ x[51];
  assign t[56] = t[78] ^ x[54];
  assign t[57] = t[79] ^ x[57];
  assign t[58] = t[80] ^ x[60];
  assign t[59] = t[81] ^ x[63];
  assign t[5] = ~(t[9]);
  assign t[60] = t[82] ^ x[66];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[4] & x[5]);
  assign t[63] = (x[7] & x[8]);
  assign t[64] = (x[10] & x[11]);
  assign t[65] = (x[13] & x[14]);
  assign t[66] = (x[16] & x[17]);
  assign t[67] = (x[19] & x[20]);
  assign t[68] = (x[22] & x[23]);
  assign t[69] = (x[25] & x[26]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[28] & x[29]);
  assign t[71] = (x[31] & x[32]);
  assign t[72] = (x[34] & x[35]);
  assign t[73] = (x[37] & x[38]);
  assign t[74] = (x[40] & x[41]);
  assign t[75] = (x[43] & x[44]);
  assign t[76] = (x[46] & x[47]);
  assign t[77] = (x[49] & x[50]);
  assign t[78] = (x[52] & x[53]);
  assign t[79] = (x[55] & x[56]);
  assign t[7] = ~(t[11]);
  assign t[80] = (x[58] & x[59]);
  assign t[81] = (x[61] & x[62]);
  assign t[82] = (x[64] & x[65]);
  assign t[8] = t[12] ? t[13] : t[40];
  assign t[9] = t[41] & t[14];
  assign y = t[0] ? t[1] : t[39];
endmodule

module R1ind370(x, y);
 input [60:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[39]);
  assign t[12] = ~(t[16]);
  assign t[13] = t[17] ? t[40] : t[18];
  assign t[14] = t[19] & t[20];
  assign t[15] = ~(t[39] & t[21]);
  assign t[16] = ~(t[22]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24] ^ t[25]);
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = t[3] ? t[37] : t[4];
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[41] | t[30]);
  assign t[22] = ~(t[31] | t[32]);
  assign t[23] = ~(t[19]);
  assign t[24] = t[42] ^ t[33];
  assign t[25] = ~(t[43] ^ t[44]);
  assign t[26] = ~(t[45] & t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[21]);
  assign t[29] = ~(t[49] & t[34]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[35] & t[36]);
  assign t[31] = ~(t[50]);
  assign t[32] = ~(t[39]);
  assign t[33] = t[38] ^ t[51];
  assign t[34] = ~(t[52]);
  assign t[35] = ~(t[53] | t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = t[57] ^ x[2];
  assign t[38] = t[58] ^ x[6];
  assign t[39] = t[59] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[60] ^ x[12];
  assign t[41] = t[61] ^ x[15];
  assign t[42] = t[62] ^ x[18];
  assign t[43] = t[63] ^ x[21];
  assign t[44] = t[64] ^ x[24];
  assign t[45] = t[65] ^ x[27];
  assign t[46] = t[66] ^ x[30];
  assign t[47] = t[67] ^ x[33];
  assign t[48] = t[68] ^ x[36];
  assign t[49] = t[69] ^ x[39];
  assign t[4] = t[7] ? t[8] : x[3];
  assign t[50] = t[70] ^ x[42];
  assign t[51] = t[71] ^ x[45];
  assign t[52] = t[72] ^ x[48];
  assign t[53] = t[73] ^ x[51];
  assign t[54] = t[74] ^ x[54];
  assign t[55] = t[75] ^ x[57];
  assign t[56] = t[76] ^ x[60];
  assign t[57] = (x[0] & x[1]);
  assign t[58] = (x[4] & x[5]);
  assign t[59] = (x[7] & x[8]);
  assign t[5] = ~(t[9]);
  assign t[60] = (x[10] & x[11]);
  assign t[61] = (x[13] & x[14]);
  assign t[62] = (x[16] & x[17]);
  assign t[63] = (x[19] & x[20]);
  assign t[64] = (x[22] & x[23]);
  assign t[65] = (x[25] & x[26]);
  assign t[66] = (x[28] & x[29]);
  assign t[67] = (x[31] & x[32]);
  assign t[68] = (x[34] & x[35]);
  assign t[69] = (x[37] & x[38]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[40] & x[41]);
  assign t[71] = (x[43] & x[44]);
  assign t[72] = (x[46] & x[47]);
  assign t[73] = (x[49] & x[50]);
  assign t[74] = (x[52] & x[53]);
  assign t[75] = (x[55] & x[56]);
  assign t[76] = (x[58] & x[59]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ? t[13] : t[38];
  assign t[9] = t[39] & t[14];
  assign y = t[0] ? t[1] : t[37];
endmodule

module R1ind371(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind372(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind373(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind374(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind375(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind376(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind377(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind378(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind379(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind380(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind381(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind382(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind383(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind384(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind385(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind386(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind387(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind388(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind389(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind390(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind391(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind392(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind393(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind394(x, y);
 input [42:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[26]);
  assign t[11] = t[13] & t[14];
  assign t[12] = ~(t[26] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[27] | t[20]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[15]);
  assign t[19] = ~(t[32] & t[21]);
  assign t[1] = t[3] ? t[24] : t[4];
  assign t[20] = ~(t[22] & t[23]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = t[38] ^ x[2];
  assign t[25] = t[39] ^ x[6];
  assign t[26] = t[40] ^ x[9];
  assign t[27] = t[41] ^ x[12];
  assign t[28] = t[42] ^ x[15];
  assign t[29] = t[43] ^ x[18];
  assign t[2] = ~(t[5]);
  assign t[30] = t[44] ^ x[21];
  assign t[31] = t[45] ^ x[24];
  assign t[32] = t[46] ^ x[27];
  assign t[33] = t[47] ^ x[30];
  assign t[34] = t[48] ^ x[33];
  assign t[35] = t[49] ^ x[36];
  assign t[36] = t[50] ^ x[39];
  assign t[37] = t[51] ^ x[42];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[4] & x[5]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[7] & x[8]);
  assign t[41] = (x[10] & x[11]);
  assign t[42] = (x[13] & x[14]);
  assign t[43] = (x[16] & x[17]);
  assign t[44] = (x[19] & x[20]);
  assign t[45] = (x[22] & x[23]);
  assign t[46] = (x[25] & x[26]);
  assign t[47] = (x[28] & x[29]);
  assign t[48] = (x[31] & x[32]);
  assign t[49] = (x[34] & x[35]);
  assign t[4] = t[7] ? t[25] : x[3];
  assign t[50] = (x[37] & x[38]);
  assign t[51] = (x[40] & x[41]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = t[26] & t[11];
  assign t[9] = ~(t[12]);
  assign y = t[0] ? t[1] : t[24];
endmodule

module R1ind395(x, y);
 input [17:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[5] & t[1]);
  assign t[10] = t[16] ^ x[17];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[3] & x[4]);
  assign t[13] = (x[6] & x[7]);
  assign t[14] = (x[9] & x[10]);
  assign t[15] = (x[12] & x[13]);
  assign t[16] = (x[15] & x[16]);
  assign t[1] = ~(t[6] | t[2]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[4] = ~(t[9] | t[10]);
  assign t[5] = t[11] ^ x[2];
  assign t[6] = t[12] ^ x[5];
  assign t[7] = t[13] ^ x[8];
  assign t[8] = t[14] ^ x[11];
  assign t[9] = t[15] ^ x[14];
  assign y = ~(t[0]);
endmodule

module R1ind396(x, y);
 input [26:0] x;
 output y;

 wire [26:0] t;
  assign t[0] = ~(t[2] & t[9]);
  assign t[10] = t[19] ^ x[5];
  assign t[11] = t[20] ^ x[8];
  assign t[12] = t[21] ^ x[11];
  assign t[13] = t[22] ^ x[14];
  assign t[14] = t[23] ^ x[17];
  assign t[15] = t[24] ^ x[20];
  assign t[16] = t[25] ^ x[23];
  assign t[17] = t[26] ^ x[26];
  assign t[18] = (x[0] & x[1]);
  assign t[19] = (x[3] & x[4]);
  assign t[1] = ~(t[10] & t[3]);
  assign t[20] = (x[6] & x[7]);
  assign t[21] = (x[9] & x[10]);
  assign t[22] = (x[12] & x[13]);
  assign t[23] = (x[15] & x[16]);
  assign t[24] = (x[18] & x[19]);
  assign t[25] = (x[21] & x[22]);
  assign t[26] = (x[24] & x[25]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[11] | t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[12] | t[13]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[14] | t[15]);
  assign t[8] = ~(t[16] | t[17]);
  assign t[9] = t[18] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind397(x, y);
 input [35:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[21] & t[22]);
  assign t[11] = ~(t[23] & t[24]);
  assign t[12] = ~(t[5]);
  assign t[13] = ~(t[18] & t[16]);
  assign t[14] = ~(t[25] | t[26]);
  assign t[15] = ~(t[27] | t[28]);
  assign t[16] = ~(t[17]);
  assign t[17] = t[29] ^ x[2];
  assign t[18] = t[30] ^ x[5];
  assign t[19] = t[31] ^ x[8];
  assign t[1] = t[3] & t[18];
  assign t[20] = t[32] ^ x[11];
  assign t[21] = t[33] ^ x[14];
  assign t[22] = t[34] ^ x[17];
  assign t[23] = t[35] ^ x[20];
  assign t[24] = t[36] ^ x[23];
  assign t[25] = t[37] ^ x[26];
  assign t[26] = t[38] ^ x[29];
  assign t[27] = t[39] ^ x[32];
  assign t[28] = t[40] ^ x[35];
  assign t[29] = (x[0] & x[1]);
  assign t[2] = t[19] & t[4];
  assign t[30] = (x[3] & x[4]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[9] & x[10]);
  assign t[33] = (x[12] & x[13]);
  assign t[34] = (x[15] & x[16]);
  assign t[35] = (x[18] & x[19]);
  assign t[36] = (x[21] & x[22]);
  assign t[37] = (x[24] & x[25]);
  assign t[38] = (x[27] & x[28]);
  assign t[39] = (x[30] & x[31]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = (x[33] & x[34]);
  assign t[4] = t[7] & t[8];
  assign t[5] = ~(t[20] | t[9]);
  assign t[6] = ~(t[19]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[14] & t[15]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind398(x, y);
 input [35:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15] & t[16]);
  assign t[11] = ~(t[21] & t[22]);
  assign t[12] = ~(t[23] & t[24]);
  assign t[13] = ~(t[6]);
  assign t[14] = ~(t[17] & t[4]);
  assign t[15] = ~(t[25] | t[26]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = t[29] ^ x[2];
  assign t[18] = t[30] ^ x[5];
  assign t[19] = t[31] ^ x[8];
  assign t[1] = ~(t[3] & ~t[4]);
  assign t[20] = t[32] ^ x[11];
  assign t[21] = t[33] ^ x[14];
  assign t[22] = t[34] ^ x[17];
  assign t[23] = t[35] ^ x[20];
  assign t[24] = t[36] ^ x[23];
  assign t[25] = t[37] ^ x[26];
  assign t[26] = t[38] ^ x[29];
  assign t[27] = t[39] ^ x[32];
  assign t[28] = t[40] ^ x[35];
  assign t[29] = (x[0] & x[1]);
  assign t[2] = t[18] & t[5];
  assign t[30] = (x[3] & x[4]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[9] & x[10]);
  assign t[33] = (x[12] & x[13]);
  assign t[34] = (x[15] & x[16]);
  assign t[35] = (x[18] & x[19]);
  assign t[36] = (x[21] & x[22]);
  assign t[37] = (x[24] & x[25]);
  assign t[38] = (x[27] & x[28]);
  assign t[39] = (x[30] & x[31]);
  assign t[3] = ~(t[6] | t[7]);
  assign t[40] = (x[33] & x[34]);
  assign t[4] = ~(t[19]);
  assign t[5] = t[8] & t[9];
  assign t[6] = ~(t[20] | t[10]);
  assign t[7] = ~(t[18]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[13] | t[14]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind399(x, y);
 input [35:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[23] | t[12]);
  assign t[11] = ~(t[24]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[25] | t[17]);
  assign t[14] = ~(t[26] | t[15]);
  assign t[15] = t[27] ^ x[2];
  assign t[16] = t[28] ^ x[5];
  assign t[17] = t[29] ^ x[8];
  assign t[18] = t[30] ^ x[11];
  assign t[19] = t[31] ^ x[14];
  assign t[1] = ~(t[16] & ~t[17]);
  assign t[20] = t[32] ^ x[17];
  assign t[21] = t[33] ^ x[20];
  assign t[22] = t[34] ^ x[23];
  assign t[23] = t[35] ^ x[26];
  assign t[24] = t[36] ^ x[29];
  assign t[25] = t[37] ^ x[32];
  assign t[26] = t[38] ^ x[35];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[3] & x[4]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = t[16] & t[3];
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[21] & x[22]);
  assign t[35] = (x[24] & x[25]);
  assign t[36] = (x[27] & x[28]);
  assign t[37] = (x[30] & x[31]);
  assign t[38] = (x[33] & x[34]);
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = ~(t[10]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind400(x, y);
 input [35:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[23] | t[12]);
  assign t[11] = ~(t[24]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[25] | t[15]);
  assign t[14] = ~(t[17] | t[26]);
  assign t[15] = t[27] ^ x[2];
  assign t[16] = t[28] ^ x[5];
  assign t[17] = t[29] ^ x[8];
  assign t[18] = t[30] ^ x[11];
  assign t[19] = t[31] ^ x[14];
  assign t[1] = t[16] & t[17];
  assign t[20] = t[32] ^ x[17];
  assign t[21] = t[33] ^ x[20];
  assign t[22] = t[34] ^ x[23];
  assign t[23] = t[35] ^ x[26];
  assign t[24] = t[36] ^ x[29];
  assign t[25] = t[37] ^ x[32];
  assign t[26] = t[38] ^ x[35];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[3] & x[4]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = t[16] & t[3];
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[21] & x[22]);
  assign t[35] = (x[24] & x[25]);
  assign t[36] = (x[27] & x[28]);
  assign t[37] = (x[30] & x[31]);
  assign t[38] = (x[33] & x[34]);
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = ~(t[10]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind401(x, y);
 input [35:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[17] | t[12]);
  assign t[11] = ~(t[23]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[24] | t[25]);
  assign t[14] = ~(t[15] | t[26]);
  assign t[15] = t[27] ^ x[2];
  assign t[16] = t[28] ^ x[5];
  assign t[17] = t[29] ^ x[8];
  assign t[18] = t[30] ^ x[11];
  assign t[19] = t[31] ^ x[14];
  assign t[1] = ~(t[16] & ~t[17]);
  assign t[20] = t[32] ^ x[17];
  assign t[21] = t[33] ^ x[20];
  assign t[22] = t[34] ^ x[23];
  assign t[23] = t[35] ^ x[26];
  assign t[24] = t[36] ^ x[29];
  assign t[25] = t[37] ^ x[32];
  assign t[26] = t[38] ^ x[35];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[3] & x[4]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = t[16] & t[3];
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[21] & x[22]);
  assign t[35] = (x[24] & x[25]);
  assign t[36] = (x[27] & x[28]);
  assign t[37] = (x[30] & x[31]);
  assign t[38] = (x[33] & x[34]);
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = ~(t[10]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind402(x, y);
 input [35:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[15] | t[12]);
  assign t[11] = ~(t[23]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[17] | t[24]);
  assign t[14] = ~(t[25] | t[26]);
  assign t[15] = t[27] ^ x[2];
  assign t[16] = t[28] ^ x[5];
  assign t[17] = t[29] ^ x[8];
  assign t[18] = t[30] ^ x[11];
  assign t[19] = t[31] ^ x[14];
  assign t[1] = t[16] & t[17];
  assign t[20] = t[32] ^ x[17];
  assign t[21] = t[33] ^ x[20];
  assign t[22] = t[34] ^ x[23];
  assign t[23] = t[35] ^ x[26];
  assign t[24] = t[36] ^ x[29];
  assign t[25] = t[37] ^ x[32];
  assign t[26] = t[38] ^ x[35];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[3] & x[4]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = t[16] & t[3];
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[21] & x[22]);
  assign t[35] = (x[24] & x[25]);
  assign t[36] = (x[27] & x[28]);
  assign t[37] = (x[30] & x[31]);
  assign t[38] = (x[33] & x[34]);
  assign t[3] = t[4] & t[5];
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = ~(t[10]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind403(x, y);
 input [35:0] x;
 output y;

 wire [39:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[24] | t[13]);
  assign t[12] = ~(t[25]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[16] | t[26]);
  assign t[15] = ~(t[27] | t[18]);
  assign t[16] = t[28] ^ x[2];
  assign t[17] = t[29] ^ x[5];
  assign t[18] = t[30] ^ x[8];
  assign t[19] = t[31] ^ x[11];
  assign t[1] = ~(t[17] & ~t[3]);
  assign t[20] = t[32] ^ x[14];
  assign t[21] = t[33] ^ x[17];
  assign t[22] = t[34] ^ x[20];
  assign t[23] = t[35] ^ x[23];
  assign t[24] = t[36] ^ x[26];
  assign t[25] = t[37] ^ x[29];
  assign t[26] = t[38] ^ x[32];
  assign t[27] = t[39] ^ x[35];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[3] & x[4]);
  assign t[2] = t[17] & t[4];
  assign t[30] = (x[6] & x[7]);
  assign t[31] = (x[9] & x[10]);
  assign t[32] = (x[12] & x[13]);
  assign t[33] = (x[15] & x[16]);
  assign t[34] = (x[18] & x[19]);
  assign t[35] = (x[21] & x[22]);
  assign t[36] = (x[24] & x[25]);
  assign t[37] = (x[27] & x[28]);
  assign t[38] = (x[30] & x[31]);
  assign t[39] = (x[33] & x[34]);
  assign t[3] = ~(t[18] ^ t[16]);
  assign t[4] = t[5] & t[6];
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[9] = ~(t[11]);
  assign y = t[0] ? t[1] : t[16];
endmodule

module R1_ind(x, y);
 input [1081:0] x;
 output [403:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[8], x[7], x[6]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[11], x[10], x[9]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[14], x[13], x[12]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[17], x[16], x[15]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[20], x[19], x[18]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[23], x[22], x[21]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[26], x[25], x[24]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[29], x[28], x[27]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[32], x[31], x[30]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[35], x[34], x[33]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[38], x[37], x[36]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[41], x[40], x[39]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[44], x[43], x[42]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[47], x[46], x[45]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[50], x[49], x[48]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[53], x[52], x[51]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[56], x[55], x[54]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[59], x[58], x[57]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[62], x[61], x[60]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[65], x[64], x[63]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[68], x[67], x[66]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[71], x[70], x[69]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[74], x[73], x[72]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[77], x[76], x[75]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[80], x[79], x[78]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[83], x[82], x[81]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[86], x[85], x[84]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[89], x[88], x[87]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[92], x[91], x[90]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[95], x[94], x[93]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[98], x[97], x[96]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[101], x[100], x[99]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[104], x[103], x[102]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[107], x[106], x[105]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[110], x[109], x[108]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[113], x[112], x[111]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[116], x[115], x[114]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[119], x[118], x[117]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[122], x[121], x[120]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[125], x[124], x[123]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[128], x[127], x[126]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[131], x[130], x[129]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[134], x[133], x[132]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[137], x[136], x[135]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[140], x[139], x[138]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[143], x[142], x[141]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[146], x[145], x[144]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[149], x[148], x[147]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[152], x[151], x[150]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[155], x[154], x[153]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[158], x[157], x[156]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[161], x[160], x[159]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[164], x[163], x[162]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[167], x[166], x[165]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[170], x[169], x[168]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[173], x[172], x[171]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[176], x[175], x[174]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[179], x[178], x[177]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[182], x[181], x[180]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[185], x[184], x[183]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[188], x[187], x[186]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[191], x[190], x[189]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[194], x[193], x[192]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[197], x[196], x[195]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[200], x[199], x[198]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[203], x[202], x[201]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[206], x[205], x[204]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[209], x[208], x[207]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[212], x[211], x[210]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[215], x[214], x[213]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[218], x[217], x[216]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[221], x[220], x[219]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[224], x[223], x[222]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[227], x[226], x[225]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[230], x[229], x[228]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[233], x[232], x[231]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[236], x[235], x[234]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[239], x[238], x[237]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[242], x[241], x[240]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[245], x[244], x[243]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[248], x[247], x[246]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[251], x[250], x[249]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[254], x[253], x[252]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[257], x[256], x[255]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[260], x[259], x[258]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[263], x[262], x[261]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[266], x[265], x[264]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[269], x[268], x[267]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[272], x[271], x[270]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[275], x[274], x[273]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[278], x[277], x[276]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[281], x[280], x[279]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[284], x[283], x[282]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[287], x[286], x[285]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[290], x[289], x[288]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[293], x[292], x[291]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[296], x[295], x[294]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[299], x[298], x[297]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[302], x[301], x[300]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[305], x[304], x[303]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[308], x[307], x[306]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[311], x[310], x[309]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[314], x[313], x[312]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[317], x[316], x[315]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[320], x[319], x[318]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[323], x[322], x[321]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[326], x[325], x[324]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[329], x[328], x[327]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[332], x[331], x[330]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[335], x[334], x[333]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[338], x[337], x[336]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[341], x[340], x[339]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[344], x[343], x[342]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[347], x[346], x[345]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[350], x[349], x[348]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[353], x[352], x[351]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[356], x[355], x[354]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[359], x[358], x[357]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[362], x[361], x[360]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[365], x[364], x[363]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[368], x[367], x[366]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[371], x[370], x[369]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[374], x[373], x[372]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[377], x[376], x[375]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[380], x[379], x[378]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[383], x[382], x[381]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[386], x[385], x[384]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[389], x[388], x[387]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x(x[423]), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[429], x[428], x[427], x[426], x[425], x[424], x[389], x[388], x[387]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[395], x[394], x[393], x[426], x[425], x[424]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[398], x[397], x[396], x[395], x[394], x[393]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[429], x[428], x[427], x[432], x[431], x[430], x[398], x[397], x[396]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[432], x[431], x[430], x[401], x[400], x[399], x[429], x[428], x[427], x[389], x[388], x[387]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[398], x[397], x[396], x[395], x[394], x[393], x[407], x[406], x[405], x[401], x[400], x[399], x[392], x[391], x[390], x[389], x[388], x[387]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[407], x[406], x[405], x[389], x[388], x[387], x[429], x[428], x[427], x[435], x[434], x[433], x[392], x[391], x[390]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[435], x[434], x[433], x[429], x[428], x[427], x[389], x[388], x[387]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[458], x[457], x[456], x[455], x[454], x[453], x[452], x[451], x[450], x[449]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[468], x[467], x[466], x[465], x[464], x[463], x[462], x[461], x[460], x[459]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[478], x[477], x[476], x[475], x[474], x[473], x[472], x[471], x[470], x[469]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[488], x[487], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[479]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[498], x[497], x[496], x[495], x[494], x[493], x[492], x[491], x[490], x[489]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[508], x[507], x[506], x[505], x[504], x[503], x[502], x[501], x[500], x[499]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[518], x[517], x[516], x[515], x[514], x[513], x[512], x[511], x[510], x[509]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[438], x[437], x[436], x[525], x[524], x[523], x[522], x[521], x[520], x[519]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[451], x[450], x[449], x[532], x[531], x[530], x[529], x[528], x[527], x[526]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[461], x[460], x[459], x[539], x[538], x[537], x[536], x[535], x[534], x[533]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[471], x[470], x[469], x[546], x[545], x[544], x[543], x[542], x[541], x[540]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[481], x[480], x[479], x[553], x[552], x[551], x[550], x[549], x[548], x[547]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[491], x[490], x[489], x[560], x[559], x[558], x[557], x[556], x[555], x[554]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[501], x[500], x[499], x[567], x[566], x[565], x[564], x[563], x[562], x[561]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[511], x[510], x[509], x[574], x[573], x[572], x[571], x[570], x[569], x[568]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[521], x[520], x[519], x[581], x[580], x[579], x[578], x[577], x[576], x[575]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[528], x[527], x[526], x[588], x[587], x[586], x[585], x[584], x[583], x[582]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[535], x[534], x[533], x[595], x[594], x[593], x[592], x[591], x[590], x[589]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[542], x[541], x[540], x[602], x[601], x[600], x[599], x[598], x[597], x[596]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[549], x[548], x[547], x[609], x[608], x[607], x[606], x[605], x[604], x[603]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[556], x[555], x[554], x[616], x[615], x[614], x[613], x[612], x[611], x[610]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[563], x[562], x[561], x[623], x[622], x[621], x[620], x[619], x[618], x[617]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[570], x[569], x[568], x[630], x[629], x[628], x[627], x[626], x[625], x[624]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[458], x[457], x[456], x[23], x[22], x[21], x[518], x[517], x[516], x[5], x[4], x[3], x[468], x[467], x[466], x[20], x[19], x[18], x[508], x[507], x[506], x[8], x[7], x[6], x[488], x[487], x[486], x[14], x[13], x[12], x[661], x[660], x[659], x[658], x[657], x[656], x[26], x[25], x[24], x[655], x[654], x[653], x[652], x[651], x[650], x[649], x[648], x[647], x[646], x[645], x[644], x[498], x[497], x[496], x[11], x[10], x[9], x[478], x[477], x[476], x[17], x[16], x[15], x[643], x[642], x[641], x[640], x[639], x[638], x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[637], x[636], x[635], x[429], x[428], x[427], x[448], x[447], x[446], x[389], x[388], x[387], x[445], x[444], x[443], x[577], x[576], x[575], x[634], x[633], x[632], x[631]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[488], x[487], x[486], x[14], x[13], x[12], x[518], x[517], x[516], x[5], x[4], x[3], x[508], x[507], x[506], x[8], x[7], x[6], x[468], x[467], x[466], x[20], x[19], x[18], x[23], x[22], x[21], x[649], x[648], x[647], x[478], x[477], x[476], x[17], x[16], x[15], x[658], x[657], x[656], x[652], x[651], x[650], x[655], x[654], x[653], x[661], x[660], x[659], x[498], x[497], x[496], x[11], x[10], x[9], x[445], x[444], x[443], x[26], x[25], x[24], x[640], x[639], x[638], x[643], x[642], x[641], x[646], x[645], x[644], x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[637], x[636], x[635], x[426], x[425], x[424], x[448], x[447], x[446], x[389], x[388], x[387], x[458], x[457], x[456], x[584], x[583], x[582], x[665], x[664], x[663], x[662]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[488], x[487], x[486], x[14], x[13], x[12], x[20], x[19], x[18], x[458], x[457], x[456], x[23], x[22], x[21], x[478], x[477], x[476], x[17], x[16], x[15], x[649], x[648], x[647], x[518], x[517], x[516], x[5], x[4], x[3], x[508], x[507], x[506], x[8], x[7], x[6], x[655], x[654], x[653], x[661], x[660], x[659], x[640], x[639], x[638], x[658], x[657], x[656], x[652], x[651], x[650], x[498], x[497], x[496], x[11], x[10], x[9], x[445], x[444], x[443], x[26], x[25], x[24], x[643], x[642], x[641], x[646], x[645], x[644], x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[637], x[636], x[635], x[395], x[394], x[393], x[389], x[388], x[387], x[468], x[467], x[466], x[591], x[590], x[589], x[669], x[668], x[667], x[666]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[458], x[457], x[456], x[23], x[22], x[21], x[468], x[467], x[466], x[20], x[19], x[18], x[508], x[507], x[506], x[8], x[7], x[6], x[488], x[487], x[486], x[14], x[13], x[12], x[661], x[660], x[659], x[518], x[517], x[516], x[5], x[4], x[3], x[445], x[444], x[443], x[26], x[25], x[24], x[655], x[654], x[653], x[652], x[651], x[650], x[649], x[648], x[647], x[658], x[657], x[656], x[646], x[645], x[644], x[498], x[497], x[496], x[11], x[10], x[9], x[17], x[16], x[15], x[643], x[642], x[641], x[640], x[639], x[638], x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[637], x[636], x[635], x[398], x[397], x[396], x[389], x[388], x[387], x[478], x[477], x[476], x[598], x[597], x[596], x[673], x[672], x[671], x[670]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[14], x[13], x[12], x[508], x[507], x[506], x[8], x[7], x[6], x[649], x[648], x[647], x[468], x[467], x[466], x[20], x[19], x[18], x[458], x[457], x[456], x[23], x[22], x[21], x[652], x[651], x[650], x[655], x[654], x[653], x[661], x[660], x[659], x[498], x[497], x[496], x[11], x[10], x[9], x[478], x[477], x[476], x[17], x[16], x[15], x[445], x[444], x[443], x[26], x[25], x[24], x[518], x[517], x[516], x[5], x[4], x[3], x[643], x[642], x[641], x[640], x[639], x[638], x[646], x[645], x[644], x[658], x[657], x[656], x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[637], x[636], x[635], x[432], x[431], x[430], x[448], x[447], x[446], x[389], x[388], x[387], x[488], x[487], x[486], x[605], x[604], x[603], x[677], x[676], x[675], x[674]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[488], x[487], x[486], x[14], x[13], x[12], x[458], x[457], x[456], x[23], x[22], x[21], x[508], x[507], x[506], x[8], x[7], x[6], x[468], x[467], x[466], x[20], x[19], x[18], x[445], x[444], x[443], x[26], x[25], x[24], x[649], x[648], x[647], x[661], x[660], x[659], x[518], x[517], x[516], x[5], x[4], x[3], x[652], x[651], x[650], x[655], x[654], x[653], x[646], x[645], x[644], x[11], x[10], x[9], x[478], x[477], x[476], x[17], x[16], x[15], x[658], x[657], x[656], x[643], x[642], x[641], x[640], x[639], x[638], x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[637], x[636], x[635], x[401], x[400], x[399], x[448], x[447], x[446], x[389], x[388], x[387], x[498], x[497], x[496], x[612], x[611], x[610], x[681], x[680], x[679], x[678]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[488], x[487], x[486], x[14], x[13], x[12], x[8], x[7], x[6], x[649], x[648], x[647], x[652], x[651], x[650], x[498], x[497], x[496], x[11], x[10], x[9], x[478], x[477], x[476], x[17], x[16], x[15], x[445], x[444], x[443], x[26], x[25], x[24], x[468], x[467], x[466], x[20], x[19], x[18], x[458], x[457], x[456], x[23], x[22], x[21], x[643], x[642], x[641], x[640], x[639], x[638], x[646], x[645], x[644], x[655], x[654], x[653], x[661], x[660], x[659], x[518], x[517], x[516], x[5], x[4], x[3], x[658], x[657], x[656], x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[407], x[406], x[405], x[637], x[636], x[635], x[392], x[391], x[390], x[448], x[447], x[446], x[389], x[388], x[387], x[508], x[507], x[506], x[619], x[618], x[617], x[685], x[684], x[683], x[682]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[458], x[457], x[456], x[23], x[22], x[21], x[661], x[660], x[659], x[468], x[467], x[466], x[20], x[19], x[18], x[488], x[487], x[486], x[14], x[13], x[12], x[508], x[507], x[506], x[8], x[7], x[6], x[445], x[444], x[443], x[26], x[25], x[24], x[655], x[654], x[653], x[649], x[648], x[647], x[5], x[4], x[3], x[652], x[651], x[650], x[646], x[645], x[644], x[498], x[497], x[496], x[11], x[10], x[9], x[478], x[477], x[476], x[17], x[16], x[15], x[658], x[657], x[656], x[643], x[642], x[641], x[640], x[639], x[638], x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[637], x[636], x[635], x[435], x[434], x[433], x[448], x[447], x[446], x[389], x[388], x[387], x[518], x[517], x[516], x[626], x[625], x[624], x[689], x[688], x[687], x[686]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[633], x[632], x[631], x[693], x[438], x[437], x[436], x[692], x[691], x[690]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[664], x[663], x[662], x[697], x[451], x[450], x[449], x[696], x[695], x[694]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[668], x[667], x[666], x[701], x[461], x[460], x[459], x[700], x[699], x[698]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[672], x[671], x[670], x[705], x[471], x[470], x[469], x[704], x[703], x[702]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[676], x[675], x[674], x[709], x[481], x[480], x[479], x[708], x[707], x[706]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[680], x[679], x[678], x[713], x[491], x[490], x[489], x[712], x[711], x[710]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[684], x[683], x[682], x[717], x[501], x[500], x[499], x[716], x[715], x[714]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[688], x[687], x[686], x[721], x[511], x[510], x[509], x[720], x[719], x[718]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[692], x[691], x[690], x[725], x[521], x[520], x[519], x[724], x[723], x[722]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[696], x[695], x[694], x[729], x[528], x[527], x[526], x[728], x[727], x[726]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[700], x[699], x[698], x[733], x[535], x[534], x[533], x[732], x[731], x[730]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[704], x[703], x[702], x[737], x[542], x[541], x[540], x[736], x[735], x[734]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[708], x[707], x[706], x[741], x[549], x[548], x[547], x[740], x[739], x[738]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[712], x[711], x[710], x[745], x[556], x[555], x[554], x[744], x[743], x[742]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[716], x[715], x[714], x[749], x[563], x[562], x[561], x[748], x[747], x[746]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[720], x[719], x[718], x[753], x[570], x[569], x[568], x[752], x[751], x[750]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[724], x[723], x[722], x[757], x[577], x[576], x[575], x[756], x[755], x[754]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[728], x[727], x[726], x[761], x[584], x[583], x[582], x[760], x[759], x[758]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[732], x[731], x[730], x[765], x[591], x[590], x[589], x[764], x[763], x[762]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[736], x[735], x[734], x[769], x[598], x[597], x[596], x[768], x[767], x[766]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[740], x[739], x[738], x[773], x[605], x[604], x[603], x[772], x[771], x[770]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[744], x[743], x[742], x[777], x[612], x[611], x[610], x[776], x[775], x[774]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[748], x[747], x[746], x[781], x[619], x[618], x[617], x[780], x[779], x[778]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[752], x[751], x[750], x[785], x[626], x[625], x[624], x[784], x[783], x[782]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[756], x[755], x[754], x[789], x[633], x[632], x[631], x[788], x[787], x[786]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[760], x[759], x[758], x[793], x[664], x[663], x[662], x[792], x[791], x[790]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[764], x[763], x[762], x[797], x[668], x[667], x[666], x[796], x[795], x[794]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[768], x[767], x[766], x[801], x[672], x[671], x[670], x[800], x[799], x[798]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[772], x[771], x[770], x[805], x[676], x[675], x[674], x[804], x[803], x[802]}), .y(y[199]));
  R1ind200 R1ind200_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[776], x[775], x[774], x[809], x[680], x[679], x[678], x[808], x[807], x[806]}), .y(y[200]));
  R1ind201 R1ind201_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[780], x[779], x[778], x[813], x[684], x[683], x[682], x[812], x[811], x[810]}), .y(y[201]));
  R1ind202 R1ind202_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[784], x[783], x[782], x[817], x[688], x[687], x[686], x[816], x[815], x[814]}), .y(y[202]));
  R1ind203 R1ind203_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[788], x[787], x[786], x[818], x[692], x[691], x[690], x[646], x[645], x[644]}), .y(y[203]));
  R1ind204 R1ind204_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[792], x[791], x[790], x[819], x[696], x[695], x[694], x[661], x[660], x[659]}), .y(y[204]));
  R1ind205 R1ind205_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[796], x[795], x[794], x[820], x[700], x[699], x[698], x[655], x[654], x[653]}), .y(y[205]));
  R1ind206 R1ind206_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[800], x[799], x[798], x[821], x[704], x[703], x[702], x[640], x[639], x[638]}), .y(y[206]));
  R1ind207 R1ind207_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[804], x[803], x[802], x[822], x[708], x[707], x[706], x[649], x[648], x[647]}), .y(y[207]));
  R1ind208 R1ind208_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[808], x[807], x[806], x[823], x[712], x[711], x[710], x[643], x[642], x[641]}), .y(y[208]));
  R1ind209 R1ind209_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[812], x[811], x[810], x[824], x[716], x[715], x[714], x[652], x[651], x[650]}), .y(y[209]));
  R1ind210 R1ind210_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[816], x[815], x[814], x[825], x[720], x[719], x[718], x[658], x[657], x[656]}), .y(y[210]));
  R1ind211 R1ind211_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[646], x[645], x[644], x[829], x[724], x[723], x[722], x[828], x[827], x[826]}), .y(y[211]));
  R1ind212 R1ind212_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[661], x[660], x[659], x[833], x[728], x[727], x[726], x[832], x[831], x[830]}), .y(y[212]));
  R1ind213 R1ind213_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[655], x[654], x[653], x[837], x[732], x[731], x[730], x[836], x[835], x[834]}), .y(y[213]));
  R1ind214 R1ind214_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[640], x[639], x[638], x[841], x[736], x[735], x[734], x[840], x[839], x[838]}), .y(y[214]));
  R1ind215 R1ind215_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[649], x[648], x[647], x[845], x[740], x[739], x[738], x[844], x[843], x[842]}), .y(y[215]));
  R1ind216 R1ind216_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[643], x[642], x[641], x[849], x[744], x[743], x[742], x[848], x[847], x[846]}), .y(y[216]));
  R1ind217 R1ind217_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[652], x[651], x[650], x[853], x[748], x[747], x[746], x[852], x[851], x[850]}), .y(y[217]));
  R1ind218 R1ind218_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[658], x[657], x[656], x[857], x[752], x[751], x[750], x[856], x[855], x[854]}), .y(y[218]));
  R1ind219 R1ind219_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[828], x[827], x[826], x[861], x[756], x[755], x[754], x[860], x[859], x[858]}), .y(y[219]));
  R1ind220 R1ind220_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[832], x[831], x[830], x[865], x[760], x[759], x[758], x[864], x[863], x[862]}), .y(y[220]));
  R1ind221 R1ind221_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[836], x[835], x[834], x[869], x[764], x[763], x[762], x[868], x[867], x[866]}), .y(y[221]));
  R1ind222 R1ind222_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[840], x[839], x[838], x[873], x[768], x[767], x[766], x[872], x[871], x[870]}), .y(y[222]));
  R1ind223 R1ind223_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[844], x[843], x[842], x[877], x[772], x[771], x[770], x[876], x[875], x[874]}), .y(y[223]));
  R1ind224 R1ind224_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[848], x[847], x[846], x[881], x[776], x[775], x[774], x[880], x[879], x[878]}), .y(y[224]));
  R1ind225 R1ind225_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[852], x[851], x[850], x[885], x[780], x[779], x[778], x[884], x[883], x[882]}), .y(y[225]));
  R1ind226 R1ind226_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[856], x[855], x[854], x[889], x[784], x[783], x[782], x[888], x[887], x[886]}), .y(y[226]));
  R1ind227 R1ind227_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[860], x[859], x[858], x[893], x[788], x[787], x[786], x[892], x[891], x[890]}), .y(y[227]));
  R1ind228 R1ind228_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[864], x[863], x[862], x[897], x[792], x[791], x[790], x[896], x[895], x[894]}), .y(y[228]));
  R1ind229 R1ind229_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[868], x[867], x[866], x[901], x[796], x[795], x[794], x[900], x[899], x[898]}), .y(y[229]));
  R1ind230 R1ind230_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[872], x[871], x[870], x[905], x[800], x[799], x[798], x[904], x[903], x[902]}), .y(y[230]));
  R1ind231 R1ind231_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[876], x[875], x[874], x[909], x[804], x[803], x[802], x[908], x[907], x[906]}), .y(y[231]));
  R1ind232 R1ind232_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[880], x[879], x[878], x[913], x[808], x[807], x[806], x[912], x[911], x[910]}), .y(y[232]));
  R1ind233 R1ind233_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[884], x[883], x[882], x[917], x[812], x[811], x[810], x[916], x[915], x[914]}), .y(y[233]));
  R1ind234 R1ind234_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[888], x[887], x[886], x[921], x[816], x[815], x[814], x[920], x[919], x[918]}), .y(y[234]));
  R1ind235 R1ind235_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[892], x[891], x[890], x[922], x[646], x[645], x[644], x[441], x[440], x[439]}), .y(y[235]));
  R1ind236 R1ind236_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[896], x[895], x[894], x[923], x[661], x[660], x[659], x[454], x[453], x[452]}), .y(y[236]));
  R1ind237 R1ind237_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[900], x[899], x[898], x[924], x[655], x[654], x[653], x[464], x[463], x[462]}), .y(y[237]));
  R1ind238 R1ind238_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[904], x[903], x[902], x[925], x[640], x[639], x[638], x[474], x[473], x[472]}), .y(y[238]));
  R1ind239 R1ind239_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[908], x[907], x[906], x[926], x[649], x[648], x[647], x[484], x[483], x[482]}), .y(y[239]));
  R1ind240 R1ind240_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[912], x[911], x[910], x[927], x[643], x[642], x[641], x[494], x[493], x[492]}), .y(y[240]));
  R1ind241 R1ind241_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[916], x[915], x[914], x[928], x[652], x[651], x[650], x[504], x[503], x[502]}), .y(y[241]));
  R1ind242 R1ind242_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[920], x[919], x[918], x[929], x[658], x[657], x[656], x[514], x[513], x[512]}), .y(y[242]));
  R1ind243 R1ind243_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[441], x[440], x[439], x[930], x[828], x[827], x[826], x[524], x[523], x[522]}), .y(y[243]));
  R1ind244 R1ind244_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[454], x[453], x[452], x[931], x[832], x[831], x[830], x[531], x[530], x[529]}), .y(y[244]));
  R1ind245 R1ind245_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[464], x[463], x[462], x[932], x[836], x[835], x[834], x[538], x[537], x[536]}), .y(y[245]));
  R1ind246 R1ind246_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[474], x[473], x[472], x[933], x[840], x[839], x[838], x[545], x[544], x[543]}), .y(y[246]));
  R1ind247 R1ind247_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[484], x[483], x[482], x[934], x[844], x[843], x[842], x[552], x[551], x[550]}), .y(y[247]));
  R1ind248 R1ind248_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[494], x[493], x[492], x[935], x[848], x[847], x[846], x[559], x[558], x[557]}), .y(y[248]));
  R1ind249 R1ind249_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[504], x[503], x[502], x[936], x[852], x[851], x[850], x[566], x[565], x[564]}), .y(y[249]));
  R1ind250 R1ind250_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[514], x[513], x[512], x[937], x[856], x[855], x[854], x[573], x[572], x[571]}), .y(y[250]));
  R1ind251 R1ind251_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[524], x[523], x[522], x[938], x[860], x[859], x[858], x[580], x[579], x[578]}), .y(y[251]));
  R1ind252 R1ind252_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[531], x[530], x[529], x[939], x[864], x[863], x[862], x[587], x[586], x[585]}), .y(y[252]));
  R1ind253 R1ind253_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[538], x[537], x[536], x[940], x[868], x[867], x[866], x[594], x[593], x[592]}), .y(y[253]));
  R1ind254 R1ind254_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[545], x[544], x[543], x[941], x[872], x[871], x[870], x[601], x[600], x[599]}), .y(y[254]));
  R1ind255 R1ind255_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[552], x[551], x[550], x[942], x[876], x[875], x[874], x[608], x[607], x[606]}), .y(y[255]));
  R1ind256 R1ind256_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[559], x[558], x[557], x[943], x[880], x[879], x[878], x[615], x[614], x[613]}), .y(y[256]));
  R1ind257 R1ind257_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[566], x[565], x[564], x[944], x[884], x[883], x[882], x[622], x[621], x[620]}), .y(y[257]));
  R1ind258 R1ind258_inst(.x({x[410], x[409], x[408], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[573], x[572], x[571], x[945], x[888], x[887], x[886], x[629], x[628], x[627]}), .y(y[258]));
  R1ind259 R1ind259_inst(.x({x[432], x[431], x[430], x[435], x[434], x[433], x[426], x[425], x[424], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[429], x[428], x[427], x[401], x[400], x[399], x[392], x[391], x[390], x[404], x[403], x[402], x[410], x[409], x[408], x[395], x[394], x[393], x[398], x[397], x[396], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[580], x[579], x[578], x[946], x[892], x[891], x[890], x[445], x[444], x[443]}), .y(y[259]));
  R1ind260 R1ind260_inst(.x({x[432], x[431], x[430], x[435], x[434], x[433], x[426], x[425], x[424], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[429], x[428], x[427], x[401], x[400], x[399], x[392], x[391], x[390], x[404], x[403], x[402], x[410], x[409], x[408], x[395], x[394], x[393], x[398], x[397], x[396], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[587], x[586], x[585], x[947], x[896], x[895], x[894], x[458], x[457], x[456]}), .y(y[260]));
  R1ind261 R1ind261_inst(.x({x[432], x[431], x[430], x[435], x[434], x[433], x[426], x[425], x[424], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[429], x[428], x[427], x[401], x[400], x[399], x[392], x[391], x[390], x[404], x[403], x[402], x[410], x[409], x[408], x[395], x[394], x[393], x[398], x[397], x[396], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[594], x[593], x[592], x[948], x[900], x[899], x[898], x[468], x[467], x[466]}), .y(y[261]));
  R1ind262 R1ind262_inst(.x({x[432], x[431], x[430], x[435], x[434], x[433], x[426], x[425], x[424], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[429], x[428], x[427], x[401], x[400], x[399], x[392], x[391], x[390], x[404], x[403], x[402], x[410], x[409], x[408], x[395], x[394], x[393], x[398], x[397], x[396], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[601], x[600], x[599], x[949], x[904], x[903], x[902], x[478], x[477], x[476]}), .y(y[262]));
  R1ind263 R1ind263_inst(.x({x[432], x[431], x[430], x[435], x[434], x[433], x[426], x[425], x[424], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[429], x[428], x[427], x[401], x[400], x[399], x[392], x[391], x[390], x[404], x[403], x[402], x[410], x[409], x[408], x[395], x[394], x[393], x[398], x[397], x[396], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[608], x[607], x[606], x[950], x[908], x[907], x[906], x[488], x[487], x[486]}), .y(y[263]));
  R1ind264 R1ind264_inst(.x({x[432], x[431], x[430], x[435], x[434], x[433], x[426], x[425], x[424], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[429], x[428], x[427], x[401], x[400], x[399], x[392], x[391], x[390], x[404], x[403], x[402], x[410], x[409], x[408], x[395], x[394], x[393], x[398], x[397], x[396], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[615], x[614], x[613], x[951], x[912], x[911], x[910], x[498], x[497], x[496]}), .y(y[264]));
  R1ind265 R1ind265_inst(.x({x[432], x[431], x[430], x[435], x[434], x[433], x[426], x[425], x[424], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[429], x[428], x[427], x[401], x[400], x[399], x[392], x[391], x[390], x[404], x[403], x[402], x[410], x[409], x[408], x[395], x[394], x[393], x[398], x[397], x[396], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[622], x[621], x[620], x[952], x[916], x[915], x[914], x[508], x[507], x[506]}), .y(y[265]));
  R1ind266 R1ind266_inst(.x({x[432], x[431], x[430], x[435], x[434], x[433], x[426], x[425], x[424], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[429], x[428], x[427], x[401], x[400], x[399], x[392], x[391], x[390], x[404], x[403], x[402], x[410], x[409], x[408], x[395], x[394], x[393], x[398], x[397], x[396], x[407], x[406], x[405], x[448], x[447], x[446], x[389], x[388], x[387], x[629], x[628], x[627], x[953], x[920], x[919], x[918], x[518], x[517], x[516]}), .y(y[266]));
  R1ind267 R1ind267_inst(.x({x[458], x[457], x[456], x[518], x[517], x[516], x[5], x[4], x[3], x[468], x[467], x[466], x[20], x[19], x[18], x[508], x[507], x[506], x[8], x[7], x[6], x[488], x[487], x[486], x[14], x[13], x[12], x[661], x[660], x[659], x[658], x[657], x[656], x[655], x[654], x[653], x[652], x[651], x[650], x[649], x[648], x[647], x[646], x[645], x[644], x[498], x[497], x[496], x[11], x[10], x[9], x[478], x[477], x[476], x[17], x[16], x[15], x[643], x[642], x[641], x[640], x[639], x[638], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[23], x[22], x[21], x[448], x[447], x[446], x[404], x[403], x[402], x[218], x[217], x[216], x[122], x[121], x[120], x[311], x[310], x[309], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[445], x[444], x[443], x[26], x[25], x[24], x[314], x[313], x[312], x[389], x[388], x[387], x[954], x[362], x[361], x[360], x[386], x[385], x[384]}), .y(y[267]));
  R1ind268 R1ind268_inst(.x({x[488], x[487], x[486], x[14], x[13], x[12], x[518], x[517], x[516], x[5], x[4], x[3], x[508], x[507], x[506], x[8], x[7], x[6], x[468], x[467], x[466], x[649], x[648], x[647], x[478], x[477], x[476], x[17], x[16], x[15], x[658], x[657], x[656], x[652], x[651], x[650], x[655], x[654], x[653], x[661], x[660], x[659], x[498], x[497], x[496], x[11], x[10], x[9], x[445], x[444], x[443], x[26], x[25], x[24], x[640], x[639], x[638], x[643], x[642], x[641], x[646], x[645], x[644], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[20], x[19], x[18], x[448], x[447], x[446], x[404], x[403], x[402], x[215], x[214], x[213], x[119], x[118], x[117], x[308], x[307], x[306], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[458], x[457], x[456], x[23], x[22], x[21], x[311], x[310], x[309], x[389], x[388], x[387], x[955], x[359], x[358], x[357], x[383], x[382], x[381]}), .y(y[268]));
  R1ind269 R1ind269_inst(.x({x[488], x[487], x[486], x[14], x[13], x[12], x[458], x[457], x[456], x[23], x[22], x[21], x[478], x[477], x[476], x[649], x[648], x[647], x[518], x[517], x[516], x[5], x[4], x[3], x[508], x[507], x[506], x[8], x[7], x[6], x[655], x[654], x[653], x[661], x[660], x[659], x[640], x[639], x[638], x[658], x[657], x[656], x[652], x[651], x[650], x[498], x[497], x[496], x[11], x[10], x[9], x[445], x[444], x[443], x[26], x[25], x[24], x[643], x[642], x[641], x[646], x[645], x[644], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[17], x[16], x[15], x[448], x[447], x[446], x[404], x[403], x[402], x[212], x[211], x[210], x[116], x[115], x[114], x[305], x[304], x[303], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[468], x[467], x[466], x[20], x[19], x[18], x[308], x[307], x[306], x[389], x[388], x[387], x[956], x[356], x[355], x[354], x[380], x[379], x[378]}), .y(y[269]));
  R1ind270 R1ind270_inst(.x({x[458], x[457], x[456], x[23], x[22], x[21], x[468], x[467], x[466], x[20], x[19], x[18], x[508], x[507], x[506], x[8], x[7], x[6], x[488], x[487], x[486], x[661], x[660], x[659], x[518], x[517], x[516], x[5], x[4], x[3], x[445], x[444], x[443], x[655], x[654], x[653], x[652], x[651], x[650], x[649], x[648], x[647], x[658], x[657], x[656], x[646], x[645], x[644], x[498], x[497], x[496], x[11], x[10], x[9], x[643], x[642], x[641], x[640], x[639], x[638], x[14], x[13], x[12], x[26], x[25], x[24], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[302], x[301], x[300], x[314], x[313], x[312], x[448], x[447], x[446], x[404], x[403], x[402], x[209], x[208], x[207], x[113], x[112], x[111], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[478], x[477], x[476], x[17], x[16], x[15], x[305], x[304], x[303], x[389], x[388], x[387], x[957], x[353], x[352], x[351], x[377], x[376], x[375]}), .y(y[270]));
  R1ind271 R1ind271_inst(.x({x[508], x[507], x[506], x[8], x[7], x[6], x[649], x[648], x[647], x[468], x[467], x[466], x[20], x[19], x[18], x[458], x[457], x[456], x[23], x[22], x[21], x[652], x[651], x[650], x[655], x[654], x[653], x[661], x[660], x[659], x[498], x[497], x[496], x[478], x[477], x[476], x[17], x[16], x[15], x[445], x[444], x[443], x[518], x[517], x[516], x[5], x[4], x[3], x[643], x[642], x[641], x[640], x[639], x[638], x[646], x[645], x[644], x[658], x[657], x[656], x[11], x[10], x[9], x[26], x[25], x[24], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[299], x[298], x[297], x[314], x[313], x[312], x[448], x[447], x[446], x[404], x[403], x[402], x[206], x[205], x[204], x[110], x[109], x[108], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[488], x[487], x[486], x[14], x[13], x[12], x[302], x[301], x[300], x[389], x[388], x[387], x[958], x[350], x[349], x[348], x[374], x[373], x[372]}), .y(y[271]));
  R1ind272 R1ind272_inst(.x({x[488], x[487], x[486], x[14], x[13], x[12], x[458], x[457], x[456], x[23], x[22], x[21], x[508], x[507], x[506], x[468], x[467], x[466], x[20], x[19], x[18], x[445], x[444], x[443], x[26], x[25], x[24], x[649], x[648], x[647], x[661], x[660], x[659], x[518], x[517], x[516], x[5], x[4], x[3], x[652], x[651], x[650], x[655], x[654], x[653], x[646], x[645], x[644], x[478], x[477], x[476], x[17], x[16], x[15], x[658], x[657], x[656], x[643], x[642], x[641], x[640], x[639], x[638], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[8], x[7], x[6], x[448], x[447], x[446], x[404], x[403], x[402], x[203], x[202], x[201], x[107], x[106], x[105], x[296], x[295], x[294], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[498], x[497], x[496], x[11], x[10], x[9], x[299], x[298], x[297], x[389], x[388], x[387], x[959], x[347], x[346], x[345], x[371], x[370], x[369]}), .y(y[272]));
  R1ind273 R1ind273_inst(.x({x[488], x[487], x[486], x[14], x[13], x[12], x[649], x[648], x[647], x[652], x[651], x[650], x[498], x[497], x[496], x[11], x[10], x[9], x[478], x[477], x[476], x[17], x[16], x[15], x[445], x[444], x[443], x[468], x[467], x[466], x[20], x[19], x[18], x[458], x[457], x[456], x[23], x[22], x[21], x[643], x[642], x[641], x[640], x[639], x[638], x[646], x[645], x[644], x[655], x[654], x[653], x[661], x[660], x[659], x[518], x[517], x[516], x[658], x[657], x[656], x[5], x[4], x[3], x[26], x[25], x[24], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[293], x[292], x[291], x[314], x[313], x[312], x[448], x[447], x[446], x[404], x[403], x[402], x[104], x[103], x[102], x[200], x[199], x[198], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[508], x[507], x[506], x[8], x[7], x[6], x[296], x[295], x[294], x[389], x[388], x[387], x[960], x[344], x[343], x[342], x[368], x[367], x[366]}), .y(y[273]));
  R1ind274 R1ind274_inst(.x({x[458], x[457], x[456], x[23], x[22], x[21], x[661], x[660], x[659], x[468], x[467], x[466], x[20], x[19], x[18], x[488], x[487], x[486], x[14], x[13], x[12], x[508], x[507], x[506], x[8], x[7], x[6], x[445], x[444], x[443], x[655], x[654], x[653], x[649], x[648], x[647], x[652], x[651], x[650], x[646], x[645], x[644], x[498], x[497], x[496], x[11], x[10], x[9], x[478], x[477], x[476], x[17], x[16], x[15], x[658], x[657], x[656], x[643], x[642], x[641], x[640], x[639], x[638], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[26], x[25], x[24], x[448], x[447], x[446], x[404], x[403], x[402], x[101], x[100], x[99], x[197], x[196], x[195], x[314], x[313], x[312], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[518], x[517], x[516], x[5], x[4], x[3], x[293], x[292], x[291], x[389], x[388], x[387], x[961], x[341], x[340], x[339], x[365], x[364], x[363]}), .y(y[274]));
  R1ind275 R1ind275_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[386], x[385], x[384], x[962], x[338], x[337], x[336], x[362], x[361], x[360]}), .y(y[275]));
  R1ind276 R1ind276_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[383], x[382], x[381], x[963], x[335], x[334], x[333], x[359], x[358], x[357]}), .y(y[276]));
  R1ind277 R1ind277_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[380], x[379], x[378], x[964], x[332], x[331], x[330], x[356], x[355], x[354]}), .y(y[277]));
  R1ind278 R1ind278_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[377], x[376], x[375], x[965], x[329], x[328], x[327], x[353], x[352], x[351]}), .y(y[278]));
  R1ind279 R1ind279_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[374], x[373], x[372], x[966], x[326], x[325], x[324], x[350], x[349], x[348]}), .y(y[279]));
  R1ind280 R1ind280_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[371], x[370], x[369], x[967], x[323], x[322], x[321], x[347], x[346], x[345]}), .y(y[280]));
  R1ind281 R1ind281_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[368], x[367], x[366], x[968], x[320], x[319], x[318], x[344], x[343], x[342]}), .y(y[281]));
  R1ind282 R1ind282_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[365], x[364], x[363], x[969], x[317], x[316], x[315], x[341], x[340], x[339]}), .y(y[282]));
  R1ind283 R1ind283_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[362], x[361], x[360], x[970], x[314], x[313], x[312], x[338], x[337], x[336]}), .y(y[283]));
  R1ind284 R1ind284_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[359], x[358], x[357], x[971], x[311], x[310], x[309], x[335], x[334], x[333]}), .y(y[284]));
  R1ind285 R1ind285_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[356], x[355], x[354], x[972], x[308], x[307], x[306], x[332], x[331], x[330]}), .y(y[285]));
  R1ind286 R1ind286_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[353], x[352], x[351], x[973], x[305], x[304], x[303], x[329], x[328], x[327]}), .y(y[286]));
  R1ind287 R1ind287_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[350], x[349], x[348], x[974], x[302], x[301], x[300], x[326], x[325], x[324]}), .y(y[287]));
  R1ind288 R1ind288_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[347], x[346], x[345], x[975], x[299], x[298], x[297], x[323], x[322], x[321]}), .y(y[288]));
  R1ind289 R1ind289_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[344], x[343], x[342], x[976], x[296], x[295], x[294], x[320], x[319], x[318]}), .y(y[289]));
  R1ind290 R1ind290_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[341], x[340], x[339], x[977], x[293], x[292], x[291], x[317], x[316], x[315]}), .y(y[290]));
  R1ind291 R1ind291_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[338], x[337], x[336], x[978], x[386], x[385], x[384], x[314], x[313], x[312]}), .y(y[291]));
  R1ind292 R1ind292_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[335], x[334], x[333], x[979], x[383], x[382], x[381], x[311], x[310], x[309]}), .y(y[292]));
  R1ind293 R1ind293_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[332], x[331], x[330], x[980], x[380], x[379], x[378], x[308], x[307], x[306]}), .y(y[293]));
  R1ind294 R1ind294_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[329], x[328], x[327], x[981], x[377], x[376], x[375], x[305], x[304], x[303]}), .y(y[294]));
  R1ind295 R1ind295_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[326], x[325], x[324], x[982], x[374], x[373], x[372], x[302], x[301], x[300]}), .y(y[295]));
  R1ind296 R1ind296_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[323], x[322], x[321], x[983], x[371], x[370], x[369], x[299], x[298], x[297]}), .y(y[296]));
  R1ind297 R1ind297_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[320], x[319], x[318], x[984], x[368], x[367], x[366], x[296], x[295], x[294]}), .y(y[297]));
  R1ind298 R1ind298_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[317], x[316], x[315], x[985], x[365], x[364], x[363], x[293], x[292], x[291]}), .y(y[298]));
  R1ind299 R1ind299_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[311], x[310], x[309], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[122], x[121], x[120], x[26], x[25], x[24], x[215], x[214], x[213], x[407], x[406], x[405], x[218], x[217], x[216], x[389], x[388], x[387], x[314], x[313], x[312], x[986], x[242], x[241], x[240], x[290], x[289], x[288]}), .y(y[299]));
  R1ind300 R1ind300_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[308], x[307], x[306], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[119], x[118], x[117], x[23], x[22], x[21], x[212], x[211], x[210], x[407], x[406], x[405], x[215], x[214], x[213], x[389], x[388], x[387], x[311], x[310], x[309], x[987], x[239], x[238], x[237], x[287], x[286], x[285]}), .y(y[300]));
  R1ind301 R1ind301_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[305], x[304], x[303], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[116], x[115], x[114], x[20], x[19], x[18], x[209], x[208], x[207], x[407], x[406], x[405], x[212], x[211], x[210], x[389], x[388], x[387], x[308], x[307], x[306], x[988], x[236], x[235], x[234], x[284], x[283], x[282]}), .y(y[301]));
  R1ind302 R1ind302_inst(.x({x[302], x[301], x[300], x[314], x[313], x[312], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[206], x[205], x[204], x[218], x[217], x[216], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[113], x[112], x[111], x[17], x[16], x[15], x[407], x[406], x[405], x[209], x[208], x[207], x[389], x[388], x[387], x[305], x[304], x[303], x[989], x[233], x[232], x[231], x[281], x[280], x[279]}), .y(y[302]));
  R1ind303 R1ind303_inst(.x({x[299], x[298], x[297], x[314], x[313], x[312], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[203], x[202], x[201], x[218], x[217], x[216], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[110], x[109], x[108], x[14], x[13], x[12], x[407], x[406], x[405], x[206], x[205], x[204], x[389], x[388], x[387], x[302], x[301], x[300], x[990], x[230], x[229], x[228], x[278], x[277], x[276]}), .y(y[303]));
  R1ind304 R1ind304_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[296], x[295], x[294], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[107], x[106], x[105], x[11], x[10], x[9], x[200], x[199], x[198], x[407], x[406], x[405], x[203], x[202], x[201], x[389], x[388], x[387], x[299], x[298], x[297], x[991], x[227], x[226], x[225], x[275], x[274], x[273]}), .y(y[304]));
  R1ind305 R1ind305_inst(.x({x[293], x[292], x[291], x[314], x[313], x[312], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[197], x[196], x[195], x[218], x[217], x[216], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[8], x[7], x[6], x[104], x[103], x[102], x[407], x[406], x[405], x[200], x[199], x[198], x[389], x[388], x[387], x[296], x[295], x[294], x[992], x[224], x[223], x[222], x[272], x[271], x[270]}), .y(y[305]));
  R1ind306 R1ind306_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[314], x[313], x[312], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[5], x[4], x[3], x[101], x[100], x[99], x[218], x[217], x[216], x[407], x[406], x[405], x[197], x[196], x[195], x[389], x[388], x[387], x[293], x[292], x[291], x[993], x[221], x[220], x[219], x[269], x[268], x[267]}), .y(y[306]));
  R1ind307 R1ind307_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[290], x[289], x[288], x[994], x[218], x[217], x[216], x[266], x[265], x[264]}), .y(y[307]));
  R1ind308 R1ind308_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[287], x[286], x[285], x[995], x[215], x[214], x[213], x[263], x[262], x[261]}), .y(y[308]));
  R1ind309 R1ind309_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[284], x[283], x[282], x[996], x[212], x[211], x[210], x[260], x[259], x[258]}), .y(y[309]));
  R1ind310 R1ind310_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[281], x[280], x[279], x[997], x[209], x[208], x[207], x[257], x[256], x[255]}), .y(y[310]));
  R1ind311 R1ind311_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[278], x[277], x[276], x[998], x[206], x[205], x[204], x[254], x[253], x[252]}), .y(y[311]));
  R1ind312 R1ind312_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[275], x[274], x[273], x[999], x[203], x[202], x[201], x[251], x[250], x[249]}), .y(y[312]));
  R1ind313 R1ind313_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[272], x[271], x[270], x[1000], x[200], x[199], x[198], x[248], x[247], x[246]}), .y(y[313]));
  R1ind314 R1ind314_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[269], x[268], x[267], x[1001], x[197], x[196], x[195], x[245], x[244], x[243]}), .y(y[314]));
  R1ind315 R1ind315_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[266], x[265], x[264], x[1002], x[290], x[289], x[288], x[242], x[241], x[240]}), .y(y[315]));
  R1ind316 R1ind316_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[263], x[262], x[261], x[1003], x[287], x[286], x[285], x[239], x[238], x[237]}), .y(y[316]));
  R1ind317 R1ind317_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[260], x[259], x[258], x[1004], x[284], x[283], x[282], x[236], x[235], x[234]}), .y(y[317]));
  R1ind318 R1ind318_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[257], x[256], x[255], x[1005], x[281], x[280], x[279], x[233], x[232], x[231]}), .y(y[318]));
  R1ind319 R1ind319_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[254], x[253], x[252], x[1006], x[278], x[277], x[276], x[230], x[229], x[228]}), .y(y[319]));
  R1ind320 R1ind320_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[251], x[250], x[249], x[1007], x[275], x[274], x[273], x[227], x[226], x[225]}), .y(y[320]));
  R1ind321 R1ind321_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[248], x[247], x[246], x[1008], x[272], x[271], x[270], x[224], x[223], x[222]}), .y(y[321]));
  R1ind322 R1ind322_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[245], x[244], x[243], x[1009], x[269], x[268], x[267], x[221], x[220], x[219]}), .y(y[322]));
  R1ind323 R1ind323_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[242], x[241], x[240], x[1010], x[266], x[265], x[264], x[218], x[217], x[216]}), .y(y[323]));
  R1ind324 R1ind324_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[239], x[238], x[237], x[1011], x[263], x[262], x[261], x[215], x[214], x[213]}), .y(y[324]));
  R1ind325 R1ind325_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[236], x[235], x[234], x[1012], x[260], x[259], x[258], x[212], x[211], x[210]}), .y(y[325]));
  R1ind326 R1ind326_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[233], x[232], x[231], x[1013], x[257], x[256], x[255], x[209], x[208], x[207]}), .y(y[326]));
  R1ind327 R1ind327_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[230], x[229], x[228], x[1014], x[254], x[253], x[252], x[206], x[205], x[204]}), .y(y[327]));
  R1ind328 R1ind328_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[227], x[226], x[225], x[1015], x[251], x[250], x[249], x[203], x[202], x[201]}), .y(y[328]));
  R1ind329 R1ind329_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[224], x[223], x[222], x[1016], x[248], x[247], x[246], x[200], x[199], x[198]}), .y(y[329]));
  R1ind330 R1ind330_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[221], x[220], x[219], x[1017], x[245], x[244], x[243], x[197], x[196], x[195]}), .y(y[330]));
  R1ind331 R1ind331_inst(.x({x[410], x[409], x[408], x[215], x[214], x[213], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[26], x[25], x[24], x[314], x[313], x[312], x[119], x[118], x[117], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[218], x[217], x[216], x[389], x[388], x[387], x[1018], x[122], x[121], x[120], x[194], x[193], x[192]}), .y(y[331]));
  R1ind332 R1ind332_inst(.x({x[410], x[409], x[408], x[212], x[211], x[210], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[23], x[22], x[21], x[311], x[310], x[309], x[116], x[115], x[114], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[215], x[214], x[213], x[389], x[388], x[387], x[1019], x[119], x[118], x[117], x[191], x[190], x[189]}), .y(y[332]));
  R1ind333 R1ind333_inst(.x({x[410], x[409], x[408], x[209], x[208], x[207], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[20], x[19], x[18], x[308], x[307], x[306], x[113], x[112], x[111], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[212], x[211], x[210], x[389], x[388], x[387], x[1020], x[116], x[115], x[114], x[188], x[187], x[186]}), .y(y[333]));
  R1ind334 R1ind334_inst(.x({x[206], x[205], x[204], x[218], x[217], x[216], x[410], x[409], x[408], x[110], x[109], x[108], x[122], x[121], x[120], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[17], x[16], x[15], x[305], x[304], x[303], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[209], x[208], x[207], x[389], x[388], x[387], x[1021], x[113], x[112], x[111], x[185], x[184], x[183]}), .y(y[334]));
  R1ind335 R1ind335_inst(.x({x[203], x[202], x[201], x[218], x[217], x[216], x[410], x[409], x[408], x[107], x[106], x[105], x[122], x[121], x[120], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[14], x[13], x[12], x[302], x[301], x[300], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[206], x[205], x[204], x[389], x[388], x[387], x[1022], x[110], x[109], x[108], x[182], x[181], x[180]}), .y(y[335]));
  R1ind336 R1ind336_inst(.x({x[410], x[409], x[408], x[200], x[199], x[198], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[11], x[10], x[9], x[299], x[298], x[297], x[104], x[103], x[102], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[203], x[202], x[201], x[389], x[388], x[387], x[1023], x[107], x[106], x[105], x[179], x[178], x[177]}), .y(y[336]));
  R1ind337 R1ind337_inst(.x({x[197], x[196], x[195], x[218], x[217], x[216], x[410], x[409], x[408], x[101], x[100], x[99], x[122], x[121], x[120], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[296], x[295], x[294], x[8], x[7], x[6], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[200], x[199], x[198], x[389], x[388], x[387], x[1024], x[104], x[103], x[102], x[176], x[175], x[174]}), .y(y[337]));
  R1ind338 R1ind338_inst(.x({x[410], x[409], x[408], x[218], x[217], x[216], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[293], x[292], x[291], x[5], x[4], x[3], x[122], x[121], x[120], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[197], x[196], x[195], x[389], x[388], x[387], x[1025], x[101], x[100], x[99], x[173], x[172], x[171]}), .y(y[338]));
  R1ind339 R1ind339_inst(.x({x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387], x[1026], x[194], x[193], x[192], x[170], x[169], x[168]}), .y(y[339]));
  R1ind340 R1ind340_inst(.x({x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387], x[1027], x[191], x[190], x[189], x[167], x[166], x[165]}), .y(y[340]));
  R1ind341 R1ind341_inst(.x({x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387], x[1028], x[188], x[187], x[186], x[164], x[163], x[162]}), .y(y[341]));
  R1ind342 R1ind342_inst(.x({x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387], x[1029], x[185], x[184], x[183], x[161], x[160], x[159]}), .y(y[342]));
  R1ind343 R1ind343_inst(.x({x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387], x[1030], x[182], x[181], x[180], x[158], x[157], x[156]}), .y(y[343]));
  R1ind344 R1ind344_inst(.x({x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387], x[1031], x[179], x[178], x[177], x[155], x[154], x[153]}), .y(y[344]));
  R1ind345 R1ind345_inst(.x({x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387], x[1032], x[176], x[175], x[174], x[152], x[151], x[150]}), .y(y[345]));
  R1ind346 R1ind346_inst(.x({x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387], x[1033], x[173], x[172], x[171], x[149], x[148], x[147]}), .y(y[346]));
  R1ind347 R1ind347_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1034], x[170], x[169], x[168], x[146], x[145], x[144]}), .y(y[347]));
  R1ind348 R1ind348_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1035], x[167], x[166], x[165], x[143], x[142], x[141]}), .y(y[348]));
  R1ind349 R1ind349_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1036], x[164], x[163], x[162], x[140], x[139], x[138]}), .y(y[349]));
  R1ind350 R1ind350_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1037], x[161], x[160], x[159], x[137], x[136], x[135]}), .y(y[350]));
  R1ind351 R1ind351_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1038], x[158], x[157], x[156], x[134], x[133], x[132]}), .y(y[351]));
  R1ind352 R1ind352_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1039], x[155], x[154], x[153], x[131], x[130], x[129]}), .y(y[352]));
  R1ind353 R1ind353_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1040], x[152], x[151], x[150], x[128], x[127], x[126]}), .y(y[353]));
  R1ind354 R1ind354_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1041], x[149], x[148], x[147], x[125], x[124], x[123]}), .y(y[354]));
  R1ind355 R1ind355_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1042], x[146], x[145], x[144], x[122], x[121], x[120]}), .y(y[355]));
  R1ind356 R1ind356_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1043], x[143], x[142], x[141], x[119], x[118], x[117]}), .y(y[356]));
  R1ind357 R1ind357_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1044], x[140], x[139], x[138], x[116], x[115], x[114]}), .y(y[357]));
  R1ind358 R1ind358_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1045], x[137], x[136], x[135], x[113], x[112], x[111]}), .y(y[358]));
  R1ind359 R1ind359_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1046], x[134], x[133], x[132], x[110], x[109], x[108]}), .y(y[359]));
  R1ind360 R1ind360_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1047], x[131], x[130], x[129], x[107], x[106], x[105]}), .y(y[360]));
  R1ind361 R1ind361_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1048], x[128], x[127], x[126], x[104], x[103], x[102]}), .y(y[361]));
  R1ind362 R1ind362_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[1049], x[125], x[124], x[123], x[101], x[100], x[99]}), .y(y[362]));
  R1ind363 R1ind363_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[119], x[118], x[117], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[314], x[313], x[312], x[218], x[217], x[216], x[23], x[22], x[21], x[407], x[406], x[405], x[26], x[25], x[24], x[389], x[388], x[387], x[122], x[121], x[120], x[1050], x[98], x[97], x[96]}), .y(y[363]));
  R1ind364 R1ind364_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[116], x[115], x[114], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[311], x[310], x[309], x[215], x[214], x[213], x[20], x[19], x[18], x[407], x[406], x[405], x[23], x[22], x[21], x[389], x[388], x[387], x[119], x[118], x[117], x[1051], x[95], x[94], x[93]}), .y(y[364]));
  R1ind365 R1ind365_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[113], x[112], x[111], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[308], x[307], x[306], x[212], x[211], x[210], x[17], x[16], x[15], x[407], x[406], x[405], x[20], x[19], x[18], x[389], x[388], x[387], x[116], x[115], x[114], x[1052], x[92], x[91], x[90]}), .y(y[365]));
  R1ind366 R1ind366_inst(.x({x[110], x[109], x[108], x[122], x[121], x[120], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[14], x[13], x[12], x[26], x[25], x[24], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[305], x[304], x[303], x[209], x[208], x[207], x[407], x[406], x[405], x[17], x[16], x[15], x[389], x[388], x[387], x[113], x[112], x[111], x[1053], x[89], x[88], x[87]}), .y(y[366]));
  R1ind367 R1ind367_inst(.x({x[107], x[106], x[105], x[122], x[121], x[120], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[11], x[10], x[9], x[26], x[25], x[24], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[302], x[301], x[300], x[206], x[205], x[204], x[407], x[406], x[405], x[14], x[13], x[12], x[389], x[388], x[387], x[110], x[109], x[108], x[1054], x[86], x[85], x[84]}), .y(y[367]));
  R1ind368 R1ind368_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[104], x[103], x[102], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[299], x[298], x[297], x[203], x[202], x[201], x[8], x[7], x[6], x[407], x[406], x[405], x[11], x[10], x[9], x[389], x[388], x[387], x[107], x[106], x[105], x[1055], x[83], x[82], x[81]}), .y(y[368]));
  R1ind369 R1ind369_inst(.x({x[101], x[100], x[99], x[122], x[121], x[120], x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[5], x[4], x[3], x[26], x[25], x[24], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[200], x[199], x[198], x[296], x[295], x[294], x[407], x[406], x[405], x[8], x[7], x[6], x[389], x[388], x[387], x[104], x[103], x[102], x[1056], x[80], x[79], x[78]}), .y(y[369]));
  R1ind370 R1ind370_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[122], x[121], x[120], x[448], x[447], x[446], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[197], x[196], x[195], x[293], x[292], x[291], x[26], x[25], x[24], x[407], x[406], x[405], x[5], x[4], x[3], x[389], x[388], x[387], x[101], x[100], x[99], x[1057], x[77], x[76], x[75]}), .y(y[370]));
  R1ind371 R1ind371_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[98], x[97], x[96], x[1058], x[74], x[73], x[72]}), .y(y[371]));
  R1ind372 R1ind372_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[95], x[94], x[93], x[1059], x[71], x[70], x[69]}), .y(y[372]));
  R1ind373 R1ind373_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[92], x[91], x[90], x[1060], x[68], x[67], x[66]}), .y(y[373]));
  R1ind374 R1ind374_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[89], x[88], x[87], x[1061], x[65], x[64], x[63]}), .y(y[374]));
  R1ind375 R1ind375_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[86], x[85], x[84], x[1062], x[62], x[61], x[60]}), .y(y[375]));
  R1ind376 R1ind376_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[83], x[82], x[81], x[1063], x[59], x[58], x[57]}), .y(y[376]));
  R1ind377 R1ind377_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[80], x[79], x[78], x[1064], x[56], x[55], x[54]}), .y(y[377]));
  R1ind378 R1ind378_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[77], x[76], x[75], x[1065], x[53], x[52], x[51]}), .y(y[378]));
  R1ind379 R1ind379_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[74], x[73], x[72], x[1066], x[50], x[49], x[48]}), .y(y[379]));
  R1ind380 R1ind380_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[71], x[70], x[69], x[1067], x[47], x[46], x[45]}), .y(y[380]));
  R1ind381 R1ind381_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[68], x[67], x[66], x[1068], x[44], x[43], x[42]}), .y(y[381]));
  R1ind382 R1ind382_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[65], x[64], x[63], x[1069], x[41], x[40], x[39]}), .y(y[382]));
  R1ind383 R1ind383_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[62], x[61], x[60], x[1070], x[38], x[37], x[36]}), .y(y[383]));
  R1ind384 R1ind384_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[59], x[58], x[57], x[1071], x[35], x[34], x[33]}), .y(y[384]));
  R1ind385 R1ind385_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[56], x[55], x[54], x[1072], x[32], x[31], x[30]}), .y(y[385]));
  R1ind386 R1ind386_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[53], x[52], x[51], x[1073], x[29], x[28], x[27]}), .y(y[386]));
  R1ind387 R1ind387_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[50], x[49], x[48], x[1074], x[26], x[25], x[24]}), .y(y[387]));
  R1ind388 R1ind388_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[47], x[46], x[45], x[1075], x[23], x[22], x[21]}), .y(y[388]));
  R1ind389 R1ind389_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[44], x[43], x[42], x[1076], x[20], x[19], x[18]}), .y(y[389]));
  R1ind390 R1ind390_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[41], x[40], x[39], x[1077], x[17], x[16], x[15]}), .y(y[390]));
  R1ind391 R1ind391_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[38], x[37], x[36], x[1078], x[14], x[13], x[12]}), .y(y[391]));
  R1ind392 R1ind392_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[35], x[34], x[33], x[1079], x[11], x[10], x[9]}), .y(y[392]));
  R1ind393 R1ind393_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[32], x[31], x[30], x[1080], x[8], x[7], x[6]}), .y(y[393]));
  R1ind394 R1ind394_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[29], x[28], x[27], x[1081], x[5], x[4], x[3]}), .y(y[394]));
  R1ind395 R1ind395_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[407], x[406], x[405], x[389], x[388], x[387]}), .y(y[395]));
  R1ind396 R1ind396_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[404], x[403], x[402], x[410], x[409], x[408], x[407], x[406], x[405], x[389], x[388], x[387], x[448], x[447], x[446]}), .y(y[396]));
  R1ind397 R1ind397_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[404], x[403], x[402], x[410], x[409], x[408]}), .y(y[397]));
  R1ind398 R1ind398_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[413], x[412], x[411], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[410], x[409], x[408], x[389], x[388], x[387], x[404], x[403], x[402]}), .y(y[398]));
  R1ind399 R1ind399_inst(.x({x[419], x[418], x[417], x[413], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[416], x[415], x[414], x[389], x[388], x[387], x[422], x[421], x[420]}), .y(y[399]));
  R1ind400 R1ind400_inst(.x({x[422], x[421], x[420], x[413], x[412], x[411], x[410], x[409], x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[419], x[418], x[417], x[389], x[388], x[387], x[416], x[415], x[414]}), .y(y[400]));
  R1ind401 R1ind401_inst(.x({x[422], x[421], x[420], x[416], x[415], x[414], x[413], x[412], x[411], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[407], x[406], x[405], x[389], x[388], x[387], x[419], x[418], x[417]}), .y(y[401]));
  R1ind402 R1ind402_inst(.x({x[422], x[421], x[420], x[419], x[418], x[417], x[416], x[415], x[414], x[410], x[409], x[408], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[413], x[412], x[411], x[389], x[388], x[387], x[407], x[406], x[405]}), .y(y[402]));
  R1ind403 R1ind403_inst(.x({x[419], x[418], x[417], x[416], x[415], x[414], x[410], x[409], x[408], x[407], x[406], x[405], x[404], x[403], x[402], x[401], x[400], x[399], x[398], x[397], x[396], x[395], x[394], x[393], x[392], x[391], x[390], x[422], x[421], x[420], x[389], x[388], x[387], x[413], x[412], x[411]}), .y(y[403]));
endmodule

module R2ind0(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (t[2] & ~t[3]);
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[1];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [35:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[13] & t[1];
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[21] | t[22]);
  assign t[12] = ~(t[23] | t[24]);
  assign t[13] = (t[25]);
  assign t[14] = (t[26]);
  assign t[15] = (t[27]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = t[2] & t[3];
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = t[37] ^ x[2];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[8];
  assign t[28] = t[40] ^ x[11];
  assign t[29] = t[41] ^ x[14];
  assign t[2] = ~(t[4] | t[5]);
  assign t[30] = t[42] ^ x[17];
  assign t[31] = t[43] ^ x[20];
  assign t[32] = t[44] ^ x[23];
  assign t[33] = t[45] ^ x[26];
  assign t[34] = t[46] ^ x[29];
  assign t[35] = t[47] ^ x[32];
  assign t[36] = t[48] ^ x[35];
  assign t[37] = (t[49] & ~t[50]);
  assign t[38] = (t[51] & ~t[52]);
  assign t[39] = (t[53] & ~t[54]);
  assign t[3] = ~(t[6] | t[7]);
  assign t[40] = (t[55] & ~t[56]);
  assign t[41] = (t[57] & ~t[58]);
  assign t[42] = (t[59] & ~t[60]);
  assign t[43] = (t[61] & ~t[62]);
  assign t[44] = (t[63] & ~t[64]);
  assign t[45] = (t[65] & ~t[66]);
  assign t[46] = (t[67] & ~t[68]);
  assign t[47] = (t[69] & ~t[70]);
  assign t[48] = (t[71] & ~t[72]);
  assign t[49] = t[73] ^ x[2];
  assign t[4] = ~(t[14] & t[15]);
  assign t[50] = t[74] ^ x[1];
  assign t[51] = t[75] ^ x[5];
  assign t[52] = t[76] ^ x[4];
  assign t[53] = t[77] ^ x[8];
  assign t[54] = t[78] ^ x[7];
  assign t[55] = t[79] ^ x[11];
  assign t[56] = t[80] ^ x[10];
  assign t[57] = t[81] ^ x[14];
  assign t[58] = t[82] ^ x[13];
  assign t[59] = t[83] ^ x[17];
  assign t[5] = ~(t[16] & t[17]);
  assign t[60] = t[84] ^ x[16];
  assign t[61] = t[85] ^ x[20];
  assign t[62] = t[86] ^ x[19];
  assign t[63] = t[87] ^ x[23];
  assign t[64] = t[88] ^ x[22];
  assign t[65] = t[89] ^ x[26];
  assign t[66] = t[90] ^ x[25];
  assign t[67] = t[91] ^ x[29];
  assign t[68] = t[92] ^ x[28];
  assign t[69] = t[93] ^ x[32];
  assign t[6] = ~(t[8]);
  assign t[70] = t[94] ^ x[31];
  assign t[71] = t[95] ^ x[35];
  assign t[72] = t[96] ^ x[34];
  assign t[73] = (x[0]);
  assign t[74] = (x[0]);
  assign t[75] = (x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[6]);
  assign t[78] = (x[6]);
  assign t[79] = (x[9]);
  assign t[7] = ~(t[18] & t[9]);
  assign t[80] = (x[9]);
  assign t[81] = (x[12]);
  assign t[82] = (x[12]);
  assign t[83] = (x[15]);
  assign t[84] = (x[15]);
  assign t[85] = (x[18]);
  assign t[86] = (x[18]);
  assign t[87] = (x[21]);
  assign t[88] = (x[21]);
  assign t[89] = (x[24]);
  assign t[8] = ~(t[19] | t[10]);
  assign t[90] = (x[24]);
  assign t[91] = (x[27]);
  assign t[92] = (x[27]);
  assign t[93] = (x[30]);
  assign t[94] = (x[30]);
  assign t[95] = (x[33]);
  assign t[96] = (x[33]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind3(x, y);
 input [35:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[13] & t[1];
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[21] | t[22]);
  assign t[12] = ~(t[23] | t[24]);
  assign t[13] = (t[25]);
  assign t[14] = (t[26]);
  assign t[15] = (t[27]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = t[2] & t[3];
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = t[37] ^ x[2];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[8];
  assign t[28] = t[40] ^ x[11];
  assign t[29] = t[41] ^ x[14];
  assign t[2] = ~(t[4] | t[5]);
  assign t[30] = t[42] ^ x[17];
  assign t[31] = t[43] ^ x[20];
  assign t[32] = t[44] ^ x[23];
  assign t[33] = t[45] ^ x[26];
  assign t[34] = t[46] ^ x[29];
  assign t[35] = t[47] ^ x[32];
  assign t[36] = t[48] ^ x[35];
  assign t[37] = (t[49] & ~t[50]);
  assign t[38] = (t[51] & ~t[52]);
  assign t[39] = (t[53] & ~t[54]);
  assign t[3] = ~(t[6] | t[7]);
  assign t[40] = (t[55] & ~t[56]);
  assign t[41] = (t[57] & ~t[58]);
  assign t[42] = (t[59] & ~t[60]);
  assign t[43] = (t[61] & ~t[62]);
  assign t[44] = (t[63] & ~t[64]);
  assign t[45] = (t[65] & ~t[66]);
  assign t[46] = (t[67] & ~t[68]);
  assign t[47] = (t[69] & ~t[70]);
  assign t[48] = (t[71] & ~t[72]);
  assign t[49] = t[73] ^ x[2];
  assign t[4] = ~(t[14] & t[15]);
  assign t[50] = t[74] ^ x[1];
  assign t[51] = t[75] ^ x[5];
  assign t[52] = t[76] ^ x[4];
  assign t[53] = t[77] ^ x[8];
  assign t[54] = t[78] ^ x[7];
  assign t[55] = t[79] ^ x[11];
  assign t[56] = t[80] ^ x[10];
  assign t[57] = t[81] ^ x[14];
  assign t[58] = t[82] ^ x[13];
  assign t[59] = t[83] ^ x[17];
  assign t[5] = ~(t[16] & t[17]);
  assign t[60] = t[84] ^ x[16];
  assign t[61] = t[85] ^ x[20];
  assign t[62] = t[86] ^ x[19];
  assign t[63] = t[87] ^ x[23];
  assign t[64] = t[88] ^ x[22];
  assign t[65] = t[89] ^ x[26];
  assign t[66] = t[90] ^ x[25];
  assign t[67] = t[91] ^ x[29];
  assign t[68] = t[92] ^ x[28];
  assign t[69] = t[93] ^ x[32];
  assign t[6] = ~(t[8]);
  assign t[70] = t[94] ^ x[31];
  assign t[71] = t[95] ^ x[35];
  assign t[72] = t[96] ^ x[34];
  assign t[73] = (x[0]);
  assign t[74] = (x[0]);
  assign t[75] = (x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[6]);
  assign t[78] = (x[6]);
  assign t[79] = (x[9]);
  assign t[7] = ~(t[18] & t[9]);
  assign t[80] = (x[9]);
  assign t[81] = (x[12]);
  assign t[82] = (x[12]);
  assign t[83] = (x[15]);
  assign t[84] = (x[15]);
  assign t[85] = (x[18]);
  assign t[86] = (x[18]);
  assign t[87] = (x[21]);
  assign t[88] = (x[21]);
  assign t[89] = (x[24]);
  assign t[8] = ~(t[19] | t[10]);
  assign t[90] = (x[24]);
  assign t[91] = (x[27]);
  assign t[92] = (x[27]);
  assign t[93] = (x[30]);
  assign t[94] = (x[30]);
  assign t[95] = (x[33]);
  assign t[96] = (x[33]);
  assign t[9] = ~(t[20]);
  assign y = (t[0]);
endmodule

module R2ind4(x, y);
 input x;
 output y;

 wire t;
  assign t = ~(x);
  assign y = (t);
endmodule

module R2ind5(x, y);
 input x;
 output y;

 wire t;
  assign t = ~(x);
  assign y = (t);
endmodule

module R2ind6(x, y);
 input [17:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[2];
  assign t[13] = t[19] ^ x[5];
  assign t[14] = t[20] ^ x[8];
  assign t[15] = t[21] ^ x[11];
  assign t[16] = t[22] ^ x[14];
  assign t[17] = t[23] ^ x[17];
  assign t[18] = (t[24] & ~t[25]);
  assign t[19] = (t[26] & ~t[27]);
  assign t[1] = ~(t[6] & t[2]);
  assign t[20] = (t[28] & ~t[29]);
  assign t[21] = (t[30] & ~t[31]);
  assign t[22] = (t[32] & ~t[33]);
  assign t[23] = (t[34] & ~t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[1];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[4];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[7];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[10];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[13];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[16];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[46] = (x[15]);
  assign t[47] = (x[15]);
  assign t[4] = ~(t[8] | t[9]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind7(x, y);
 input [17:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = t[18] ^ x[2];
  assign t[13] = t[19] ^ x[5];
  assign t[14] = t[20] ^ x[8];
  assign t[15] = t[21] ^ x[11];
  assign t[16] = t[22] ^ x[14];
  assign t[17] = t[23] ^ x[17];
  assign t[18] = (t[24] & ~t[25]);
  assign t[19] = (t[26] & ~t[27]);
  assign t[1] = ~(t[6] & t[2]);
  assign t[20] = (t[28] & ~t[29]);
  assign t[21] = (t[30] & ~t[31]);
  assign t[22] = (t[32] & ~t[33]);
  assign t[23] = (t[34] & ~t[35]);
  assign t[24] = t[36] ^ x[2];
  assign t[25] = t[37] ^ x[1];
  assign t[26] = t[38] ^ x[5];
  assign t[27] = t[39] ^ x[4];
  assign t[28] = t[40] ^ x[8];
  assign t[29] = t[41] ^ x[7];
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = t[42] ^ x[11];
  assign t[31] = t[43] ^ x[10];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[13];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[16];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[46] = (x[15]);
  assign t[47] = (x[15]);
  assign t[4] = ~(t[8] | t[9]);
  assign t[5] = ~(t[10] | t[11]);
  assign t[6] = (t[12]);
  assign t[7] = (t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind8(x, y);
 input [26:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = t[28] ^ x[2];
  assign t[1] = ~(t[3] & t[10]);
  assign t[20] = t[29] ^ x[5];
  assign t[21] = t[30] ^ x[8];
  assign t[22] = t[31] ^ x[11];
  assign t[23] = t[32] ^ x[14];
  assign t[24] = t[33] ^ x[17];
  assign t[25] = t[34] ^ x[20];
  assign t[26] = t[35] ^ x[23];
  assign t[27] = t[36] ^ x[26];
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = (t[39] & ~t[40]);
  assign t[2] = ~(t[11] & t[4]);
  assign t[30] = (t[41] & ~t[42]);
  assign t[31] = (t[43] & ~t[44]);
  assign t[32] = (t[45] & ~t[46]);
  assign t[33] = (t[47] & ~t[48]);
  assign t[34] = (t[49] & ~t[50]);
  assign t[35] = (t[51] & ~t[52]);
  assign t[36] = (t[53] & ~t[54]);
  assign t[37] = t[55] ^ x[2];
  assign t[38] = t[56] ^ x[1];
  assign t[39] = t[57] ^ x[5];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[58] ^ x[4];
  assign t[41] = t[59] ^ x[8];
  assign t[42] = t[60] ^ x[7];
  assign t[43] = t[61] ^ x[11];
  assign t[44] = t[62] ^ x[10];
  assign t[45] = t[63] ^ x[14];
  assign t[46] = t[64] ^ x[13];
  assign t[47] = t[65] ^ x[17];
  assign t[48] = t[66] ^ x[16];
  assign t[49] = t[67] ^ x[20];
  assign t[4] = ~(t[12] | t[7]);
  assign t[50] = t[68] ^ x[19];
  assign t[51] = t[69] ^ x[23];
  assign t[52] = t[70] ^ x[22];
  assign t[53] = t[71] ^ x[26];
  assign t[54] = t[72] ^ x[25];
  assign t[55] = (x[0]);
  assign t[56] = (x[0]);
  assign t[57] = (x[3]);
  assign t[58] = (x[3]);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[6]);
  assign t[61] = (x[9]);
  assign t[62] = (x[9]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[15]);
  assign t[66] = (x[15]);
  assign t[67] = (x[18]);
  assign t[68] = (x[18]);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[13] | t[14]);
  assign t[70] = (x[21]);
  assign t[71] = (x[24]);
  assign t[72] = (x[24]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[15] | t[16]);
  assign t[9] = ~(t[17] | t[18]);
  assign y = (t[0]);
endmodule

module R2ind9(x, y);
 input [26:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = t[28] ^ x[2];
  assign t[1] = ~(t[3] & t[10]);
  assign t[20] = t[29] ^ x[5];
  assign t[21] = t[30] ^ x[8];
  assign t[22] = t[31] ^ x[11];
  assign t[23] = t[32] ^ x[14];
  assign t[24] = t[33] ^ x[17];
  assign t[25] = t[34] ^ x[20];
  assign t[26] = t[35] ^ x[23];
  assign t[27] = t[36] ^ x[26];
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = (t[39] & ~t[40]);
  assign t[2] = ~(t[11] & t[4]);
  assign t[30] = (t[41] & ~t[42]);
  assign t[31] = (t[43] & ~t[44]);
  assign t[32] = (t[45] & ~t[46]);
  assign t[33] = (t[47] & ~t[48]);
  assign t[34] = (t[49] & ~t[50]);
  assign t[35] = (t[51] & ~t[52]);
  assign t[36] = (t[53] & ~t[54]);
  assign t[37] = t[55] ^ x[2];
  assign t[38] = t[56] ^ x[1];
  assign t[39] = t[57] ^ x[5];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[58] ^ x[4];
  assign t[41] = t[59] ^ x[8];
  assign t[42] = t[60] ^ x[7];
  assign t[43] = t[61] ^ x[11];
  assign t[44] = t[62] ^ x[10];
  assign t[45] = t[63] ^ x[14];
  assign t[46] = t[64] ^ x[13];
  assign t[47] = t[65] ^ x[17];
  assign t[48] = t[66] ^ x[16];
  assign t[49] = t[67] ^ x[20];
  assign t[4] = ~(t[12] | t[7]);
  assign t[50] = t[68] ^ x[19];
  assign t[51] = t[69] ^ x[23];
  assign t[52] = t[70] ^ x[22];
  assign t[53] = t[71] ^ x[26];
  assign t[54] = t[72] ^ x[25];
  assign t[55] = (x[0]);
  assign t[56] = (x[0]);
  assign t[57] = (x[3]);
  assign t[58] = (x[3]);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[6]);
  assign t[61] = (x[9]);
  assign t[62] = (x[9]);
  assign t[63] = (x[12]);
  assign t[64] = (x[12]);
  assign t[65] = (x[15]);
  assign t[66] = (x[15]);
  assign t[67] = (x[18]);
  assign t[68] = (x[18]);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[13] | t[14]);
  assign t[70] = (x[21]);
  assign t[71] = (x[24]);
  assign t[72] = (x[24]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[15] | t[16]);
  assign t[9] = ~(t[17] | t[18]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [41:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[22] & t[1]);
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[15]);
  assign t[103] = (x[15]);
  assign t[104] = (x[18]);
  assign t[105] = (x[18]);
  assign t[106] = (x[21]);
  assign t[107] = (x[21]);
  assign t[108] = (x[24]);
  assign t[109] = (x[24]);
  assign t[10] = t[12] & t[13];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[30]);
  assign t[113] = (x[30]);
  assign t[114] = (x[33]);
  assign t[115] = (x[33]);
  assign t[116] = (x[36]);
  assign t[117] = (x[36]);
  assign t[118] = (x[39]);
  assign t[119] = (x[39]);
  assign t[11] = ~(t[25] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[11]);
  assign t[18] = ~(t[30] & t[21]);
  assign t[19] = ~(t[31] | t[32]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[20] = ~(t[33] | t[34]);
  assign t[21] = ~(t[35]);
  assign t[22] = (t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = t[50] ^ x[2];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[11];
  assign t[3] = ~(t[23]);
  assign t[40] = t[54] ^ x[14];
  assign t[41] = t[55] ^ x[17];
  assign t[42] = t[56] ^ x[20];
  assign t[43] = t[57] ^ x[23];
  assign t[44] = t[58] ^ x[26];
  assign t[45] = t[59] ^ x[29];
  assign t[46] = t[60] ^ x[32];
  assign t[47] = t[61] ^ x[35];
  assign t[48] = t[62] ^ x[38];
  assign t[49] = t[63] ^ x[41];
  assign t[4] = ~(t[24]);
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = (t[76] & ~t[77]);
  assign t[57] = (t[78] & ~t[79]);
  assign t[58] = (t[80] & ~t[81]);
  assign t[59] = (t[82] & ~t[83]);
  assign t[5] = t[6] & t[7];
  assign t[60] = (t[84] & ~t[85]);
  assign t[61] = (t[86] & ~t[87]);
  assign t[62] = (t[88] & ~t[89]);
  assign t[63] = (t[90] & ~t[91]);
  assign t[64] = t[92] ^ x[2];
  assign t[65] = t[93] ^ x[1];
  assign t[66] = t[94] ^ x[5];
  assign t[67] = t[95] ^ x[4];
  assign t[68] = t[96] ^ x[8];
  assign t[69] = t[97] ^ x[7];
  assign t[6] = ~(t[8]);
  assign t[70] = t[98] ^ x[11];
  assign t[71] = t[99] ^ x[10];
  assign t[72] = t[100] ^ x[14];
  assign t[73] = t[101] ^ x[13];
  assign t[74] = t[102] ^ x[17];
  assign t[75] = t[103] ^ x[16];
  assign t[76] = t[104] ^ x[20];
  assign t[77] = t[105] ^ x[19];
  assign t[78] = t[106] ^ x[23];
  assign t[79] = t[107] ^ x[22];
  assign t[7] = ~(t[9]);
  assign t[80] = t[108] ^ x[26];
  assign t[81] = t[109] ^ x[25];
  assign t[82] = t[110] ^ x[29];
  assign t[83] = t[111] ^ x[28];
  assign t[84] = t[112] ^ x[32];
  assign t[85] = t[113] ^ x[31];
  assign t[86] = t[114] ^ x[35];
  assign t[87] = t[115] ^ x[34];
  assign t[88] = t[116] ^ x[38];
  assign t[89] = t[117] ^ x[37];
  assign t[8] = t[22] & t[10];
  assign t[90] = t[118] ^ x[41];
  assign t[91] = t[119] ^ x[40];
  assign t[92] = (x[0]);
  assign t[93] = (x[0]);
  assign t[94] = (x[3]);
  assign t[95] = (x[3]);
  assign t[96] = (x[6]);
  assign t[97] = (x[6]);
  assign t[98] = (x[9]);
  assign t[99] = (x[9]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind11(x, y);
 input [41:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[22] & t[1]);
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[15]);
  assign t[103] = (x[15]);
  assign t[104] = (x[18]);
  assign t[105] = (x[18]);
  assign t[106] = (x[21]);
  assign t[107] = (x[21]);
  assign t[108] = (x[24]);
  assign t[109] = (x[24]);
  assign t[10] = t[12] & t[13];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[30]);
  assign t[113] = (x[30]);
  assign t[114] = (x[33]);
  assign t[115] = (x[33]);
  assign t[116] = (x[36]);
  assign t[117] = (x[36]);
  assign t[118] = (x[39]);
  assign t[119] = (x[39]);
  assign t[11] = ~(t[25] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[11]);
  assign t[18] = ~(t[30] & t[21]);
  assign t[19] = ~(t[31] | t[32]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[20] = ~(t[33] | t[34]);
  assign t[21] = ~(t[35]);
  assign t[22] = (t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = t[50] ^ x[2];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[11];
  assign t[3] = ~(t[23]);
  assign t[40] = t[54] ^ x[14];
  assign t[41] = t[55] ^ x[17];
  assign t[42] = t[56] ^ x[20];
  assign t[43] = t[57] ^ x[23];
  assign t[44] = t[58] ^ x[26];
  assign t[45] = t[59] ^ x[29];
  assign t[46] = t[60] ^ x[32];
  assign t[47] = t[61] ^ x[35];
  assign t[48] = t[62] ^ x[38];
  assign t[49] = t[63] ^ x[41];
  assign t[4] = ~(t[24]);
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = (t[76] & ~t[77]);
  assign t[57] = (t[78] & ~t[79]);
  assign t[58] = (t[80] & ~t[81]);
  assign t[59] = (t[82] & ~t[83]);
  assign t[5] = t[6] & t[7];
  assign t[60] = (t[84] & ~t[85]);
  assign t[61] = (t[86] & ~t[87]);
  assign t[62] = (t[88] & ~t[89]);
  assign t[63] = (t[90] & ~t[91]);
  assign t[64] = t[92] ^ x[2];
  assign t[65] = t[93] ^ x[1];
  assign t[66] = t[94] ^ x[5];
  assign t[67] = t[95] ^ x[4];
  assign t[68] = t[96] ^ x[8];
  assign t[69] = t[97] ^ x[7];
  assign t[6] = ~(t[8]);
  assign t[70] = t[98] ^ x[11];
  assign t[71] = t[99] ^ x[10];
  assign t[72] = t[100] ^ x[14];
  assign t[73] = t[101] ^ x[13];
  assign t[74] = t[102] ^ x[17];
  assign t[75] = t[103] ^ x[16];
  assign t[76] = t[104] ^ x[20];
  assign t[77] = t[105] ^ x[19];
  assign t[78] = t[106] ^ x[23];
  assign t[79] = t[107] ^ x[22];
  assign t[7] = ~(t[9]);
  assign t[80] = t[108] ^ x[26];
  assign t[81] = t[109] ^ x[25];
  assign t[82] = t[110] ^ x[29];
  assign t[83] = t[111] ^ x[28];
  assign t[84] = t[112] ^ x[32];
  assign t[85] = t[113] ^ x[31];
  assign t[86] = t[114] ^ x[35];
  assign t[87] = t[115] ^ x[34];
  assign t[88] = t[116] ^ x[38];
  assign t[89] = t[117] ^ x[37];
  assign t[8] = t[22] & t[10];
  assign t[90] = t[118] ^ x[41];
  assign t[91] = t[119] ^ x[40];
  assign t[92] = (x[0]);
  assign t[93] = (x[0]);
  assign t[94] = (x[3]);
  assign t[95] = (x[3]);
  assign t[96] = (x[6]);
  assign t[97] = (x[6]);
  assign t[98] = (x[9]);
  assign t[99] = (x[9]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind12(x, y);
 input [38:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18]);
  assign t[102] = (x[18]);
  assign t[103] = (x[21]);
  assign t[104] = (x[21]);
  assign t[105] = (x[24]);
  assign t[106] = (x[24]);
  assign t[107] = (x[27]);
  assign t[108] = (x[27]);
  assign t[109] = (x[30]);
  assign t[10] = t[26] & t[12];
  assign t[110] = (x[30]);
  assign t[111] = (x[33]);
  assign t[112] = (x[33]);
  assign t[113] = (x[36]);
  assign t[114] = (x[36]);
  assign t[11] = ~(t[26] & t[13]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] | t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[28] & t[25]);
  assign t[18] = ~(t[29] & t[30]);
  assign t[19] = ~(t[13]);
  assign t[1] = ~(t[24] & t[3]);
  assign t[20] = ~(t[31] & t[23]);
  assign t[21] = ~(t[32] | t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36]);
  assign t[24] = (t[37]);
  assign t[25] = (t[38]);
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[25] & t[4]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = t[50] ^ x[2];
  assign t[38] = t[51] ^ x[5];
  assign t[39] = t[52] ^ x[8];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[53] ^ x[11];
  assign t[41] = t[54] ^ x[14];
  assign t[42] = t[55] ^ x[17];
  assign t[43] = t[56] ^ x[20];
  assign t[44] = t[57] ^ x[23];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[29];
  assign t[47] = t[60] ^ x[32];
  assign t[48] = t[61] ^ x[35];
  assign t[49] = t[62] ^ x[38];
  assign t[4] = ~(t[7] | t[6]);
  assign t[50] = (t[63] & ~t[64]);
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = t[89] ^ x[2];
  assign t[64] = t[90] ^ x[1];
  assign t[65] = t[91] ^ x[5];
  assign t[66] = t[92] ^ x[4];
  assign t[67] = t[93] ^ x[8];
  assign t[68] = t[94] ^ x[7];
  assign t[69] = t[95] ^ x[11];
  assign t[6] = ~(t[26]);
  assign t[70] = t[96] ^ x[10];
  assign t[71] = t[97] ^ x[14];
  assign t[72] = t[98] ^ x[13];
  assign t[73] = t[99] ^ x[17];
  assign t[74] = t[100] ^ x[16];
  assign t[75] = t[101] ^ x[20];
  assign t[76] = t[102] ^ x[19];
  assign t[77] = t[103] ^ x[23];
  assign t[78] = t[104] ^ x[22];
  assign t[79] = t[105] ^ x[26];
  assign t[7] = ~(t[5]);
  assign t[80] = t[106] ^ x[25];
  assign t[81] = t[107] ^ x[29];
  assign t[82] = t[108] ^ x[28];
  assign t[83] = t[109] ^ x[32];
  assign t[84] = t[110] ^ x[31];
  assign t[85] = t[111] ^ x[35];
  assign t[86] = t[112] ^ x[34];
  assign t[87] = t[113] ^ x[38];
  assign t[88] = t[114] ^ x[37];
  assign t[89] = (x[0]);
  assign t[8] = ~(t[10]);
  assign t[90] = (x[0]);
  assign t[91] = (x[3]);
  assign t[92] = (x[3]);
  assign t[93] = (x[6]);
  assign t[94] = (x[6]);
  assign t[95] = (x[9]);
  assign t[96] = (x[9]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[15]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind13(x, y);
 input [38:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[15]);
  assign t[101] = (x[18]);
  assign t[102] = (x[18]);
  assign t[103] = (x[21]);
  assign t[104] = (x[21]);
  assign t[105] = (x[24]);
  assign t[106] = (x[24]);
  assign t[107] = (x[27]);
  assign t[108] = (x[27]);
  assign t[109] = (x[30]);
  assign t[10] = t[26] & t[12];
  assign t[110] = (x[30]);
  assign t[111] = (x[33]);
  assign t[112] = (x[33]);
  assign t[113] = (x[36]);
  assign t[114] = (x[36]);
  assign t[11] = ~(t[26] & t[13]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] | t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[28] & t[25]);
  assign t[18] = ~(t[29] & t[30]);
  assign t[19] = ~(t[13]);
  assign t[1] = ~(t[24] & t[3]);
  assign t[20] = ~(t[31] & t[23]);
  assign t[21] = ~(t[32] | t[33]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36]);
  assign t[24] = (t[37]);
  assign t[25] = (t[38]);
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = ~(t[25] & t[4]);
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = (t[48]);
  assign t[36] = (t[49]);
  assign t[37] = t[50] ^ x[2];
  assign t[38] = t[51] ^ x[5];
  assign t[39] = t[52] ^ x[8];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[53] ^ x[11];
  assign t[41] = t[54] ^ x[14];
  assign t[42] = t[55] ^ x[17];
  assign t[43] = t[56] ^ x[20];
  assign t[44] = t[57] ^ x[23];
  assign t[45] = t[58] ^ x[26];
  assign t[46] = t[59] ^ x[29];
  assign t[47] = t[60] ^ x[32];
  assign t[48] = t[61] ^ x[35];
  assign t[49] = t[62] ^ x[38];
  assign t[4] = ~(t[7] | t[6]);
  assign t[50] = (t[63] & ~t[64]);
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] & t[9];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = t[89] ^ x[2];
  assign t[64] = t[90] ^ x[1];
  assign t[65] = t[91] ^ x[5];
  assign t[66] = t[92] ^ x[4];
  assign t[67] = t[93] ^ x[8];
  assign t[68] = t[94] ^ x[7];
  assign t[69] = t[95] ^ x[11];
  assign t[6] = ~(t[26]);
  assign t[70] = t[96] ^ x[10];
  assign t[71] = t[97] ^ x[14];
  assign t[72] = t[98] ^ x[13];
  assign t[73] = t[99] ^ x[17];
  assign t[74] = t[100] ^ x[16];
  assign t[75] = t[101] ^ x[20];
  assign t[76] = t[102] ^ x[19];
  assign t[77] = t[103] ^ x[23];
  assign t[78] = t[104] ^ x[22];
  assign t[79] = t[105] ^ x[26];
  assign t[7] = ~(t[5]);
  assign t[80] = t[106] ^ x[25];
  assign t[81] = t[107] ^ x[29];
  assign t[82] = t[108] ^ x[28];
  assign t[83] = t[109] ^ x[32];
  assign t[84] = t[110] ^ x[31];
  assign t[85] = t[111] ^ x[35];
  assign t[86] = t[112] ^ x[34];
  assign t[87] = t[113] ^ x[38];
  assign t[88] = t[114] ^ x[37];
  assign t[89] = (x[0]);
  assign t[8] = ~(t[10]);
  assign t[90] = (x[0]);
  assign t[91] = (x[3]);
  assign t[92] = (x[3]);
  assign t[93] = (x[6]);
  assign t[94] = (x[6]);
  assign t[95] = (x[9]);
  assign t[96] = (x[9]);
  assign t[97] = (x[12]);
  assign t[98] = (x[12]);
  assign t[99] = (x[15]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind14(x, y);
 input [35:0] x;
 output y;

 wire [107:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[24]);
  assign t[101] = (x[24]);
  assign t[102] = (x[27]);
  assign t[103] = (x[27]);
  assign t[104] = (x[30]);
  assign t[105] = (x[30]);
  assign t[106] = (x[33]);
  assign t[107] = (x[33]);
  assign t[10] = t[26] & t[12];
  assign t[11] = ~(t[26] & t[13]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] | t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[28] & t[24]);
  assign t[18] = ~(t[25] & t[29]);
  assign t[19] = ~(t[13]);
  assign t[1] = ~(t[24] & t[3]);
  assign t[20] = ~(t[30] & t[23]);
  assign t[21] = ~(t[31] | t[32]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[23] = ~(t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = (t[41]);
  assign t[2] = ~(t[25] & t[4]);
  assign t[30] = (t[42]);
  assign t[31] = (t[43]);
  assign t[32] = (t[44]);
  assign t[33] = (t[45]);
  assign t[34] = (t[46]);
  assign t[35] = (t[47]);
  assign t[36] = t[48] ^ x[2];
  assign t[37] = t[49] ^ x[5];
  assign t[38] = t[50] ^ x[8];
  assign t[39] = t[51] ^ x[11];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[52] ^ x[14];
  assign t[41] = t[53] ^ x[17];
  assign t[42] = t[54] ^ x[20];
  assign t[43] = t[55] ^ x[23];
  assign t[44] = t[56] ^ x[26];
  assign t[45] = t[57] ^ x[29];
  assign t[46] = t[58] ^ x[32];
  assign t[47] = t[59] ^ x[35];
  assign t[48] = (t[60] & ~t[61]);
  assign t[49] = (t[62] & ~t[63]);
  assign t[4] = ~(t[7] | t[6]);
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = (t[76] & ~t[77]);
  assign t[57] = (t[78] & ~t[79]);
  assign t[58] = (t[80] & ~t[81]);
  assign t[59] = (t[82] & ~t[83]);
  assign t[5] = t[8] & t[9];
  assign t[60] = t[84] ^ x[2];
  assign t[61] = t[85] ^ x[1];
  assign t[62] = t[86] ^ x[5];
  assign t[63] = t[87] ^ x[4];
  assign t[64] = t[88] ^ x[8];
  assign t[65] = t[89] ^ x[7];
  assign t[66] = t[90] ^ x[11];
  assign t[67] = t[91] ^ x[10];
  assign t[68] = t[92] ^ x[14];
  assign t[69] = t[93] ^ x[13];
  assign t[6] = ~(t[26]);
  assign t[70] = t[94] ^ x[17];
  assign t[71] = t[95] ^ x[16];
  assign t[72] = t[96] ^ x[20];
  assign t[73] = t[97] ^ x[19];
  assign t[74] = t[98] ^ x[23];
  assign t[75] = t[99] ^ x[22];
  assign t[76] = t[100] ^ x[26];
  assign t[77] = t[101] ^ x[25];
  assign t[78] = t[102] ^ x[29];
  assign t[79] = t[103] ^ x[28];
  assign t[7] = ~(t[5]);
  assign t[80] = t[104] ^ x[32];
  assign t[81] = t[105] ^ x[31];
  assign t[82] = t[106] ^ x[35];
  assign t[83] = t[107] ^ x[34];
  assign t[84] = (x[0]);
  assign t[85] = (x[0]);
  assign t[86] = (x[3]);
  assign t[87] = (x[3]);
  assign t[88] = (x[6]);
  assign t[89] = (x[6]);
  assign t[8] = ~(t[10]);
  assign t[90] = (x[9]);
  assign t[91] = (x[9]);
  assign t[92] = (x[12]);
  assign t[93] = (x[12]);
  assign t[94] = (x[15]);
  assign t[95] = (x[15]);
  assign t[96] = (x[18]);
  assign t[97] = (x[18]);
  assign t[98] = (x[21]);
  assign t[99] = (x[21]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [35:0] x;
 output y;

 wire [107:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[24]);
  assign t[101] = (x[24]);
  assign t[102] = (x[27]);
  assign t[103] = (x[27]);
  assign t[104] = (x[30]);
  assign t[105] = (x[30]);
  assign t[106] = (x[33]);
  assign t[107] = (x[33]);
  assign t[10] = t[26] & t[12];
  assign t[11] = ~(t[26] & t[13]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] | t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[21] & t[22]);
  assign t[17] = ~(t[28] & t[24]);
  assign t[18] = ~(t[25] & t[29]);
  assign t[19] = ~(t[13]);
  assign t[1] = ~(t[24] & t[3]);
  assign t[20] = ~(t[30] & t[23]);
  assign t[21] = ~(t[31] | t[32]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[23] = ~(t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = (t[41]);
  assign t[2] = ~(t[25] & t[4]);
  assign t[30] = (t[42]);
  assign t[31] = (t[43]);
  assign t[32] = (t[44]);
  assign t[33] = (t[45]);
  assign t[34] = (t[46]);
  assign t[35] = (t[47]);
  assign t[36] = t[48] ^ x[2];
  assign t[37] = t[49] ^ x[5];
  assign t[38] = t[50] ^ x[8];
  assign t[39] = t[51] ^ x[11];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[52] ^ x[14];
  assign t[41] = t[53] ^ x[17];
  assign t[42] = t[54] ^ x[20];
  assign t[43] = t[55] ^ x[23];
  assign t[44] = t[56] ^ x[26];
  assign t[45] = t[57] ^ x[29];
  assign t[46] = t[58] ^ x[32];
  assign t[47] = t[59] ^ x[35];
  assign t[48] = (t[60] & ~t[61]);
  assign t[49] = (t[62] & ~t[63]);
  assign t[4] = ~(t[7] | t[6]);
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = (t[76] & ~t[77]);
  assign t[57] = (t[78] & ~t[79]);
  assign t[58] = (t[80] & ~t[81]);
  assign t[59] = (t[82] & ~t[83]);
  assign t[5] = t[8] & t[9];
  assign t[60] = t[84] ^ x[2];
  assign t[61] = t[85] ^ x[1];
  assign t[62] = t[86] ^ x[5];
  assign t[63] = t[87] ^ x[4];
  assign t[64] = t[88] ^ x[8];
  assign t[65] = t[89] ^ x[7];
  assign t[66] = t[90] ^ x[11];
  assign t[67] = t[91] ^ x[10];
  assign t[68] = t[92] ^ x[14];
  assign t[69] = t[93] ^ x[13];
  assign t[6] = ~(t[26]);
  assign t[70] = t[94] ^ x[17];
  assign t[71] = t[95] ^ x[16];
  assign t[72] = t[96] ^ x[20];
  assign t[73] = t[97] ^ x[19];
  assign t[74] = t[98] ^ x[23];
  assign t[75] = t[99] ^ x[22];
  assign t[76] = t[100] ^ x[26];
  assign t[77] = t[101] ^ x[25];
  assign t[78] = t[102] ^ x[29];
  assign t[79] = t[103] ^ x[28];
  assign t[7] = ~(t[5]);
  assign t[80] = t[104] ^ x[32];
  assign t[81] = t[105] ^ x[31];
  assign t[82] = t[106] ^ x[35];
  assign t[83] = t[107] ^ x[34];
  assign t[84] = (x[0]);
  assign t[85] = (x[0]);
  assign t[86] = (x[3]);
  assign t[87] = (x[3]);
  assign t[88] = (x[6]);
  assign t[89] = (x[6]);
  assign t[8] = ~(t[10]);
  assign t[90] = (x[9]);
  assign t[91] = (x[9]);
  assign t[92] = (x[12]);
  assign t[93] = (x[12]);
  assign t[94] = (x[15]);
  assign t[95] = (x[15]);
  assign t[96] = (x[18]);
  assign t[97] = (x[18]);
  assign t[98] = (x[21]);
  assign t[99] = (x[21]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind16(x, y);
 input [41:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = t[11] & t[12];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[12] = ~(t[14]);
  assign t[13] = t[30] & t[15];
  assign t[14] = ~(t[30] & t[16]);
  assign t[15] = t[17] & t[18];
  assign t[16] = ~(t[31] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[32] & t[33]);
  assign t[21] = ~(t[27] & t[34]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[35] & t[26]);
  assign t[24] = ~(t[36] | t[37]);
  assign t[25] = ~(t[38] | t[39]);
  assign t[26] = ~(t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[27] & t[5]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = t[6] ^ t[7];
  assign t[40] = (t[54]);
  assign t[41] = t[55] ^ x[2];
  assign t[42] = t[56] ^ x[5];
  assign t[43] = t[57] ^ x[8];
  assign t[44] = t[58] ^ x[11];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[20];
  assign t[48] = t[62] ^ x[23];
  assign t[49] = t[63] ^ x[26];
  assign t[4] = ~(t[8] | t[9]);
  assign t[50] = t[64] ^ x[29];
  assign t[51] = t[65] ^ x[32];
  assign t[52] = t[66] ^ x[35];
  assign t[53] = t[67] ^ x[38];
  assign t[54] = t[68] ^ x[41];
  assign t[55] = (t[69] & ~t[70]);
  assign t[56] = (t[71] & ~t[72]);
  assign t[57] = (t[73] & ~t[74]);
  assign t[58] = (t[75] & ~t[76]);
  assign t[59] = (t[77] & ~t[78]);
  assign t[5] = ~(t[10] | t[9]);
  assign t[60] = (t[79] & ~t[80]);
  assign t[61] = (t[81] & ~t[82]);
  assign t[62] = (t[83] & ~t[84]);
  assign t[63] = (t[85] & ~t[86]);
  assign t[64] = (t[87] & ~t[88]);
  assign t[65] = (t[89] & ~t[90]);
  assign t[66] = (t[91] & ~t[92]);
  assign t[67] = (t[93] & ~t[94]);
  assign t[68] = (t[95] & ~t[96]);
  assign t[69] = t[97] ^ x[2];
  assign t[6] = ~(t[28]);
  assign t[70] = t[98] ^ x[1];
  assign t[71] = t[99] ^ x[5];
  assign t[72] = t[100] ^ x[4];
  assign t[73] = t[101] ^ x[8];
  assign t[74] = t[102] ^ x[7];
  assign t[75] = t[103] ^ x[11];
  assign t[76] = t[104] ^ x[10];
  assign t[77] = t[105] ^ x[14];
  assign t[78] = t[106] ^ x[13];
  assign t[79] = t[107] ^ x[17];
  assign t[7] = ~(t[29]);
  assign t[80] = t[108] ^ x[16];
  assign t[81] = t[109] ^ x[20];
  assign t[82] = t[110] ^ x[19];
  assign t[83] = t[111] ^ x[23];
  assign t[84] = t[112] ^ x[22];
  assign t[85] = t[113] ^ x[26];
  assign t[86] = t[114] ^ x[25];
  assign t[87] = t[115] ^ x[29];
  assign t[88] = t[116] ^ x[28];
  assign t[89] = t[117] ^ x[32];
  assign t[8] = ~(t[10]);
  assign t[90] = t[118] ^ x[31];
  assign t[91] = t[119] ^ x[35];
  assign t[92] = t[120] ^ x[34];
  assign t[93] = t[121] ^ x[38];
  assign t[94] = t[122] ^ x[37];
  assign t[95] = t[123] ^ x[41];
  assign t[96] = t[124] ^ x[40];
  assign t[97] = (x[0]);
  assign t[98] = (x[0]);
  assign t[99] = (x[3]);
  assign t[9] = ~(t[30]);
  assign y = (t[0]);
endmodule

module R2ind17(x, y);
 input [41:0] x;
 output y;

 wire [124:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[3]);
  assign t[101] = (x[6]);
  assign t[102] = (x[6]);
  assign t[103] = (x[9]);
  assign t[104] = (x[9]);
  assign t[105] = (x[12]);
  assign t[106] = (x[12]);
  assign t[107] = (x[15]);
  assign t[108] = (x[15]);
  assign t[109] = (x[18]);
  assign t[10] = t[11] & t[12];
  assign t[110] = (x[18]);
  assign t[111] = (x[21]);
  assign t[112] = (x[21]);
  assign t[113] = (x[24]);
  assign t[114] = (x[24]);
  assign t[115] = (x[27]);
  assign t[116] = (x[27]);
  assign t[117] = (x[30]);
  assign t[118] = (x[30]);
  assign t[119] = (x[33]);
  assign t[11] = ~(t[13]);
  assign t[120] = (x[33]);
  assign t[121] = (x[36]);
  assign t[122] = (x[36]);
  assign t[123] = (x[39]);
  assign t[124] = (x[39]);
  assign t[12] = ~(t[14]);
  assign t[13] = t[30] & t[15];
  assign t[14] = ~(t[30] & t[16]);
  assign t[15] = t[17] & t[18];
  assign t[16] = ~(t[31] | t[19]);
  assign t[17] = ~(t[20] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[32] & t[33]);
  assign t[21] = ~(t[27] & t[34]);
  assign t[22] = ~(t[16]);
  assign t[23] = ~(t[35] & t[26]);
  assign t[24] = ~(t[36] | t[37]);
  assign t[25] = ~(t[38] | t[39]);
  assign t[26] = ~(t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[27] & t[5]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = t[6] ^ t[7];
  assign t[40] = (t[54]);
  assign t[41] = t[55] ^ x[2];
  assign t[42] = t[56] ^ x[5];
  assign t[43] = t[57] ^ x[8];
  assign t[44] = t[58] ^ x[11];
  assign t[45] = t[59] ^ x[14];
  assign t[46] = t[60] ^ x[17];
  assign t[47] = t[61] ^ x[20];
  assign t[48] = t[62] ^ x[23];
  assign t[49] = t[63] ^ x[26];
  assign t[4] = ~(t[8] | t[9]);
  assign t[50] = t[64] ^ x[29];
  assign t[51] = t[65] ^ x[32];
  assign t[52] = t[66] ^ x[35];
  assign t[53] = t[67] ^ x[38];
  assign t[54] = t[68] ^ x[41];
  assign t[55] = (t[69] & ~t[70]);
  assign t[56] = (t[71] & ~t[72]);
  assign t[57] = (t[73] & ~t[74]);
  assign t[58] = (t[75] & ~t[76]);
  assign t[59] = (t[77] & ~t[78]);
  assign t[5] = ~(t[10] | t[9]);
  assign t[60] = (t[79] & ~t[80]);
  assign t[61] = (t[81] & ~t[82]);
  assign t[62] = (t[83] & ~t[84]);
  assign t[63] = (t[85] & ~t[86]);
  assign t[64] = (t[87] & ~t[88]);
  assign t[65] = (t[89] & ~t[90]);
  assign t[66] = (t[91] & ~t[92]);
  assign t[67] = (t[93] & ~t[94]);
  assign t[68] = (t[95] & ~t[96]);
  assign t[69] = t[97] ^ x[2];
  assign t[6] = ~(t[28]);
  assign t[70] = t[98] ^ x[1];
  assign t[71] = t[99] ^ x[5];
  assign t[72] = t[100] ^ x[4];
  assign t[73] = t[101] ^ x[8];
  assign t[74] = t[102] ^ x[7];
  assign t[75] = t[103] ^ x[11];
  assign t[76] = t[104] ^ x[10];
  assign t[77] = t[105] ^ x[14];
  assign t[78] = t[106] ^ x[13];
  assign t[79] = t[107] ^ x[17];
  assign t[7] = ~(t[29]);
  assign t[80] = t[108] ^ x[16];
  assign t[81] = t[109] ^ x[20];
  assign t[82] = t[110] ^ x[19];
  assign t[83] = t[111] ^ x[23];
  assign t[84] = t[112] ^ x[22];
  assign t[85] = t[113] ^ x[26];
  assign t[86] = t[114] ^ x[25];
  assign t[87] = t[115] ^ x[29];
  assign t[88] = t[116] ^ x[28];
  assign t[89] = t[117] ^ x[32];
  assign t[8] = ~(t[10]);
  assign t[90] = t[118] ^ x[31];
  assign t[91] = t[119] ^ x[35];
  assign t[92] = t[120] ^ x[34];
  assign t[93] = t[121] ^ x[38];
  assign t[94] = t[122] ^ x[37];
  assign t[95] = t[123] ^ x[41];
  assign t[96] = t[124] ^ x[40];
  assign t[97] = (x[0]);
  assign t[98] = (x[0]);
  assign t[99] = (x[3]);
  assign t[9] = ~(t[30]);
  assign y = (t[0]);
endmodule

module R2ind18(x, y);
 input [41:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[22] & t[1]);
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[15]);
  assign t[103] = (x[15]);
  assign t[104] = (x[18]);
  assign t[105] = (x[18]);
  assign t[106] = (x[21]);
  assign t[107] = (x[21]);
  assign t[108] = (x[24]);
  assign t[109] = (x[24]);
  assign t[10] = t[12] & t[13];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[30]);
  assign t[113] = (x[30]);
  assign t[114] = (x[33]);
  assign t[115] = (x[33]);
  assign t[116] = (x[36]);
  assign t[117] = (x[36]);
  assign t[118] = (x[39]);
  assign t[119] = (x[39]);
  assign t[11] = ~(t[26] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[27] & t[28]);
  assign t[16] = ~(t[29] & t[24]);
  assign t[17] = ~(t[11]);
  assign t[18] = ~(t[30] & t[21]);
  assign t[19] = ~(t[31] | t[32]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[20] = ~(t[33] | t[34]);
  assign t[21] = ~(t[35]);
  assign t[22] = (t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = t[50] ^ x[2];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[11];
  assign t[3] = ~(t[23] ^ t[24]);
  assign t[40] = t[54] ^ x[14];
  assign t[41] = t[55] ^ x[17];
  assign t[42] = t[56] ^ x[20];
  assign t[43] = t[57] ^ x[23];
  assign t[44] = t[58] ^ x[26];
  assign t[45] = t[59] ^ x[29];
  assign t[46] = t[60] ^ x[32];
  assign t[47] = t[61] ^ x[35];
  assign t[48] = t[62] ^ x[38];
  assign t[49] = t[63] ^ x[41];
  assign t[4] = ~(t[25]);
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = (t[76] & ~t[77]);
  assign t[57] = (t[78] & ~t[79]);
  assign t[58] = (t[80] & ~t[81]);
  assign t[59] = (t[82] & ~t[83]);
  assign t[5] = t[6] & t[7];
  assign t[60] = (t[84] & ~t[85]);
  assign t[61] = (t[86] & ~t[87]);
  assign t[62] = (t[88] & ~t[89]);
  assign t[63] = (t[90] & ~t[91]);
  assign t[64] = t[92] ^ x[2];
  assign t[65] = t[93] ^ x[1];
  assign t[66] = t[94] ^ x[5];
  assign t[67] = t[95] ^ x[4];
  assign t[68] = t[96] ^ x[8];
  assign t[69] = t[97] ^ x[7];
  assign t[6] = ~(t[8]);
  assign t[70] = t[98] ^ x[11];
  assign t[71] = t[99] ^ x[10];
  assign t[72] = t[100] ^ x[14];
  assign t[73] = t[101] ^ x[13];
  assign t[74] = t[102] ^ x[17];
  assign t[75] = t[103] ^ x[16];
  assign t[76] = t[104] ^ x[20];
  assign t[77] = t[105] ^ x[19];
  assign t[78] = t[106] ^ x[23];
  assign t[79] = t[107] ^ x[22];
  assign t[7] = ~(t[9]);
  assign t[80] = t[108] ^ x[26];
  assign t[81] = t[109] ^ x[25];
  assign t[82] = t[110] ^ x[29];
  assign t[83] = t[111] ^ x[28];
  assign t[84] = t[112] ^ x[32];
  assign t[85] = t[113] ^ x[31];
  assign t[86] = t[114] ^ x[35];
  assign t[87] = t[115] ^ x[34];
  assign t[88] = t[116] ^ x[38];
  assign t[89] = t[117] ^ x[37];
  assign t[8] = t[22] & t[10];
  assign t[90] = t[118] ^ x[41];
  assign t[91] = t[119] ^ x[40];
  assign t[92] = (x[0]);
  assign t[93] = (x[0]);
  assign t[94] = (x[3]);
  assign t[95] = (x[3]);
  assign t[96] = (x[6]);
  assign t[97] = (x[6]);
  assign t[98] = (x[9]);
  assign t[99] = (x[9]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind19(x, y);
 input [41:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[22] & t[1]);
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[15]);
  assign t[103] = (x[15]);
  assign t[104] = (x[18]);
  assign t[105] = (x[18]);
  assign t[106] = (x[21]);
  assign t[107] = (x[21]);
  assign t[108] = (x[24]);
  assign t[109] = (x[24]);
  assign t[10] = t[12] & t[13];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[30]);
  assign t[113] = (x[30]);
  assign t[114] = (x[33]);
  assign t[115] = (x[33]);
  assign t[116] = (x[36]);
  assign t[117] = (x[36]);
  assign t[118] = (x[39]);
  assign t[119] = (x[39]);
  assign t[11] = ~(t[26] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[27] & t[28]);
  assign t[16] = ~(t[29] & t[24]);
  assign t[17] = ~(t[11]);
  assign t[18] = ~(t[30] & t[21]);
  assign t[19] = ~(t[31] | t[32]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[20] = ~(t[33] | t[34]);
  assign t[21] = ~(t[35]);
  assign t[22] = (t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = t[50] ^ x[2];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[11];
  assign t[3] = ~(t[23] ^ t[24]);
  assign t[40] = t[54] ^ x[14];
  assign t[41] = t[55] ^ x[17];
  assign t[42] = t[56] ^ x[20];
  assign t[43] = t[57] ^ x[23];
  assign t[44] = t[58] ^ x[26];
  assign t[45] = t[59] ^ x[29];
  assign t[46] = t[60] ^ x[32];
  assign t[47] = t[61] ^ x[35];
  assign t[48] = t[62] ^ x[38];
  assign t[49] = t[63] ^ x[41];
  assign t[4] = ~(t[25]);
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = (t[76] & ~t[77]);
  assign t[57] = (t[78] & ~t[79]);
  assign t[58] = (t[80] & ~t[81]);
  assign t[59] = (t[82] & ~t[83]);
  assign t[5] = t[6] & t[7];
  assign t[60] = (t[84] & ~t[85]);
  assign t[61] = (t[86] & ~t[87]);
  assign t[62] = (t[88] & ~t[89]);
  assign t[63] = (t[90] & ~t[91]);
  assign t[64] = t[92] ^ x[2];
  assign t[65] = t[93] ^ x[1];
  assign t[66] = t[94] ^ x[5];
  assign t[67] = t[95] ^ x[4];
  assign t[68] = t[96] ^ x[8];
  assign t[69] = t[97] ^ x[7];
  assign t[6] = ~(t[8]);
  assign t[70] = t[98] ^ x[11];
  assign t[71] = t[99] ^ x[10];
  assign t[72] = t[100] ^ x[14];
  assign t[73] = t[101] ^ x[13];
  assign t[74] = t[102] ^ x[17];
  assign t[75] = t[103] ^ x[16];
  assign t[76] = t[104] ^ x[20];
  assign t[77] = t[105] ^ x[19];
  assign t[78] = t[106] ^ x[23];
  assign t[79] = t[107] ^ x[22];
  assign t[7] = ~(t[9]);
  assign t[80] = t[108] ^ x[26];
  assign t[81] = t[109] ^ x[25];
  assign t[82] = t[110] ^ x[29];
  assign t[83] = t[111] ^ x[28];
  assign t[84] = t[112] ^ x[32];
  assign t[85] = t[113] ^ x[31];
  assign t[86] = t[114] ^ x[35];
  assign t[87] = t[115] ^ x[34];
  assign t[88] = t[116] ^ x[38];
  assign t[89] = t[117] ^ x[37];
  assign t[8] = t[22] & t[10];
  assign t[90] = t[118] ^ x[41];
  assign t[91] = t[119] ^ x[40];
  assign t[92] = (x[0]);
  assign t[93] = (x[0]);
  assign t[94] = (x[3]);
  assign t[95] = (x[3]);
  assign t[96] = (x[6]);
  assign t[97] = (x[6]);
  assign t[98] = (x[9]);
  assign t[99] = (x[9]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [35:0] x;
 output y;

 wire [105:0] t;
  assign t[0] = ~(t[22] & t[1]);
  assign t[100] = (x[27]);
  assign t[101] = (x[27]);
  assign t[102] = (x[30]);
  assign t[103] = (x[30]);
  assign t[104] = (x[33]);
  assign t[105] = (x[33]);
  assign t[10] = t[12] & t[13];
  assign t[11] = ~(t[25] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[23] & t[26]);
  assign t[16] = ~(t[27] & t[24]);
  assign t[17] = ~(t[11]);
  assign t[18] = ~(t[28] & t[21]);
  assign t[19] = ~(t[29] | t[30]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[20] = ~(t[31] | t[32]);
  assign t[21] = ~(t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = (t[41]);
  assign t[2] = ~(t[5]);
  assign t[30] = (t[42]);
  assign t[31] = (t[43]);
  assign t[32] = (t[44]);
  assign t[33] = (t[45]);
  assign t[34] = t[46] ^ x[2];
  assign t[35] = t[47] ^ x[5];
  assign t[36] = t[48] ^ x[8];
  assign t[37] = t[49] ^ x[11];
  assign t[38] = t[50] ^ x[14];
  assign t[39] = t[51] ^ x[17];
  assign t[3] = ~(t[23]);
  assign t[40] = t[52] ^ x[20];
  assign t[41] = t[53] ^ x[23];
  assign t[42] = t[54] ^ x[26];
  assign t[43] = t[55] ^ x[29];
  assign t[44] = t[56] ^ x[32];
  assign t[45] = t[57] ^ x[35];
  assign t[46] = (t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[61]);
  assign t[48] = (t[62] & ~t[63]);
  assign t[49] = (t[64] & ~t[65]);
  assign t[4] = ~(t[24]);
  assign t[50] = (t[66] & ~t[67]);
  assign t[51] = (t[68] & ~t[69]);
  assign t[52] = (t[70] & ~t[71]);
  assign t[53] = (t[72] & ~t[73]);
  assign t[54] = (t[74] & ~t[75]);
  assign t[55] = (t[76] & ~t[77]);
  assign t[56] = (t[78] & ~t[79]);
  assign t[57] = (t[80] & ~t[81]);
  assign t[58] = t[82] ^ x[2];
  assign t[59] = t[83] ^ x[1];
  assign t[5] = t[6] & t[7];
  assign t[60] = t[84] ^ x[5];
  assign t[61] = t[85] ^ x[4];
  assign t[62] = t[86] ^ x[8];
  assign t[63] = t[87] ^ x[7];
  assign t[64] = t[88] ^ x[11];
  assign t[65] = t[89] ^ x[10];
  assign t[66] = t[90] ^ x[14];
  assign t[67] = t[91] ^ x[13];
  assign t[68] = t[92] ^ x[17];
  assign t[69] = t[93] ^ x[16];
  assign t[6] = ~(t[8]);
  assign t[70] = t[94] ^ x[20];
  assign t[71] = t[95] ^ x[19];
  assign t[72] = t[96] ^ x[23];
  assign t[73] = t[97] ^ x[22];
  assign t[74] = t[98] ^ x[26];
  assign t[75] = t[99] ^ x[25];
  assign t[76] = t[100] ^ x[29];
  assign t[77] = t[101] ^ x[28];
  assign t[78] = t[102] ^ x[32];
  assign t[79] = t[103] ^ x[31];
  assign t[7] = ~(t[9]);
  assign t[80] = t[104] ^ x[35];
  assign t[81] = t[105] ^ x[34];
  assign t[82] = (x[0]);
  assign t[83] = (x[0]);
  assign t[84] = (x[3]);
  assign t[85] = (x[3]);
  assign t[86] = (x[6]);
  assign t[87] = (x[6]);
  assign t[88] = (x[9]);
  assign t[89] = (x[9]);
  assign t[8] = t[22] & t[10];
  assign t[90] = (x[12]);
  assign t[91] = (x[12]);
  assign t[92] = (x[15]);
  assign t[93] = (x[15]);
  assign t[94] = (x[18]);
  assign t[95] = (x[18]);
  assign t[96] = (x[21]);
  assign t[97] = (x[21]);
  assign t[98] = (x[24]);
  assign t[99] = (x[24]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind21(x, y);
 input [35:0] x;
 output y;

 wire [105:0] t;
  assign t[0] = ~(t[22] & t[1]);
  assign t[100] = (x[27]);
  assign t[101] = (x[27]);
  assign t[102] = (x[30]);
  assign t[103] = (x[30]);
  assign t[104] = (x[33]);
  assign t[105] = (x[33]);
  assign t[10] = t[12] & t[13];
  assign t[11] = ~(t[25] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[23] & t[26]);
  assign t[16] = ~(t[27] & t[24]);
  assign t[17] = ~(t[11]);
  assign t[18] = ~(t[28] & t[21]);
  assign t[19] = ~(t[29] | t[30]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[20] = ~(t[31] | t[32]);
  assign t[21] = ~(t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = (t[41]);
  assign t[2] = ~(t[5]);
  assign t[30] = (t[42]);
  assign t[31] = (t[43]);
  assign t[32] = (t[44]);
  assign t[33] = (t[45]);
  assign t[34] = t[46] ^ x[2];
  assign t[35] = t[47] ^ x[5];
  assign t[36] = t[48] ^ x[8];
  assign t[37] = t[49] ^ x[11];
  assign t[38] = t[50] ^ x[14];
  assign t[39] = t[51] ^ x[17];
  assign t[3] = ~(t[23]);
  assign t[40] = t[52] ^ x[20];
  assign t[41] = t[53] ^ x[23];
  assign t[42] = t[54] ^ x[26];
  assign t[43] = t[55] ^ x[29];
  assign t[44] = t[56] ^ x[32];
  assign t[45] = t[57] ^ x[35];
  assign t[46] = (t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[61]);
  assign t[48] = (t[62] & ~t[63]);
  assign t[49] = (t[64] & ~t[65]);
  assign t[4] = ~(t[24]);
  assign t[50] = (t[66] & ~t[67]);
  assign t[51] = (t[68] & ~t[69]);
  assign t[52] = (t[70] & ~t[71]);
  assign t[53] = (t[72] & ~t[73]);
  assign t[54] = (t[74] & ~t[75]);
  assign t[55] = (t[76] & ~t[77]);
  assign t[56] = (t[78] & ~t[79]);
  assign t[57] = (t[80] & ~t[81]);
  assign t[58] = t[82] ^ x[2];
  assign t[59] = t[83] ^ x[1];
  assign t[5] = t[6] & t[7];
  assign t[60] = t[84] ^ x[5];
  assign t[61] = t[85] ^ x[4];
  assign t[62] = t[86] ^ x[8];
  assign t[63] = t[87] ^ x[7];
  assign t[64] = t[88] ^ x[11];
  assign t[65] = t[89] ^ x[10];
  assign t[66] = t[90] ^ x[14];
  assign t[67] = t[91] ^ x[13];
  assign t[68] = t[92] ^ x[17];
  assign t[69] = t[93] ^ x[16];
  assign t[6] = ~(t[8]);
  assign t[70] = t[94] ^ x[20];
  assign t[71] = t[95] ^ x[19];
  assign t[72] = t[96] ^ x[23];
  assign t[73] = t[97] ^ x[22];
  assign t[74] = t[98] ^ x[26];
  assign t[75] = t[99] ^ x[25];
  assign t[76] = t[100] ^ x[29];
  assign t[77] = t[101] ^ x[28];
  assign t[78] = t[102] ^ x[32];
  assign t[79] = t[103] ^ x[31];
  assign t[7] = ~(t[9]);
  assign t[80] = t[104] ^ x[35];
  assign t[81] = t[105] ^ x[34];
  assign t[82] = (x[0]);
  assign t[83] = (x[0]);
  assign t[84] = (x[3]);
  assign t[85] = (x[3]);
  assign t[86] = (x[6]);
  assign t[87] = (x[6]);
  assign t[88] = (x[9]);
  assign t[89] = (x[9]);
  assign t[8] = t[22] & t[10];
  assign t[90] = (x[12]);
  assign t[91] = (x[12]);
  assign t[92] = (x[15]);
  assign t[93] = (x[15]);
  assign t[94] = (x[18]);
  assign t[95] = (x[18]);
  assign t[96] = (x[21]);
  assign t[97] = (x[21]);
  assign t[98] = (x[24]);
  assign t[99] = (x[24]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind22(x, y);
 input [41:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[6]);
  assign t[101] = (x[9]);
  assign t[102] = (x[9]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[15]);
  assign t[106] = (x[15]);
  assign t[107] = (x[18]);
  assign t[108] = (x[18]);
  assign t[109] = (x[21]);
  assign t[10] = ~(t[12]);
  assign t[110] = (x[21]);
  assign t[111] = (x[24]);
  assign t[112] = (x[24]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[30]);
  assign t[116] = (x[30]);
  assign t[117] = (x[33]);
  assign t[118] = (x[33]);
  assign t[119] = (x[36]);
  assign t[11] = t[28] & t[13];
  assign t[120] = (x[36]);
  assign t[121] = (x[39]);
  assign t[122] = (x[39]);
  assign t[12] = ~(t[28] & t[14]);
  assign t[13] = t[15] & t[16];
  assign t[14] = ~(t[29] | t[17]);
  assign t[15] = ~(t[18] | t[19]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[25] & t[30]);
  assign t[19] = ~(t[31] & t[32]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[14]);
  assign t[21] = ~(t[33] & t[24]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5] & t[25]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = t[26] ^ t[27];
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[8];
  assign t[42] = t[56] ^ x[11];
  assign t[43] = t[57] ^ x[14];
  assign t[44] = t[58] ^ x[17];
  assign t[45] = t[59] ^ x[20];
  assign t[46] = t[60] ^ x[23];
  assign t[47] = t[61] ^ x[26];
  assign t[48] = t[62] ^ x[29];
  assign t[49] = t[63] ^ x[32];
  assign t[4] = ~(t[6] | t[7]);
  assign t[50] = t[64] ^ x[35];
  assign t[51] = t[65] ^ x[38];
  assign t[52] = t[66] ^ x[41];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = ~(t[8] | t[7]);
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[8]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[8];
  assign t[72] = t[100] ^ x[7];
  assign t[73] = t[101] ^ x[11];
  assign t[74] = t[102] ^ x[10];
  assign t[75] = t[103] ^ x[14];
  assign t[76] = t[104] ^ x[13];
  assign t[77] = t[105] ^ x[17];
  assign t[78] = t[106] ^ x[16];
  assign t[79] = t[107] ^ x[20];
  assign t[7] = ~(t[28]);
  assign t[80] = t[108] ^ x[19];
  assign t[81] = t[109] ^ x[23];
  assign t[82] = t[110] ^ x[22];
  assign t[83] = t[111] ^ x[26];
  assign t[84] = t[112] ^ x[25];
  assign t[85] = t[113] ^ x[29];
  assign t[86] = t[114] ^ x[28];
  assign t[87] = t[115] ^ x[32];
  assign t[88] = t[116] ^ x[31];
  assign t[89] = t[117] ^ x[35];
  assign t[8] = t[9] & t[10];
  assign t[90] = t[118] ^ x[34];
  assign t[91] = t[119] ^ x[38];
  assign t[92] = t[120] ^ x[37];
  assign t[93] = t[121] ^ x[41];
  assign t[94] = t[122] ^ x[40];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[6]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind23(x, y);
 input [41:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[6]);
  assign t[101] = (x[9]);
  assign t[102] = (x[9]);
  assign t[103] = (x[12]);
  assign t[104] = (x[12]);
  assign t[105] = (x[15]);
  assign t[106] = (x[15]);
  assign t[107] = (x[18]);
  assign t[108] = (x[18]);
  assign t[109] = (x[21]);
  assign t[10] = ~(t[12]);
  assign t[110] = (x[21]);
  assign t[111] = (x[24]);
  assign t[112] = (x[24]);
  assign t[113] = (x[27]);
  assign t[114] = (x[27]);
  assign t[115] = (x[30]);
  assign t[116] = (x[30]);
  assign t[117] = (x[33]);
  assign t[118] = (x[33]);
  assign t[119] = (x[36]);
  assign t[11] = t[28] & t[13];
  assign t[120] = (x[36]);
  assign t[121] = (x[39]);
  assign t[122] = (x[39]);
  assign t[12] = ~(t[28] & t[14]);
  assign t[13] = t[15] & t[16];
  assign t[14] = ~(t[29] | t[17]);
  assign t[15] = ~(t[18] | t[19]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[22] & t[23]);
  assign t[18] = ~(t[25] & t[30]);
  assign t[19] = ~(t[31] & t[32]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[14]);
  assign t[21] = ~(t[33] & t[24]);
  assign t[22] = ~(t[34] | t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5] & t[25]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = t[26] ^ t[27];
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[8];
  assign t[42] = t[56] ^ x[11];
  assign t[43] = t[57] ^ x[14];
  assign t[44] = t[58] ^ x[17];
  assign t[45] = t[59] ^ x[20];
  assign t[46] = t[60] ^ x[23];
  assign t[47] = t[61] ^ x[26];
  assign t[48] = t[62] ^ x[29];
  assign t[49] = t[63] ^ x[32];
  assign t[4] = ~(t[6] | t[7]);
  assign t[50] = t[64] ^ x[35];
  assign t[51] = t[65] ^ x[38];
  assign t[52] = t[66] ^ x[41];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = ~(t[8] | t[7]);
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[8]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[8];
  assign t[72] = t[100] ^ x[7];
  assign t[73] = t[101] ^ x[11];
  assign t[74] = t[102] ^ x[10];
  assign t[75] = t[103] ^ x[14];
  assign t[76] = t[104] ^ x[13];
  assign t[77] = t[105] ^ x[17];
  assign t[78] = t[106] ^ x[16];
  assign t[79] = t[107] ^ x[20];
  assign t[7] = ~(t[28]);
  assign t[80] = t[108] ^ x[19];
  assign t[81] = t[109] ^ x[23];
  assign t[82] = t[110] ^ x[22];
  assign t[83] = t[111] ^ x[26];
  assign t[84] = t[112] ^ x[25];
  assign t[85] = t[113] ^ x[29];
  assign t[86] = t[114] ^ x[28];
  assign t[87] = t[115] ^ x[32];
  assign t[88] = t[116] ^ x[31];
  assign t[89] = t[117] ^ x[35];
  assign t[8] = t[9] & t[10];
  assign t[90] = t[118] ^ x[34];
  assign t[91] = t[119] ^ x[38];
  assign t[92] = t[120] ^ x[37];
  assign t[93] = t[121] ^ x[41];
  assign t[94] = t[122] ^ x[40];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[6]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind24(x, y);
 input [41:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[22] & t[1]);
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[15]);
  assign t[103] = (x[15]);
  assign t[104] = (x[18]);
  assign t[105] = (x[18]);
  assign t[106] = (x[21]);
  assign t[107] = (x[21]);
  assign t[108] = (x[24]);
  assign t[109] = (x[24]);
  assign t[10] = t[12] & t[13];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[30]);
  assign t[113] = (x[30]);
  assign t[114] = (x[33]);
  assign t[115] = (x[33]);
  assign t[116] = (x[36]);
  assign t[117] = (x[36]);
  assign t[118] = (x[39]);
  assign t[119] = (x[39]);
  assign t[11] = ~(t[25] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[11]);
  assign t[18] = ~(t[30] & t[21]);
  assign t[19] = ~(t[31] | t[32]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[20] = ~(t[33] | t[34]);
  assign t[21] = ~(t[35]);
  assign t[22] = (t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = t[50] ^ x[2];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[11];
  assign t[3] = ~(t[23]);
  assign t[40] = t[54] ^ x[14];
  assign t[41] = t[55] ^ x[17];
  assign t[42] = t[56] ^ x[20];
  assign t[43] = t[57] ^ x[23];
  assign t[44] = t[58] ^ x[26];
  assign t[45] = t[59] ^ x[29];
  assign t[46] = t[60] ^ x[32];
  assign t[47] = t[61] ^ x[35];
  assign t[48] = t[62] ^ x[38];
  assign t[49] = t[63] ^ x[41];
  assign t[4] = ~(t[24]);
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = (t[76] & ~t[77]);
  assign t[57] = (t[78] & ~t[79]);
  assign t[58] = (t[80] & ~t[81]);
  assign t[59] = (t[82] & ~t[83]);
  assign t[5] = t[6] & t[7];
  assign t[60] = (t[84] & ~t[85]);
  assign t[61] = (t[86] & ~t[87]);
  assign t[62] = (t[88] & ~t[89]);
  assign t[63] = (t[90] & ~t[91]);
  assign t[64] = t[92] ^ x[2];
  assign t[65] = t[93] ^ x[1];
  assign t[66] = t[94] ^ x[5];
  assign t[67] = t[95] ^ x[4];
  assign t[68] = t[96] ^ x[8];
  assign t[69] = t[97] ^ x[7];
  assign t[6] = ~(t[8]);
  assign t[70] = t[98] ^ x[11];
  assign t[71] = t[99] ^ x[10];
  assign t[72] = t[100] ^ x[14];
  assign t[73] = t[101] ^ x[13];
  assign t[74] = t[102] ^ x[17];
  assign t[75] = t[103] ^ x[16];
  assign t[76] = t[104] ^ x[20];
  assign t[77] = t[105] ^ x[19];
  assign t[78] = t[106] ^ x[23];
  assign t[79] = t[107] ^ x[22];
  assign t[7] = ~(t[9]);
  assign t[80] = t[108] ^ x[26];
  assign t[81] = t[109] ^ x[25];
  assign t[82] = t[110] ^ x[29];
  assign t[83] = t[111] ^ x[28];
  assign t[84] = t[112] ^ x[32];
  assign t[85] = t[113] ^ x[31];
  assign t[86] = t[114] ^ x[35];
  assign t[87] = t[115] ^ x[34];
  assign t[88] = t[116] ^ x[38];
  assign t[89] = t[117] ^ x[37];
  assign t[8] = t[22] & t[10];
  assign t[90] = t[118] ^ x[41];
  assign t[91] = t[119] ^ x[40];
  assign t[92] = (x[0]);
  assign t[93] = (x[0]);
  assign t[94] = (x[3]);
  assign t[95] = (x[3]);
  assign t[96] = (x[6]);
  assign t[97] = (x[6]);
  assign t[98] = (x[9]);
  assign t[99] = (x[9]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [41:0] x;
 output y;

 wire [119:0] t;
  assign t[0] = ~(t[22] & t[1]);
  assign t[100] = (x[12]);
  assign t[101] = (x[12]);
  assign t[102] = (x[15]);
  assign t[103] = (x[15]);
  assign t[104] = (x[18]);
  assign t[105] = (x[18]);
  assign t[106] = (x[21]);
  assign t[107] = (x[21]);
  assign t[108] = (x[24]);
  assign t[109] = (x[24]);
  assign t[10] = t[12] & t[13];
  assign t[110] = (x[27]);
  assign t[111] = (x[27]);
  assign t[112] = (x[30]);
  assign t[113] = (x[30]);
  assign t[114] = (x[33]);
  assign t[115] = (x[33]);
  assign t[116] = (x[36]);
  assign t[117] = (x[36]);
  assign t[118] = (x[39]);
  assign t[119] = (x[39]);
  assign t[11] = ~(t[25] | t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(t[19] & t[20]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[28] & t[29]);
  assign t[17] = ~(t[11]);
  assign t[18] = ~(t[30] & t[21]);
  assign t[19] = ~(t[31] | t[32]);
  assign t[1] = t[2] ? t[4] : t[3];
  assign t[20] = ~(t[33] | t[34]);
  assign t[21] = ~(t[35]);
  assign t[22] = (t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = t[50] ^ x[2];
  assign t[37] = t[51] ^ x[5];
  assign t[38] = t[52] ^ x[8];
  assign t[39] = t[53] ^ x[11];
  assign t[3] = ~(t[23]);
  assign t[40] = t[54] ^ x[14];
  assign t[41] = t[55] ^ x[17];
  assign t[42] = t[56] ^ x[20];
  assign t[43] = t[57] ^ x[23];
  assign t[44] = t[58] ^ x[26];
  assign t[45] = t[59] ^ x[29];
  assign t[46] = t[60] ^ x[32];
  assign t[47] = t[61] ^ x[35];
  assign t[48] = t[62] ^ x[38];
  assign t[49] = t[63] ^ x[41];
  assign t[4] = ~(t[24]);
  assign t[50] = (t[64] & ~t[65]);
  assign t[51] = (t[66] & ~t[67]);
  assign t[52] = (t[68] & ~t[69]);
  assign t[53] = (t[70] & ~t[71]);
  assign t[54] = (t[72] & ~t[73]);
  assign t[55] = (t[74] & ~t[75]);
  assign t[56] = (t[76] & ~t[77]);
  assign t[57] = (t[78] & ~t[79]);
  assign t[58] = (t[80] & ~t[81]);
  assign t[59] = (t[82] & ~t[83]);
  assign t[5] = t[6] & t[7];
  assign t[60] = (t[84] & ~t[85]);
  assign t[61] = (t[86] & ~t[87]);
  assign t[62] = (t[88] & ~t[89]);
  assign t[63] = (t[90] & ~t[91]);
  assign t[64] = t[92] ^ x[2];
  assign t[65] = t[93] ^ x[1];
  assign t[66] = t[94] ^ x[5];
  assign t[67] = t[95] ^ x[4];
  assign t[68] = t[96] ^ x[8];
  assign t[69] = t[97] ^ x[7];
  assign t[6] = ~(t[8]);
  assign t[70] = t[98] ^ x[11];
  assign t[71] = t[99] ^ x[10];
  assign t[72] = t[100] ^ x[14];
  assign t[73] = t[101] ^ x[13];
  assign t[74] = t[102] ^ x[17];
  assign t[75] = t[103] ^ x[16];
  assign t[76] = t[104] ^ x[20];
  assign t[77] = t[105] ^ x[19];
  assign t[78] = t[106] ^ x[23];
  assign t[79] = t[107] ^ x[22];
  assign t[7] = ~(t[9]);
  assign t[80] = t[108] ^ x[26];
  assign t[81] = t[109] ^ x[25];
  assign t[82] = t[110] ^ x[29];
  assign t[83] = t[111] ^ x[28];
  assign t[84] = t[112] ^ x[32];
  assign t[85] = t[113] ^ x[31];
  assign t[86] = t[114] ^ x[35];
  assign t[87] = t[115] ^ x[34];
  assign t[88] = t[116] ^ x[38];
  assign t[89] = t[117] ^ x[37];
  assign t[8] = t[22] & t[10];
  assign t[90] = t[118] ^ x[41];
  assign t[91] = t[119] ^ x[40];
  assign t[92] = (x[0]);
  assign t[93] = (x[0]);
  assign t[94] = (x[3]);
  assign t[95] = (x[3]);
  assign t[96] = (x[6]);
  assign t[97] = (x[6]);
  assign t[98] = (x[9]);
  assign t[99] = (x[9]);
  assign t[9] = ~(t[22] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind26(x, y);
 input [35:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[100] = (x[33]);
  assign t[101] = (x[33]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[22] & t[23]);
  assign t[13] = ~(t[24] & t[25]);
  assign t[14] = ~(t[7]);
  assign t[15] = ~(t[18] & t[5]);
  assign t[16] = ~(t[26] | t[27]);
  assign t[17] = ~(t[28] | t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = (t[41]);
  assign t[2] = ~(t[4] & ~t[5]);
  assign t[30] = t[42] ^ x[2];
  assign t[31] = t[43] ^ x[5];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[11];
  assign t[34] = t[46] ^ x[14];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[20];
  assign t[37] = t[49] ^ x[23];
  assign t[38] = t[50] ^ x[26];
  assign t[39] = t[51] ^ x[29];
  assign t[3] = t[19] & t[6];
  assign t[40] = t[52] ^ x[32];
  assign t[41] = t[53] ^ x[35];
  assign t[42] = (t[54] & ~t[55]);
  assign t[43] = (t[56] & ~t[57]);
  assign t[44] = (t[58] & ~t[59]);
  assign t[45] = (t[60] & ~t[61]);
  assign t[46] = (t[62] & ~t[63]);
  assign t[47] = (t[64] & ~t[65]);
  assign t[48] = (t[66] & ~t[67]);
  assign t[49] = (t[68] & ~t[69]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[50] = (t[70] & ~t[71]);
  assign t[51] = (t[72] & ~t[73]);
  assign t[52] = (t[74] & ~t[75]);
  assign t[53] = (t[76] & ~t[77]);
  assign t[54] = t[78] ^ x[2];
  assign t[55] = t[79] ^ x[1];
  assign t[56] = t[80] ^ x[5];
  assign t[57] = t[81] ^ x[4];
  assign t[58] = t[82] ^ x[8];
  assign t[59] = t[83] ^ x[7];
  assign t[5] = ~(t[20]);
  assign t[60] = t[84] ^ x[11];
  assign t[61] = t[85] ^ x[10];
  assign t[62] = t[86] ^ x[14];
  assign t[63] = t[87] ^ x[13];
  assign t[64] = t[88] ^ x[17];
  assign t[65] = t[89] ^ x[16];
  assign t[66] = t[90] ^ x[20];
  assign t[67] = t[91] ^ x[19];
  assign t[68] = t[92] ^ x[23];
  assign t[69] = t[93] ^ x[22];
  assign t[6] = t[9] & t[10];
  assign t[70] = t[94] ^ x[26];
  assign t[71] = t[95] ^ x[25];
  assign t[72] = t[96] ^ x[29];
  assign t[73] = t[97] ^ x[28];
  assign t[74] = t[98] ^ x[32];
  assign t[75] = t[99] ^ x[31];
  assign t[76] = t[100] ^ x[35];
  assign t[77] = t[101] ^ x[34];
  assign t[78] = (x[0]);
  assign t[79] = (x[0]);
  assign t[7] = ~(t[21] | t[11]);
  assign t[80] = (x[3]);
  assign t[81] = (x[3]);
  assign t[82] = (x[6]);
  assign t[83] = (x[6]);
  assign t[84] = (x[9]);
  assign t[85] = (x[9]);
  assign t[86] = (x[12]);
  assign t[87] = (x[12]);
  assign t[88] = (x[15]);
  assign t[89] = (x[15]);
  assign t[8] = ~(t[19]);
  assign t[90] = (x[18]);
  assign t[91] = (x[18]);
  assign t[92] = (x[21]);
  assign t[93] = (x[21]);
  assign t[94] = (x[24]);
  assign t[95] = (x[24]);
  assign t[96] = (x[27]);
  assign t[97] = (x[27]);
  assign t[98] = (x[30]);
  assign t[99] = (x[30]);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind27(x, y);
 input [35:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[100] = (x[33]);
  assign t[101] = (x[33]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(t[16] & t[17]);
  assign t[12] = ~(t[22] & t[23]);
  assign t[13] = ~(t[24] & t[25]);
  assign t[14] = ~(t[7]);
  assign t[15] = ~(t[18] & t[5]);
  assign t[16] = ~(t[26] | t[27]);
  assign t[17] = ~(t[28] | t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = (t[41]);
  assign t[2] = ~(t[4] & ~t[5]);
  assign t[30] = t[42] ^ x[2];
  assign t[31] = t[43] ^ x[5];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[11];
  assign t[34] = t[46] ^ x[14];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[20];
  assign t[37] = t[49] ^ x[23];
  assign t[38] = t[50] ^ x[26];
  assign t[39] = t[51] ^ x[29];
  assign t[3] = t[19] & t[6];
  assign t[40] = t[52] ^ x[32];
  assign t[41] = t[53] ^ x[35];
  assign t[42] = (t[54] & ~t[55]);
  assign t[43] = (t[56] & ~t[57]);
  assign t[44] = (t[58] & ~t[59]);
  assign t[45] = (t[60] & ~t[61]);
  assign t[46] = (t[62] & ~t[63]);
  assign t[47] = (t[64] & ~t[65]);
  assign t[48] = (t[66] & ~t[67]);
  assign t[49] = (t[68] & ~t[69]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[50] = (t[70] & ~t[71]);
  assign t[51] = (t[72] & ~t[73]);
  assign t[52] = (t[74] & ~t[75]);
  assign t[53] = (t[76] & ~t[77]);
  assign t[54] = t[78] ^ x[2];
  assign t[55] = t[79] ^ x[1];
  assign t[56] = t[80] ^ x[5];
  assign t[57] = t[81] ^ x[4];
  assign t[58] = t[82] ^ x[8];
  assign t[59] = t[83] ^ x[7];
  assign t[5] = ~(t[20]);
  assign t[60] = t[84] ^ x[11];
  assign t[61] = t[85] ^ x[10];
  assign t[62] = t[86] ^ x[14];
  assign t[63] = t[87] ^ x[13];
  assign t[64] = t[88] ^ x[17];
  assign t[65] = t[89] ^ x[16];
  assign t[66] = t[90] ^ x[20];
  assign t[67] = t[91] ^ x[19];
  assign t[68] = t[92] ^ x[23];
  assign t[69] = t[93] ^ x[22];
  assign t[6] = t[9] & t[10];
  assign t[70] = t[94] ^ x[26];
  assign t[71] = t[95] ^ x[25];
  assign t[72] = t[96] ^ x[29];
  assign t[73] = t[97] ^ x[28];
  assign t[74] = t[98] ^ x[32];
  assign t[75] = t[99] ^ x[31];
  assign t[76] = t[100] ^ x[35];
  assign t[77] = t[101] ^ x[34];
  assign t[78] = (x[0]);
  assign t[79] = (x[0]);
  assign t[7] = ~(t[21] | t[11]);
  assign t[80] = (x[3]);
  assign t[81] = (x[3]);
  assign t[82] = (x[6]);
  assign t[83] = (x[6]);
  assign t[84] = (x[9]);
  assign t[85] = (x[9]);
  assign t[86] = (x[12]);
  assign t[87] = (x[12]);
  assign t[88] = (x[15]);
  assign t[89] = (x[15]);
  assign t[8] = ~(t[19]);
  assign t[90] = (x[18]);
  assign t[91] = (x[18]);
  assign t[92] = (x[21]);
  assign t[93] = (x[21]);
  assign t[94] = (x[24]);
  assign t[95] = (x[24]);
  assign t[96] = (x[27]);
  assign t[97] = (x[27]);
  assign t[98] = (x[30]);
  assign t[99] = (x[30]);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind28(x, y);
 input [35:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[100] = (x[33]);
  assign t[101] = (x[33]);
  assign t[10] = ~(t[15] & t[16]);
  assign t[11] = ~(t[22] & t[23]);
  assign t[12] = ~(t[24] & t[25]);
  assign t[13] = ~(t[6]);
  assign t[14] = ~(t[19] & t[17]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[18]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = (t[41]);
  assign t[2] = t[4] & t[19];
  assign t[30] = t[42] ^ x[2];
  assign t[31] = t[43] ^ x[5];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[11];
  assign t[34] = t[46] ^ x[14];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[20];
  assign t[37] = t[49] ^ x[23];
  assign t[38] = t[50] ^ x[26];
  assign t[39] = t[51] ^ x[29];
  assign t[3] = t[20] & t[5];
  assign t[40] = t[52] ^ x[32];
  assign t[41] = t[53] ^ x[35];
  assign t[42] = (t[54] & ~t[55]);
  assign t[43] = (t[56] & ~t[57]);
  assign t[44] = (t[58] & ~t[59]);
  assign t[45] = (t[60] & ~t[61]);
  assign t[46] = (t[62] & ~t[63]);
  assign t[47] = (t[64] & ~t[65]);
  assign t[48] = (t[66] & ~t[67]);
  assign t[49] = (t[68] & ~t[69]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[50] = (t[70] & ~t[71]);
  assign t[51] = (t[72] & ~t[73]);
  assign t[52] = (t[74] & ~t[75]);
  assign t[53] = (t[76] & ~t[77]);
  assign t[54] = t[78] ^ x[2];
  assign t[55] = t[79] ^ x[1];
  assign t[56] = t[80] ^ x[5];
  assign t[57] = t[81] ^ x[4];
  assign t[58] = t[82] ^ x[8];
  assign t[59] = t[83] ^ x[7];
  assign t[5] = t[8] & t[9];
  assign t[60] = t[84] ^ x[11];
  assign t[61] = t[85] ^ x[10];
  assign t[62] = t[86] ^ x[14];
  assign t[63] = t[87] ^ x[13];
  assign t[64] = t[88] ^ x[17];
  assign t[65] = t[89] ^ x[16];
  assign t[66] = t[90] ^ x[20];
  assign t[67] = t[91] ^ x[19];
  assign t[68] = t[92] ^ x[23];
  assign t[69] = t[93] ^ x[22];
  assign t[6] = ~(t[21] | t[10]);
  assign t[70] = t[94] ^ x[26];
  assign t[71] = t[95] ^ x[25];
  assign t[72] = t[96] ^ x[29];
  assign t[73] = t[97] ^ x[28];
  assign t[74] = t[98] ^ x[32];
  assign t[75] = t[99] ^ x[31];
  assign t[76] = t[100] ^ x[35];
  assign t[77] = t[101] ^ x[34];
  assign t[78] = (x[0]);
  assign t[79] = (x[0]);
  assign t[7] = ~(t[20]);
  assign t[80] = (x[3]);
  assign t[81] = (x[3]);
  assign t[82] = (x[6]);
  assign t[83] = (x[6]);
  assign t[84] = (x[9]);
  assign t[85] = (x[9]);
  assign t[86] = (x[12]);
  assign t[87] = (x[12]);
  assign t[88] = (x[15]);
  assign t[89] = (x[15]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[90] = (x[18]);
  assign t[91] = (x[18]);
  assign t[92] = (x[21]);
  assign t[93] = (x[21]);
  assign t[94] = (x[24]);
  assign t[95] = (x[24]);
  assign t[96] = (x[27]);
  assign t[97] = (x[27]);
  assign t[98] = (x[30]);
  assign t[99] = (x[30]);
  assign t[9] = ~(t[13] | t[14]);
  assign y = (t[0]);
endmodule

module R2ind29(x, y);
 input [35:0] x;
 output y;

 wire [101:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[100] = (x[33]);
  assign t[101] = (x[33]);
  assign t[10] = ~(t[15] & t[16]);
  assign t[11] = ~(t[22] & t[23]);
  assign t[12] = ~(t[24] & t[25]);
  assign t[13] = ~(t[6]);
  assign t[14] = ~(t[19] & t[17]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = ~(t[28] | t[29]);
  assign t[17] = ~(t[18]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = (t[41]);
  assign t[2] = t[4] & t[19];
  assign t[30] = t[42] ^ x[2];
  assign t[31] = t[43] ^ x[5];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[11];
  assign t[34] = t[46] ^ x[14];
  assign t[35] = t[47] ^ x[17];
  assign t[36] = t[48] ^ x[20];
  assign t[37] = t[49] ^ x[23];
  assign t[38] = t[50] ^ x[26];
  assign t[39] = t[51] ^ x[29];
  assign t[3] = t[20] & t[5];
  assign t[40] = t[52] ^ x[32];
  assign t[41] = t[53] ^ x[35];
  assign t[42] = (t[54] & ~t[55]);
  assign t[43] = (t[56] & ~t[57]);
  assign t[44] = (t[58] & ~t[59]);
  assign t[45] = (t[60] & ~t[61]);
  assign t[46] = (t[62] & ~t[63]);
  assign t[47] = (t[64] & ~t[65]);
  assign t[48] = (t[66] & ~t[67]);
  assign t[49] = (t[68] & ~t[69]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[50] = (t[70] & ~t[71]);
  assign t[51] = (t[72] & ~t[73]);
  assign t[52] = (t[74] & ~t[75]);
  assign t[53] = (t[76] & ~t[77]);
  assign t[54] = t[78] ^ x[2];
  assign t[55] = t[79] ^ x[1];
  assign t[56] = t[80] ^ x[5];
  assign t[57] = t[81] ^ x[4];
  assign t[58] = t[82] ^ x[8];
  assign t[59] = t[83] ^ x[7];
  assign t[5] = t[8] & t[9];
  assign t[60] = t[84] ^ x[11];
  assign t[61] = t[85] ^ x[10];
  assign t[62] = t[86] ^ x[14];
  assign t[63] = t[87] ^ x[13];
  assign t[64] = t[88] ^ x[17];
  assign t[65] = t[89] ^ x[16];
  assign t[66] = t[90] ^ x[20];
  assign t[67] = t[91] ^ x[19];
  assign t[68] = t[92] ^ x[23];
  assign t[69] = t[93] ^ x[22];
  assign t[6] = ~(t[21] | t[10]);
  assign t[70] = t[94] ^ x[26];
  assign t[71] = t[95] ^ x[25];
  assign t[72] = t[96] ^ x[29];
  assign t[73] = t[97] ^ x[28];
  assign t[74] = t[98] ^ x[32];
  assign t[75] = t[99] ^ x[31];
  assign t[76] = t[100] ^ x[35];
  assign t[77] = t[101] ^ x[34];
  assign t[78] = (x[0]);
  assign t[79] = (x[0]);
  assign t[7] = ~(t[20]);
  assign t[80] = (x[3]);
  assign t[81] = (x[3]);
  assign t[82] = (x[6]);
  assign t[83] = (x[6]);
  assign t[84] = (x[9]);
  assign t[85] = (x[9]);
  assign t[86] = (x[12]);
  assign t[87] = (x[12]);
  assign t[88] = (x[15]);
  assign t[89] = (x[15]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[90] = (x[18]);
  assign t[91] = (x[18]);
  assign t[92] = (x[21]);
  assign t[93] = (x[21]);
  assign t[94] = (x[24]);
  assign t[95] = (x[24]);
  assign t[96] = (x[27]);
  assign t[97] = (x[27]);
  assign t[98] = (x[30]);
  assign t[99] = (x[30]);
  assign t[9] = ~(t[13] | t[14]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [35:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = t[1] ? t[2] : t[17];
  assign t[100] = (x[33]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[24] & t[13]);
  assign t[12] = ~(t[25] | t[14]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[15] & t[16]);
  assign t[15] = ~(t[17] | t[27]);
  assign t[16] = ~(t[28] | t[19]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = t[41] ^ x[2];
  assign t[2] = ~(t[18] & ~t[4]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[8];
  assign t[32] = t[44] ^ x[11];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[20];
  assign t[36] = t[48] ^ x[23];
  assign t[37] = t[49] ^ x[26];
  assign t[38] = t[50] ^ x[29];
  assign t[39] = t[51] ^ x[32];
  assign t[3] = t[18] & t[5];
  assign t[40] = t[52] ^ x[35];
  assign t[41] = (t[53] & ~t[54]);
  assign t[42] = (t[55] & ~t[56]);
  assign t[43] = (t[57] & ~t[58]);
  assign t[44] = (t[59] & ~t[60]);
  assign t[45] = (t[61] & ~t[62]);
  assign t[46] = (t[63] & ~t[64]);
  assign t[47] = (t[65] & ~t[66]);
  assign t[48] = (t[67] & ~t[68]);
  assign t[49] = (t[69] & ~t[70]);
  assign t[4] = ~(t[19] ^ t[17]);
  assign t[50] = (t[71] & ~t[72]);
  assign t[51] = (t[73] & ~t[74]);
  assign t[52] = (t[75] & ~t[76]);
  assign t[53] = t[77] ^ x[2];
  assign t[54] = t[78] ^ x[1];
  assign t[55] = t[79] ^ x[5];
  assign t[56] = t[80] ^ x[4];
  assign t[57] = t[81] ^ x[8];
  assign t[58] = t[82] ^ x[7];
  assign t[59] = t[83] ^ x[11];
  assign t[5] = t[6] & t[7];
  assign t[60] = t[84] ^ x[10];
  assign t[61] = t[85] ^ x[14];
  assign t[62] = t[86] ^ x[13];
  assign t[63] = t[87] ^ x[17];
  assign t[64] = t[88] ^ x[16];
  assign t[65] = t[89] ^ x[20];
  assign t[66] = t[90] ^ x[19];
  assign t[67] = t[91] ^ x[23];
  assign t[68] = t[92] ^ x[22];
  assign t[69] = t[93] ^ x[26];
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = t[94] ^ x[25];
  assign t[71] = t[95] ^ x[29];
  assign t[72] = t[96] ^ x[28];
  assign t[73] = t[97] ^ x[32];
  assign t[74] = t[98] ^ x[31];
  assign t[75] = t[99] ^ x[35];
  assign t[76] = t[100] ^ x[34];
  assign t[77] = (x[0]);
  assign t[78] = (x[0]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[80] = (x[3]);
  assign t[81] = (x[6]);
  assign t[82] = (x[6]);
  assign t[83] = (x[9]);
  assign t[84] = (x[9]);
  assign t[85] = (x[12]);
  assign t[86] = (x[12]);
  assign t[87] = (x[15]);
  assign t[88] = (x[15]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[20] & t[21]);
  assign t[90] = (x[18]);
  assign t[91] = (x[21]);
  assign t[92] = (x[21]);
  assign t[93] = (x[24]);
  assign t[94] = (x[24]);
  assign t[95] = (x[27]);
  assign t[96] = (x[27]);
  assign t[97] = (x[30]);
  assign t[98] = (x[30]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[22] & t[23]);
  assign y = (t[0]);
endmodule

module R2ind31(x, y);
 input [35:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = t[1] ? t[2] : t[17];
  assign t[100] = (x[33]);
  assign t[10] = ~(t[12]);
  assign t[11] = ~(t[24] & t[13]);
  assign t[12] = ~(t[25] | t[14]);
  assign t[13] = ~(t[26]);
  assign t[14] = ~(t[15] & t[16]);
  assign t[15] = ~(t[17] | t[27]);
  assign t[16] = ~(t[28] | t[19]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = t[41] ^ x[2];
  assign t[2] = ~(t[18] & ~t[4]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[8];
  assign t[32] = t[44] ^ x[11];
  assign t[33] = t[45] ^ x[14];
  assign t[34] = t[46] ^ x[17];
  assign t[35] = t[47] ^ x[20];
  assign t[36] = t[48] ^ x[23];
  assign t[37] = t[49] ^ x[26];
  assign t[38] = t[50] ^ x[29];
  assign t[39] = t[51] ^ x[32];
  assign t[3] = t[18] & t[5];
  assign t[40] = t[52] ^ x[35];
  assign t[41] = (t[53] & ~t[54]);
  assign t[42] = (t[55] & ~t[56]);
  assign t[43] = (t[57] & ~t[58]);
  assign t[44] = (t[59] & ~t[60]);
  assign t[45] = (t[61] & ~t[62]);
  assign t[46] = (t[63] & ~t[64]);
  assign t[47] = (t[65] & ~t[66]);
  assign t[48] = (t[67] & ~t[68]);
  assign t[49] = (t[69] & ~t[70]);
  assign t[4] = ~(t[19] ^ t[17]);
  assign t[50] = (t[71] & ~t[72]);
  assign t[51] = (t[73] & ~t[74]);
  assign t[52] = (t[75] & ~t[76]);
  assign t[53] = t[77] ^ x[2];
  assign t[54] = t[78] ^ x[1];
  assign t[55] = t[79] ^ x[5];
  assign t[56] = t[80] ^ x[4];
  assign t[57] = t[81] ^ x[8];
  assign t[58] = t[82] ^ x[7];
  assign t[59] = t[83] ^ x[11];
  assign t[5] = t[6] & t[7];
  assign t[60] = t[84] ^ x[10];
  assign t[61] = t[85] ^ x[14];
  assign t[62] = t[86] ^ x[13];
  assign t[63] = t[87] ^ x[17];
  assign t[64] = t[88] ^ x[16];
  assign t[65] = t[89] ^ x[20];
  assign t[66] = t[90] ^ x[19];
  assign t[67] = t[91] ^ x[23];
  assign t[68] = t[92] ^ x[22];
  assign t[69] = t[93] ^ x[26];
  assign t[6] = ~(t[8] | t[9]);
  assign t[70] = t[94] ^ x[25];
  assign t[71] = t[95] ^ x[29];
  assign t[72] = t[96] ^ x[28];
  assign t[73] = t[97] ^ x[32];
  assign t[74] = t[98] ^ x[31];
  assign t[75] = t[99] ^ x[35];
  assign t[76] = t[100] ^ x[34];
  assign t[77] = (x[0]);
  assign t[78] = (x[0]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[80] = (x[3]);
  assign t[81] = (x[6]);
  assign t[82] = (x[6]);
  assign t[83] = (x[9]);
  assign t[84] = (x[9]);
  assign t[85] = (x[12]);
  assign t[86] = (x[12]);
  assign t[87] = (x[15]);
  assign t[88] = (x[15]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[20] & t[21]);
  assign t[90] = (x[18]);
  assign t[91] = (x[21]);
  assign t[92] = (x[21]);
  assign t[93] = (x[24]);
  assign t[94] = (x[24]);
  assign t[95] = (x[27]);
  assign t[96] = (x[27]);
  assign t[97] = (x[30]);
  assign t[98] = (x[30]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[22] & t[23]);
  assign y = (t[0]);
endmodule

module R2ind32(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[16] | t[13]);
  assign t[12] = ~(t[24]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[18] | t[25]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = t[17] & t[18];
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[17];
  assign t[34] = t[46] ^ x[20];
  assign t[35] = t[47] ^ x[23];
  assign t[36] = t[48] ^ x[26];
  assign t[37] = t[49] ^ x[29];
  assign t[38] = t[50] ^ x[32];
  assign t[39] = t[51] ^ x[35];
  assign t[3] = t[17] & t[4];
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[61]);
  assign t[45] = (t[62] & ~t[63]);
  assign t[46] = (t[64] & ~t[65]);
  assign t[47] = (t[66] & ~t[67]);
  assign t[48] = (t[68] & ~t[69]);
  assign t[49] = (t[70] & ~t[71]);
  assign t[4] = t[5] & t[6];
  assign t[50] = (t[72] & ~t[73]);
  assign t[51] = (t[74] & ~t[75]);
  assign t[52] = t[76] ^ x[2];
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[5];
  assign t[55] = t[79] ^ x[4];
  assign t[56] = t[80] ^ x[8];
  assign t[57] = t[81] ^ x[7];
  assign t[58] = t[82] ^ x[11];
  assign t[59] = t[83] ^ x[10];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[84] ^ x[14];
  assign t[61] = t[85] ^ x[13];
  assign t[62] = t[86] ^ x[17];
  assign t[63] = t[87] ^ x[16];
  assign t[64] = t[88] ^ x[20];
  assign t[65] = t[89] ^ x[19];
  assign t[66] = t[90] ^ x[23];
  assign t[67] = t[91] ^ x[22];
  assign t[68] = t[92] ^ x[26];
  assign t[69] = t[93] ^ x[25];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[94] ^ x[29];
  assign t[71] = t[95] ^ x[28];
  assign t[72] = t[96] ^ x[32];
  assign t[73] = t[97] ^ x[31];
  assign t[74] = t[98] ^ x[35];
  assign t[75] = t[99] ^ x[34];
  assign t[76] = (x[0]);
  assign t[77] = (x[0]);
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind33(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[16] | t[13]);
  assign t[12] = ~(t[24]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[18] | t[25]);
  assign t[15] = ~(t[26] | t[27]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = t[17] & t[18];
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[17];
  assign t[34] = t[46] ^ x[20];
  assign t[35] = t[47] ^ x[23];
  assign t[36] = t[48] ^ x[26];
  assign t[37] = t[49] ^ x[29];
  assign t[38] = t[50] ^ x[32];
  assign t[39] = t[51] ^ x[35];
  assign t[3] = t[17] & t[4];
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[61]);
  assign t[45] = (t[62] & ~t[63]);
  assign t[46] = (t[64] & ~t[65]);
  assign t[47] = (t[66] & ~t[67]);
  assign t[48] = (t[68] & ~t[69]);
  assign t[49] = (t[70] & ~t[71]);
  assign t[4] = t[5] & t[6];
  assign t[50] = (t[72] & ~t[73]);
  assign t[51] = (t[74] & ~t[75]);
  assign t[52] = t[76] ^ x[2];
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[5];
  assign t[55] = t[79] ^ x[4];
  assign t[56] = t[80] ^ x[8];
  assign t[57] = t[81] ^ x[7];
  assign t[58] = t[82] ^ x[11];
  assign t[59] = t[83] ^ x[10];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[84] ^ x[14];
  assign t[61] = t[85] ^ x[13];
  assign t[62] = t[86] ^ x[17];
  assign t[63] = t[87] ^ x[16];
  assign t[64] = t[88] ^ x[20];
  assign t[65] = t[89] ^ x[19];
  assign t[66] = t[90] ^ x[23];
  assign t[67] = t[91] ^ x[22];
  assign t[68] = t[92] ^ x[26];
  assign t[69] = t[93] ^ x[25];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[94] ^ x[29];
  assign t[71] = t[95] ^ x[28];
  assign t[72] = t[96] ^ x[32];
  assign t[73] = t[97] ^ x[31];
  assign t[74] = t[98] ^ x[35];
  assign t[75] = t[99] ^ x[34];
  assign t[76] = (x[0]);
  assign t[77] = (x[0]);
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind34(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[18] | t[13]);
  assign t[12] = ~(t[24]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[25] | t[26]);
  assign t[15] = ~(t[16] | t[27]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[17] & ~t[18]);
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[17];
  assign t[34] = t[46] ^ x[20];
  assign t[35] = t[47] ^ x[23];
  assign t[36] = t[48] ^ x[26];
  assign t[37] = t[49] ^ x[29];
  assign t[38] = t[50] ^ x[32];
  assign t[39] = t[51] ^ x[35];
  assign t[3] = t[17] & t[4];
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[61]);
  assign t[45] = (t[62] & ~t[63]);
  assign t[46] = (t[64] & ~t[65]);
  assign t[47] = (t[66] & ~t[67]);
  assign t[48] = (t[68] & ~t[69]);
  assign t[49] = (t[70] & ~t[71]);
  assign t[4] = t[5] & t[6];
  assign t[50] = (t[72] & ~t[73]);
  assign t[51] = (t[74] & ~t[75]);
  assign t[52] = t[76] ^ x[2];
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[5];
  assign t[55] = t[79] ^ x[4];
  assign t[56] = t[80] ^ x[8];
  assign t[57] = t[81] ^ x[7];
  assign t[58] = t[82] ^ x[11];
  assign t[59] = t[83] ^ x[10];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[84] ^ x[14];
  assign t[61] = t[85] ^ x[13];
  assign t[62] = t[86] ^ x[17];
  assign t[63] = t[87] ^ x[16];
  assign t[64] = t[88] ^ x[20];
  assign t[65] = t[89] ^ x[19];
  assign t[66] = t[90] ^ x[23];
  assign t[67] = t[91] ^ x[22];
  assign t[68] = t[92] ^ x[26];
  assign t[69] = t[93] ^ x[25];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[94] ^ x[29];
  assign t[71] = t[95] ^ x[28];
  assign t[72] = t[96] ^ x[32];
  assign t[73] = t[97] ^ x[31];
  assign t[74] = t[98] ^ x[35];
  assign t[75] = t[99] ^ x[34];
  assign t[76] = (x[0]);
  assign t[77] = (x[0]);
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[18] | t[13]);
  assign t[12] = ~(t[24]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[25] | t[26]);
  assign t[15] = ~(t[16] | t[27]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[17] & ~t[18]);
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[17];
  assign t[34] = t[46] ^ x[20];
  assign t[35] = t[47] ^ x[23];
  assign t[36] = t[48] ^ x[26];
  assign t[37] = t[49] ^ x[29];
  assign t[38] = t[50] ^ x[32];
  assign t[39] = t[51] ^ x[35];
  assign t[3] = t[17] & t[4];
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[61]);
  assign t[45] = (t[62] & ~t[63]);
  assign t[46] = (t[64] & ~t[65]);
  assign t[47] = (t[66] & ~t[67]);
  assign t[48] = (t[68] & ~t[69]);
  assign t[49] = (t[70] & ~t[71]);
  assign t[4] = t[5] & t[6];
  assign t[50] = (t[72] & ~t[73]);
  assign t[51] = (t[74] & ~t[75]);
  assign t[52] = t[76] ^ x[2];
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[5];
  assign t[55] = t[79] ^ x[4];
  assign t[56] = t[80] ^ x[8];
  assign t[57] = t[81] ^ x[7];
  assign t[58] = t[82] ^ x[11];
  assign t[59] = t[83] ^ x[10];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[84] ^ x[14];
  assign t[61] = t[85] ^ x[13];
  assign t[62] = t[86] ^ x[17];
  assign t[63] = t[87] ^ x[16];
  assign t[64] = t[88] ^ x[20];
  assign t[65] = t[89] ^ x[19];
  assign t[66] = t[90] ^ x[23];
  assign t[67] = t[91] ^ x[22];
  assign t[68] = t[92] ^ x[26];
  assign t[69] = t[93] ^ x[25];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[94] ^ x[29];
  assign t[71] = t[95] ^ x[28];
  assign t[72] = t[96] ^ x[32];
  assign t[73] = t[97] ^ x[31];
  assign t[74] = t[98] ^ x[35];
  assign t[75] = t[99] ^ x[34];
  assign t[76] = (x[0]);
  assign t[77] = (x[0]);
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind36(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[24] | t[13]);
  assign t[12] = ~(t[25]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[26] | t[16]);
  assign t[15] = ~(t[18] | t[27]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = t[17] & t[18];
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[17];
  assign t[34] = t[46] ^ x[20];
  assign t[35] = t[47] ^ x[23];
  assign t[36] = t[48] ^ x[26];
  assign t[37] = t[49] ^ x[29];
  assign t[38] = t[50] ^ x[32];
  assign t[39] = t[51] ^ x[35];
  assign t[3] = t[17] & t[4];
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[61]);
  assign t[45] = (t[62] & ~t[63]);
  assign t[46] = (t[64] & ~t[65]);
  assign t[47] = (t[66] & ~t[67]);
  assign t[48] = (t[68] & ~t[69]);
  assign t[49] = (t[70] & ~t[71]);
  assign t[4] = t[5] & t[6];
  assign t[50] = (t[72] & ~t[73]);
  assign t[51] = (t[74] & ~t[75]);
  assign t[52] = t[76] ^ x[2];
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[5];
  assign t[55] = t[79] ^ x[4];
  assign t[56] = t[80] ^ x[8];
  assign t[57] = t[81] ^ x[7];
  assign t[58] = t[82] ^ x[11];
  assign t[59] = t[83] ^ x[10];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[84] ^ x[14];
  assign t[61] = t[85] ^ x[13];
  assign t[62] = t[86] ^ x[17];
  assign t[63] = t[87] ^ x[16];
  assign t[64] = t[88] ^ x[20];
  assign t[65] = t[89] ^ x[19];
  assign t[66] = t[90] ^ x[23];
  assign t[67] = t[91] ^ x[22];
  assign t[68] = t[92] ^ x[26];
  assign t[69] = t[93] ^ x[25];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[94] ^ x[29];
  assign t[71] = t[95] ^ x[28];
  assign t[72] = t[96] ^ x[32];
  assign t[73] = t[97] ^ x[31];
  assign t[74] = t[98] ^ x[35];
  assign t[75] = t[99] ^ x[34];
  assign t[76] = (x[0]);
  assign t[77] = (x[0]);
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind37(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[24] | t[13]);
  assign t[12] = ~(t[25]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[26] | t[16]);
  assign t[15] = ~(t[18] | t[27]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = t[17] & t[18];
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[17];
  assign t[34] = t[46] ^ x[20];
  assign t[35] = t[47] ^ x[23];
  assign t[36] = t[48] ^ x[26];
  assign t[37] = t[49] ^ x[29];
  assign t[38] = t[50] ^ x[32];
  assign t[39] = t[51] ^ x[35];
  assign t[3] = t[17] & t[4];
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[61]);
  assign t[45] = (t[62] & ~t[63]);
  assign t[46] = (t[64] & ~t[65]);
  assign t[47] = (t[66] & ~t[67]);
  assign t[48] = (t[68] & ~t[69]);
  assign t[49] = (t[70] & ~t[71]);
  assign t[4] = t[5] & t[6];
  assign t[50] = (t[72] & ~t[73]);
  assign t[51] = (t[74] & ~t[75]);
  assign t[52] = t[76] ^ x[2];
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[5];
  assign t[55] = t[79] ^ x[4];
  assign t[56] = t[80] ^ x[8];
  assign t[57] = t[81] ^ x[7];
  assign t[58] = t[82] ^ x[11];
  assign t[59] = t[83] ^ x[10];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[84] ^ x[14];
  assign t[61] = t[85] ^ x[13];
  assign t[62] = t[86] ^ x[17];
  assign t[63] = t[87] ^ x[16];
  assign t[64] = t[88] ^ x[20];
  assign t[65] = t[89] ^ x[19];
  assign t[66] = t[90] ^ x[23];
  assign t[67] = t[91] ^ x[22];
  assign t[68] = t[92] ^ x[26];
  assign t[69] = t[93] ^ x[25];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[94] ^ x[29];
  assign t[71] = t[95] ^ x[28];
  assign t[72] = t[96] ^ x[32];
  assign t[73] = t[97] ^ x[31];
  assign t[74] = t[98] ^ x[35];
  assign t[75] = t[99] ^ x[34];
  assign t[76] = (x[0]);
  assign t[77] = (x[0]);
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind38(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[24] | t[13]);
  assign t[12] = ~(t[25]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[26] | t[18]);
  assign t[15] = ~(t[27] | t[16]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[17] & ~t[18]);
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[17];
  assign t[34] = t[46] ^ x[20];
  assign t[35] = t[47] ^ x[23];
  assign t[36] = t[48] ^ x[26];
  assign t[37] = t[49] ^ x[29];
  assign t[38] = t[50] ^ x[32];
  assign t[39] = t[51] ^ x[35];
  assign t[3] = t[17] & t[4];
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[61]);
  assign t[45] = (t[62] & ~t[63]);
  assign t[46] = (t[64] & ~t[65]);
  assign t[47] = (t[66] & ~t[67]);
  assign t[48] = (t[68] & ~t[69]);
  assign t[49] = (t[70] & ~t[71]);
  assign t[4] = t[5] & t[6];
  assign t[50] = (t[72] & ~t[73]);
  assign t[51] = (t[74] & ~t[75]);
  assign t[52] = t[76] ^ x[2];
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[5];
  assign t[55] = t[79] ^ x[4];
  assign t[56] = t[80] ^ x[8];
  assign t[57] = t[81] ^ x[7];
  assign t[58] = t[82] ^ x[11];
  assign t[59] = t[83] ^ x[10];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[84] ^ x[14];
  assign t[61] = t[85] ^ x[13];
  assign t[62] = t[86] ^ x[17];
  assign t[63] = t[87] ^ x[16];
  assign t[64] = t[88] ^ x[20];
  assign t[65] = t[89] ^ x[19];
  assign t[66] = t[90] ^ x[23];
  assign t[67] = t[91] ^ x[22];
  assign t[68] = t[92] ^ x[26];
  assign t[69] = t[93] ^ x[25];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[94] ^ x[29];
  assign t[71] = t[95] ^ x[28];
  assign t[72] = t[96] ^ x[32];
  assign t[73] = t[97] ^ x[31];
  assign t[74] = t[98] ^ x[35];
  assign t[75] = t[99] ^ x[34];
  assign t[76] = (x[0]);
  assign t[77] = (x[0]);
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind39(x, y);
 input [35:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[23] & t[12]);
  assign t[11] = ~(t[24] | t[13]);
  assign t[12] = ~(t[25]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[26] | t[18]);
  assign t[15] = ~(t[27] | t[16]);
  assign t[16] = (t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[5];
  assign t[2] = ~(t[17] & ~t[18]);
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[11];
  assign t[32] = t[44] ^ x[14];
  assign t[33] = t[45] ^ x[17];
  assign t[34] = t[46] ^ x[20];
  assign t[35] = t[47] ^ x[23];
  assign t[36] = t[48] ^ x[26];
  assign t[37] = t[49] ^ x[29];
  assign t[38] = t[50] ^ x[32];
  assign t[39] = t[51] ^ x[35];
  assign t[3] = t[17] & t[4];
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = (t[60] & ~t[61]);
  assign t[45] = (t[62] & ~t[63]);
  assign t[46] = (t[64] & ~t[65]);
  assign t[47] = (t[66] & ~t[67]);
  assign t[48] = (t[68] & ~t[69]);
  assign t[49] = (t[70] & ~t[71]);
  assign t[4] = t[5] & t[6];
  assign t[50] = (t[72] & ~t[73]);
  assign t[51] = (t[74] & ~t[75]);
  assign t[52] = t[76] ^ x[2];
  assign t[53] = t[77] ^ x[1];
  assign t[54] = t[78] ^ x[5];
  assign t[55] = t[79] ^ x[4];
  assign t[56] = t[80] ^ x[8];
  assign t[57] = t[81] ^ x[7];
  assign t[58] = t[82] ^ x[11];
  assign t[59] = t[83] ^ x[10];
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = t[84] ^ x[14];
  assign t[61] = t[85] ^ x[13];
  assign t[62] = t[86] ^ x[17];
  assign t[63] = t[87] ^ x[16];
  assign t[64] = t[88] ^ x[20];
  assign t[65] = t[89] ^ x[19];
  assign t[66] = t[90] ^ x[23];
  assign t[67] = t[91] ^ x[22];
  assign t[68] = t[92] ^ x[26];
  assign t[69] = t[93] ^ x[25];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[94] ^ x[29];
  assign t[71] = t[95] ^ x[28];
  assign t[72] = t[96] ^ x[32];
  assign t[73] = t[97] ^ x[31];
  assign t[74] = t[98] ^ x[35];
  assign t[75] = t[99] ^ x[34];
  assign t[76] = (x[0]);
  assign t[77] = (x[0]);
  assign t[78] = (x[3]);
  assign t[79] = (x[3]);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[6]);
  assign t[81] = (x[6]);
  assign t[82] = (x[9]);
  assign t[83] = (x[9]);
  assign t[84] = (x[12]);
  assign t[85] = (x[12]);
  assign t[86] = (x[15]);
  assign t[87] = (x[15]);
  assign t[88] = (x[18]);
  assign t[89] = (x[18]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[21]);
  assign t[91] = (x[21]);
  assign t[92] = (x[24]);
  assign t[93] = (x[24]);
  assign t[94] = (x[27]);
  assign t[95] = (x[27]);
  assign t[96] = (x[30]);
  assign t[97] = (x[30]);
  assign t[98] = (x[33]);
  assign t[99] = (x[33]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind41(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind46(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind51(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [60:0] x;
 output y;

 wire [181:0] t;
  assign t[0] = t[1] ? t[2] : t[42];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = t[142] ^ x[2];
  assign t[103] = t[143] ^ x[1];
  assign t[104] = t[144] ^ x[5];
  assign t[105] = t[145] ^ x[4];
  assign t[106] = t[146] ^ x[9];
  assign t[107] = t[147] ^ x[8];
  assign t[108] = t[148] ^ x[12];
  assign t[109] = t[149] ^ x[11];
  assign t[10] = ~(t[16]);
  assign t[110] = t[150] ^ x[15];
  assign t[111] = t[151] ^ x[14];
  assign t[112] = t[152] ^ x[18];
  assign t[113] = t[153] ^ x[17];
  assign t[114] = t[154] ^ x[21];
  assign t[115] = t[155] ^ x[20];
  assign t[116] = t[156] ^ x[24];
  assign t[117] = t[157] ^ x[23];
  assign t[118] = t[158] ^ x[27];
  assign t[119] = t[159] ^ x[26];
  assign t[11] = t[45] & t[17];
  assign t[120] = t[160] ^ x[30];
  assign t[121] = t[161] ^ x[29];
  assign t[122] = t[162] ^ x[33];
  assign t[123] = t[163] ^ x[32];
  assign t[124] = t[164] ^ x[36];
  assign t[125] = t[165] ^ x[35];
  assign t[126] = t[166] ^ x[39];
  assign t[127] = t[167] ^ x[38];
  assign t[128] = t[168] ^ x[42];
  assign t[129] = t[169] ^ x[41];
  assign t[12] = ~(t[18] | t[19]);
  assign t[130] = t[170] ^ x[45];
  assign t[131] = t[171] ^ x[44];
  assign t[132] = t[172] ^ x[48];
  assign t[133] = t[173] ^ x[47];
  assign t[134] = t[174] ^ x[51];
  assign t[135] = t[175] ^ x[50];
  assign t[136] = t[176] ^ x[54];
  assign t[137] = t[177] ^ x[53];
  assign t[138] = t[178] ^ x[57];
  assign t[139] = t[179] ^ x[56];
  assign t[13] = ~(t[45]);
  assign t[140] = t[180] ^ x[60];
  assign t[141] = t[181] ^ x[59];
  assign t[142] = (x[0]);
  assign t[143] = (x[0]);
  assign t[144] = (x[3]);
  assign t[145] = (x[3]);
  assign t[146] = (x[7]);
  assign t[147] = (x[7]);
  assign t[148] = (x[10]);
  assign t[149] = (x[10]);
  assign t[14] = t[20] & t[21];
  assign t[150] = (x[13]);
  assign t[151] = (x[13]);
  assign t[152] = (x[16]);
  assign t[153] = (x[16]);
  assign t[154] = (x[19]);
  assign t[155] = (x[19]);
  assign t[156] = (x[22]);
  assign t[157] = (x[22]);
  assign t[158] = (x[25]);
  assign t[159] = (x[25]);
  assign t[15] = t[44] ^ t[42];
  assign t[160] = (x[28]);
  assign t[161] = (x[28]);
  assign t[162] = (x[31]);
  assign t[163] = (x[31]);
  assign t[164] = (x[34]);
  assign t[165] = (x[34]);
  assign t[166] = (x[37]);
  assign t[167] = (x[37]);
  assign t[168] = (x[40]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[45] & t[22]);
  assign t[170] = (x[43]);
  assign t[171] = (x[43]);
  assign t[172] = (x[46]);
  assign t[173] = (x[46]);
  assign t[174] = (x[49]);
  assign t[175] = (x[49]);
  assign t[176] = (x[52]);
  assign t[177] = (x[52]);
  assign t[178] = (x[55]);
  assign t[179] = (x[55]);
  assign t[17] = t[23] & t[24];
  assign t[180] = (x[58]);
  assign t[181] = (x[58]);
  assign t[18] = ~(t[46]);
  assign t[19] = ~(t[45]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[19] | t[27]);
  assign t[22] = ~(t[47] | t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[25] = ~(t[48] | t[49]);
  assign t[26] = ~(t[33] | t[34]);
  assign t[27] = ~(t[50] | t[51]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[52] & t[49]);
  assign t[2] = t[4] ? t[43] : t[5];
  assign t[30] = ~(t[48] & t[53]);
  assign t[31] = ~(t[22]);
  assign t[32] = ~(t[51] & t[37]);
  assign t[33] = ~(t[53] & t[54]);
  assign t[34] = ~(t[38] & t[39]);
  assign t[35] = ~(t[55] | t[56]);
  assign t[36] = ~(t[57] | t[58]);
  assign t[37] = ~(t[50]);
  assign t[38] = ~(t[59] | t[40]);
  assign t[39] = ~(t[52] | t[41]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[60]);
  assign t[41] = ~(t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = (t[78]);
  assign t[59] = (t[79]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[80]);
  assign t[61] = (t[81]);
  assign t[62] = t[82] ^ x[2];
  assign t[63] = t[83] ^ x[5];
  assign t[64] = t[84] ^ x[9];
  assign t[65] = t[85] ^ x[12];
  assign t[66] = t[86] ^ x[15];
  assign t[67] = t[87] ^ x[18];
  assign t[68] = t[88] ^ x[21];
  assign t[69] = t[89] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[90] ^ x[27];
  assign t[71] = t[91] ^ x[30];
  assign t[72] = t[92] ^ x[33];
  assign t[73] = t[93] ^ x[36];
  assign t[74] = t[94] ^ x[39];
  assign t[75] = t[95] ^ x[42];
  assign t[76] = t[96] ^ x[45];
  assign t[77] = t[97] ^ x[48];
  assign t[78] = t[98] ^ x[51];
  assign t[79] = t[99] ^ x[54];
  assign t[7] = ~(t[12]);
  assign t[80] = t[100] ^ x[57];
  assign t[81] = t[101] ^ x[60];
  assign t[82] = (t[102] & ~t[103]);
  assign t[83] = (t[104] & ~t[105]);
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[13]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[14] ? t[15] : t[44];
  assign y = (t[0]);
endmodule

module R2ind56(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind61(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind66(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind71(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind76(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind81(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind86(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind91(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind96(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind101(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind106(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind111(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind116(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind121(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind126(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind131(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind136(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind141(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind146(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind151(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind156(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind161(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind166(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind171(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind176(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind181(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind186(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind191(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind196(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind201(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind206(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind211(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind216(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind221(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind226(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind231(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [123:0] x;
 output y;

 wire [422:0] t;
  assign t[0] = t[1] ? t[2] : t[136];
  assign t[100] = t[170] ^ t[171];
  assign t[101] = t[172] ^ t[173];
  assign t[102] = t[13] ? t[174] : t[111];
  assign t[103] = t[112] ^ t[113];
  assign t[104] = t[54] ^ t[114];
  assign t[105] = t[115] ^ t[116];
  assign t[106] = t[117] ^ t[118];
  assign t[107] = t[119] ^ t[120];
  assign t[108] = t[119] & t[120];
  assign t[109] = t[54] & t[121];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[122] ^ t[116];
  assign t[111] = t[175] ^ t[176];
  assign t[112] = t[104] & t[71];
  assign t[113] = t[55] & t[53];
  assign t[114] = t[87] ^ t[123];
  assign t[115] = t[124] ^ t[125];
  assign t[116] = t[126] ^ t[109];
  assign t[117] = t[114] & t[61];
  assign t[118] = t[127] & t[59];
  assign t[119] = t[69] ^ t[51];
  assign t[11] = ~(t[17]);
  assign t[120] = t[59] ^ t[87];
  assign t[121] = t[67] ^ t[128];
  assign t[122] = t[129] ^ t[130];
  assign t[123] = t[50] ^ t[61];
  assign t[124] = t[131] ^ t[113];
  assign t[125] = t[72] & t[86];
  assign t[126] = t[38] & t[132];
  assign t[127] = t[55] ^ t[38];
  assign t[128] = t[102] ^ t[51];
  assign t[129] = t[133] ^ t[118];
  assign t[12] = t[139] & t[18];
  assign t[130] = t[134] & t[135];
  assign t[131] = t[55] ^ t[53];
  assign t[132] = t[54] ^ t[68];
  assign t[133] = t[59] ^ t[128];
  assign t[134] = t[119] ^ t[72];
  assign t[135] = t[61] ^ t[59];
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = ~(t[139]);
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = (t[194]);
  assign t[154] = (t[195]);
  assign t[155] = (t[196]);
  assign t[156] = (t[197]);
  assign t[157] = (t[198]);
  assign t[158] = (t[199]);
  assign t[159] = (t[200]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[201]);
  assign t[161] = (t[202]);
  assign t[162] = (t[203]);
  assign t[163] = (t[204]);
  assign t[164] = (t[205]);
  assign t[165] = (t[206]);
  assign t[166] = (t[207]);
  assign t[167] = (t[208]);
  assign t[168] = (t[209]);
  assign t[169] = (t[210]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (t[211]);
  assign t[171] = (t[212]);
  assign t[172] = (t[213]);
  assign t[173] = (t[214]);
  assign t[174] = (t[215]);
  assign t[175] = (t[216]);
  assign t[176] = (t[217]);
  assign t[177] = t[218] ^ x[2];
  assign t[178] = t[219] ^ x[6];
  assign t[179] = t[220] ^ x[9];
  assign t[17] = ~(t[139] & t[25]);
  assign t[180] = t[221] ^ x[12];
  assign t[181] = t[222] ^ x[15];
  assign t[182] = t[223] ^ x[18];
  assign t[183] = t[224] ^ x[21];
  assign t[184] = t[225] ^ x[24];
  assign t[185] = t[226] ^ x[27];
  assign t[186] = t[227] ^ x[30];
  assign t[187] = t[228] ^ x[33];
  assign t[188] = t[229] ^ x[36];
  assign t[189] = t[230] ^ x[39];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[231] ^ x[42];
  assign t[191] = t[232] ^ x[45];
  assign t[192] = t[233] ^ x[48];
  assign t[193] = t[234] ^ x[51];
  assign t[194] = t[235] ^ x[54];
  assign t[195] = t[236] ^ x[57];
  assign t[196] = t[237] ^ x[60];
  assign t[197] = t[238] ^ x[63];
  assign t[198] = t[239] ^ x[66];
  assign t[199] = t[240] ^ x[69];
  assign t[19] = ~(t[140]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[241] ^ x[72];
  assign t[201] = t[242] ^ x[75];
  assign t[202] = t[243] ^ x[78];
  assign t[203] = t[244] ^ x[81];
  assign t[204] = t[245] ^ x[84];
  assign t[205] = t[246] ^ x[87];
  assign t[206] = t[247] ^ x[90];
  assign t[207] = t[248] ^ x[93];
  assign t[208] = t[249] ^ x[96];
  assign t[209] = t[250] ^ x[99];
  assign t[20] = ~(t[139]);
  assign t[210] = t[251] ^ x[102];
  assign t[211] = t[252] ^ x[105];
  assign t[212] = t[253] ^ x[108];
  assign t[213] = t[254] ^ x[111];
  assign t[214] = t[255] ^ x[114];
  assign t[215] = t[256] ^ x[117];
  assign t[216] = t[257] ^ x[120];
  assign t[217] = t[258] ^ x[123];
  assign t[218] = (t[259] & ~t[260]);
  assign t[219] = (t[261] & ~t[262]);
  assign t[21] = ~(t[141]);
  assign t[220] = (t[263] & ~t[264]);
  assign t[221] = (t[265] & ~t[266]);
  assign t[222] = (t[267] & ~t[268]);
  assign t[223] = (t[269] & ~t[270]);
  assign t[224] = (t[271] & ~t[272]);
  assign t[225] = (t[273] & ~t[274]);
  assign t[226] = (t[275] & ~t[276]);
  assign t[227] = (t[277] & ~t[278]);
  assign t[228] = (t[279] & ~t[280]);
  assign t[229] = (t[281] & ~t[282]);
  assign t[22] = ~(t[142]);
  assign t[230] = (t[283] & ~t[284]);
  assign t[231] = (t[285] & ~t[286]);
  assign t[232] = (t[287] & ~t[288]);
  assign t[233] = (t[289] & ~t[290]);
  assign t[234] = (t[291] & ~t[292]);
  assign t[235] = (t[293] & ~t[294]);
  assign t[236] = (t[295] & ~t[296]);
  assign t[237] = (t[297] & ~t[298]);
  assign t[238] = (t[299] & ~t[300]);
  assign t[239] = (t[301] & ~t[302]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[303] & ~t[304]);
  assign t[241] = (t[305] & ~t[306]);
  assign t[242] = (t[307] & ~t[308]);
  assign t[243] = (t[309] & ~t[310]);
  assign t[244] = (t[311] & ~t[312]);
  assign t[245] = (t[313] & ~t[314]);
  assign t[246] = (t[315] & ~t[316]);
  assign t[247] = (t[317] & ~t[318]);
  assign t[248] = (t[319] & ~t[320]);
  assign t[249] = (t[321] & ~t[322]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[323] & ~t[324]);
  assign t[251] = (t[325] & ~t[326]);
  assign t[252] = (t[327] & ~t[328]);
  assign t[253] = (t[329] & ~t[330]);
  assign t[254] = (t[331] & ~t[332]);
  assign t[255] = (t[333] & ~t[334]);
  assign t[256] = (t[335] & ~t[336]);
  assign t[257] = (t[337] & ~t[338]);
  assign t[258] = (t[339] & ~t[340]);
  assign t[259] = t[341] ^ x[2];
  assign t[25] = ~(t[143] | t[32]);
  assign t[260] = t[342] ^ x[1];
  assign t[261] = t[343] ^ x[6];
  assign t[262] = t[344] ^ x[5];
  assign t[263] = t[345] ^ x[9];
  assign t[264] = t[346] ^ x[8];
  assign t[265] = t[347] ^ x[12];
  assign t[266] = t[348] ^ x[11];
  assign t[267] = t[349] ^ x[15];
  assign t[268] = t[350] ^ x[14];
  assign t[269] = t[351] ^ x[18];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[352] ^ x[17];
  assign t[271] = t[353] ^ x[21];
  assign t[272] = t[354] ^ x[20];
  assign t[273] = t[355] ^ x[24];
  assign t[274] = t[356] ^ x[23];
  assign t[275] = t[357] ^ x[27];
  assign t[276] = t[358] ^ x[26];
  assign t[277] = t[359] ^ x[30];
  assign t[278] = t[360] ^ x[29];
  assign t[279] = t[361] ^ x[33];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[362] ^ x[32];
  assign t[281] = t[363] ^ x[36];
  assign t[282] = t[364] ^ x[35];
  assign t[283] = t[365] ^ x[39];
  assign t[284] = t[366] ^ x[38];
  assign t[285] = t[367] ^ x[42];
  assign t[286] = t[368] ^ x[41];
  assign t[287] = t[369] ^ x[45];
  assign t[288] = t[370] ^ x[44];
  assign t[289] = t[371] ^ x[48];
  assign t[28] = t[37] & t[38];
  assign t[290] = t[372] ^ x[47];
  assign t[291] = t[373] ^ x[51];
  assign t[292] = t[374] ^ x[50];
  assign t[293] = t[375] ^ x[54];
  assign t[294] = t[376] ^ x[53];
  assign t[295] = t[377] ^ x[57];
  assign t[296] = t[378] ^ x[56];
  assign t[297] = t[379] ^ x[60];
  assign t[298] = t[380] ^ x[59];
  assign t[299] = t[381] ^ x[63];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[62];
  assign t[301] = t[383] ^ x[66];
  assign t[302] = t[384] ^ x[65];
  assign t[303] = t[385] ^ x[69];
  assign t[304] = t[386] ^ x[68];
  assign t[305] = t[387] ^ x[72];
  assign t[306] = t[388] ^ x[71];
  assign t[307] = t[389] ^ x[75];
  assign t[308] = t[390] ^ x[74];
  assign t[309] = t[391] ^ x[78];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[392] ^ x[77];
  assign t[311] = t[393] ^ x[81];
  assign t[312] = t[394] ^ x[80];
  assign t[313] = t[395] ^ x[84];
  assign t[314] = t[396] ^ x[83];
  assign t[315] = t[397] ^ x[87];
  assign t[316] = t[398] ^ x[86];
  assign t[317] = t[399] ^ x[90];
  assign t[318] = t[400] ^ x[89];
  assign t[319] = t[401] ^ x[93];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[402] ^ x[92];
  assign t[321] = t[403] ^ x[96];
  assign t[322] = t[404] ^ x[95];
  assign t[323] = t[405] ^ x[99];
  assign t[324] = t[406] ^ x[98];
  assign t[325] = t[407] ^ x[102];
  assign t[326] = t[408] ^ x[101];
  assign t[327] = t[409] ^ x[105];
  assign t[328] = t[410] ^ x[104];
  assign t[329] = t[411] ^ x[108];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[412] ^ x[107];
  assign t[331] = t[413] ^ x[111];
  assign t[332] = t[414] ^ x[110];
  assign t[333] = t[415] ^ x[114];
  assign t[334] = t[416] ^ x[113];
  assign t[335] = t[417] ^ x[117];
  assign t[336] = t[418] ^ x[116];
  assign t[337] = t[419] ^ x[120];
  assign t[338] = t[420] ^ x[119];
  assign t[339] = t[421] ^ x[123];
  assign t[33] = ~(t[144] & t[145]);
  assign t[340] = t[422] ^ x[122];
  assign t[341] = (x[0]);
  assign t[342] = (x[0]);
  assign t[343] = (x[4]);
  assign t[344] = (x[4]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[146] & t[147]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[148] & t[47]);
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[49]);
  assign t[374] = (x[49]);
  assign t[375] = (x[52]);
  assign t[376] = (x[52]);
  assign t[377] = (x[55]);
  assign t[378] = (x[55]);
  assign t[379] = (x[58]);
  assign t[37] = t[48] ^ t[49];
  assign t[380] = (x[58]);
  assign t[381] = (x[61]);
  assign t[382] = (x[61]);
  assign t[383] = (x[64]);
  assign t[384] = (x[64]);
  assign t[385] = (x[67]);
  assign t[386] = (x[67]);
  assign t[387] = (x[70]);
  assign t[388] = (x[70]);
  assign t[389] = (x[73]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[73]);
  assign t[391] = (x[76]);
  assign t[392] = (x[76]);
  assign t[393] = (x[79]);
  assign t[394] = (x[79]);
  assign t[395] = (x[82]);
  assign t[396] = (x[82]);
  assign t[397] = (x[85]);
  assign t[398] = (x[85]);
  assign t[399] = (x[88]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[88]);
  assign t[401] = (x[91]);
  assign t[402] = (x[91]);
  assign t[403] = (x[94]);
  assign t[404] = (x[94]);
  assign t[405] = (x[97]);
  assign t[406] = (x[97]);
  assign t[407] = (x[100]);
  assign t[408] = (x[100]);
  assign t[409] = (x[103]);
  assign t[40] = t[48] & t[54];
  assign t[410] = (x[103]);
  assign t[411] = (x[106]);
  assign t[412] = (x[106]);
  assign t[413] = (x[109]);
  assign t[414] = (x[109]);
  assign t[415] = (x[112]);
  assign t[416] = (x[112]);
  assign t[417] = (x[115]);
  assign t[418] = (x[115]);
  assign t[419] = (x[118]);
  assign t[41] = t[52] & t[55];
  assign t[420] = (x[118]);
  assign t[421] = (x[121]);
  assign t[422] = (x[121]);
  assign t[42] = t[56] ^ t[57];
  assign t[43] = t[58] & t[59];
  assign t[44] = t[60] & t[61];
  assign t[45] = ~(t[149] | t[150]);
  assign t[46] = ~(t[151] | t[152]);
  assign t[47] = ~(t[153]);
  assign t[48] = t[62] ^ t[60];
  assign t[49] = t[63] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[13] ? t[154] : t[65];
  assign t[51] = t[13] ? t[155] : t[66];
  assign t[52] = t[62] ^ t[63];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[69] ^ t[50];
  assign t[55] = t[69] ^ t[70];
  assign t[56] = t[62] & t[71];
  assign t[57] = t[63] & t[72];
  assign t[58] = t[60] ^ t[64];
  assign t[59] = t[54] ^ t[67];
  assign t[5] = t[9] ? t[137] : x[3];
  assign t[60] = t[73] ^ t[74];
  assign t[61] = t[13] ? t[156] : t[75];
  assign t[62] = t[76] ^ t[77];
  assign t[63] = t[78] ^ t[79];
  assign t[64] = t[80] ^ t[81];
  assign t[65] = t[157] ^ t[158];
  assign t[66] = t[159] ^ t[160];
  assign t[67] = t[82] ^ t[70];
  assign t[68] = t[83] ^ t[51];
  assign t[69] = t[13] ? t[161] : t[84];
  assign t[6] = ~(t[10] ^ t[138]);
  assign t[70] = t[13] ? t[162] : t[85];
  assign t[71] = t[86] ^ t[53];
  assign t[72] = t[87] ^ t[88];
  assign t[73] = t[89] ^ t[90];
  assign t[74] = t[91] & t[92];
  assign t[75] = t[163] ^ t[138];
  assign t[76] = t[93] ^ t[94];
  assign t[77] = t[95] & t[96];
  assign t[78] = t[96] & t[97];
  assign t[79] = t[96] ^ t[98];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[92] & t[99];
  assign t[81] = t[92] ^ t[98];
  assign t[82] = t[13] ? t[164] : t[100];
  assign t[83] = t[13] ? t[165] : t[101];
  assign t[84] = t[166] ^ t[167];
  assign t[85] = t[168] ^ t[169];
  assign t[86] = t[61] ^ t[87];
  assign t[87] = t[102] ^ t[83];
  assign t[88] = t[70] ^ t[61];
  assign t[89] = t[103] ^ t[94];
  assign t[8] = ~(t[13]);
  assign t[90] = t[104] ^ t[71];
  assign t[91] = t[76] ^ t[98];
  assign t[92] = t[105] ^ t[73];
  assign t[93] = t[106] ^ t[107];
  assign t[94] = t[108] ^ t[109];
  assign t[95] = t[73] ^ t[98];
  assign t[96] = t[110] ^ t[76];
  assign t[97] = t[110] & t[73];
  assign t[98] = t[105] & t[110];
  assign t[99] = t[76] & t[105];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [123:0] x;
 output y;

 wire [422:0] t;
  assign t[0] = t[1] ? t[2] : t[136];
  assign t[100] = t[170] ^ t[171];
  assign t[101] = t[172] ^ t[173];
  assign t[102] = t[13] ? t[174] : t[111];
  assign t[103] = t[112] ^ t[113];
  assign t[104] = t[54] ^ t[114];
  assign t[105] = t[115] ^ t[116];
  assign t[106] = t[117] ^ t[118];
  assign t[107] = t[119] ^ t[120];
  assign t[108] = t[119] & t[120];
  assign t[109] = t[54] & t[121];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[122] ^ t[116];
  assign t[111] = t[175] ^ t[176];
  assign t[112] = t[104] & t[71];
  assign t[113] = t[55] & t[53];
  assign t[114] = t[87] ^ t[123];
  assign t[115] = t[124] ^ t[125];
  assign t[116] = t[126] ^ t[109];
  assign t[117] = t[114] & t[61];
  assign t[118] = t[127] & t[59];
  assign t[119] = t[69] ^ t[51];
  assign t[11] = ~(t[17]);
  assign t[120] = t[59] ^ t[87];
  assign t[121] = t[67] ^ t[128];
  assign t[122] = t[129] ^ t[130];
  assign t[123] = t[50] ^ t[61];
  assign t[124] = t[131] ^ t[113];
  assign t[125] = t[72] & t[86];
  assign t[126] = t[38] & t[132];
  assign t[127] = t[55] ^ t[38];
  assign t[128] = t[102] ^ t[51];
  assign t[129] = t[133] ^ t[118];
  assign t[12] = t[139] & t[18];
  assign t[130] = t[134] & t[135];
  assign t[131] = t[55] ^ t[53];
  assign t[132] = t[54] ^ t[68];
  assign t[133] = t[59] ^ t[128];
  assign t[134] = t[119] ^ t[72];
  assign t[135] = t[61] ^ t[59];
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = ~(t[139]);
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = (t[194]);
  assign t[154] = (t[195]);
  assign t[155] = (t[196]);
  assign t[156] = (t[197]);
  assign t[157] = (t[198]);
  assign t[158] = (t[199]);
  assign t[159] = (t[200]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[201]);
  assign t[161] = (t[202]);
  assign t[162] = (t[203]);
  assign t[163] = (t[204]);
  assign t[164] = (t[205]);
  assign t[165] = (t[206]);
  assign t[166] = (t[207]);
  assign t[167] = (t[208]);
  assign t[168] = (t[209]);
  assign t[169] = (t[210]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (t[211]);
  assign t[171] = (t[212]);
  assign t[172] = (t[213]);
  assign t[173] = (t[214]);
  assign t[174] = (t[215]);
  assign t[175] = (t[216]);
  assign t[176] = (t[217]);
  assign t[177] = t[218] ^ x[2];
  assign t[178] = t[219] ^ x[6];
  assign t[179] = t[220] ^ x[9];
  assign t[17] = ~(t[139] & t[25]);
  assign t[180] = t[221] ^ x[12];
  assign t[181] = t[222] ^ x[15];
  assign t[182] = t[223] ^ x[18];
  assign t[183] = t[224] ^ x[21];
  assign t[184] = t[225] ^ x[24];
  assign t[185] = t[226] ^ x[27];
  assign t[186] = t[227] ^ x[30];
  assign t[187] = t[228] ^ x[33];
  assign t[188] = t[229] ^ x[36];
  assign t[189] = t[230] ^ x[39];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[231] ^ x[42];
  assign t[191] = t[232] ^ x[45];
  assign t[192] = t[233] ^ x[48];
  assign t[193] = t[234] ^ x[51];
  assign t[194] = t[235] ^ x[54];
  assign t[195] = t[236] ^ x[57];
  assign t[196] = t[237] ^ x[60];
  assign t[197] = t[238] ^ x[63];
  assign t[198] = t[239] ^ x[66];
  assign t[199] = t[240] ^ x[69];
  assign t[19] = ~(t[140]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[241] ^ x[72];
  assign t[201] = t[242] ^ x[75];
  assign t[202] = t[243] ^ x[78];
  assign t[203] = t[244] ^ x[81];
  assign t[204] = t[245] ^ x[84];
  assign t[205] = t[246] ^ x[87];
  assign t[206] = t[247] ^ x[90];
  assign t[207] = t[248] ^ x[93];
  assign t[208] = t[249] ^ x[96];
  assign t[209] = t[250] ^ x[99];
  assign t[20] = ~(t[139]);
  assign t[210] = t[251] ^ x[102];
  assign t[211] = t[252] ^ x[105];
  assign t[212] = t[253] ^ x[108];
  assign t[213] = t[254] ^ x[111];
  assign t[214] = t[255] ^ x[114];
  assign t[215] = t[256] ^ x[117];
  assign t[216] = t[257] ^ x[120];
  assign t[217] = t[258] ^ x[123];
  assign t[218] = (t[259] & ~t[260]);
  assign t[219] = (t[261] & ~t[262]);
  assign t[21] = ~(t[141]);
  assign t[220] = (t[263] & ~t[264]);
  assign t[221] = (t[265] & ~t[266]);
  assign t[222] = (t[267] & ~t[268]);
  assign t[223] = (t[269] & ~t[270]);
  assign t[224] = (t[271] & ~t[272]);
  assign t[225] = (t[273] & ~t[274]);
  assign t[226] = (t[275] & ~t[276]);
  assign t[227] = (t[277] & ~t[278]);
  assign t[228] = (t[279] & ~t[280]);
  assign t[229] = (t[281] & ~t[282]);
  assign t[22] = ~(t[142]);
  assign t[230] = (t[283] & ~t[284]);
  assign t[231] = (t[285] & ~t[286]);
  assign t[232] = (t[287] & ~t[288]);
  assign t[233] = (t[289] & ~t[290]);
  assign t[234] = (t[291] & ~t[292]);
  assign t[235] = (t[293] & ~t[294]);
  assign t[236] = (t[295] & ~t[296]);
  assign t[237] = (t[297] & ~t[298]);
  assign t[238] = (t[299] & ~t[300]);
  assign t[239] = (t[301] & ~t[302]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[303] & ~t[304]);
  assign t[241] = (t[305] & ~t[306]);
  assign t[242] = (t[307] & ~t[308]);
  assign t[243] = (t[309] & ~t[310]);
  assign t[244] = (t[311] & ~t[312]);
  assign t[245] = (t[313] & ~t[314]);
  assign t[246] = (t[315] & ~t[316]);
  assign t[247] = (t[317] & ~t[318]);
  assign t[248] = (t[319] & ~t[320]);
  assign t[249] = (t[321] & ~t[322]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[323] & ~t[324]);
  assign t[251] = (t[325] & ~t[326]);
  assign t[252] = (t[327] & ~t[328]);
  assign t[253] = (t[329] & ~t[330]);
  assign t[254] = (t[331] & ~t[332]);
  assign t[255] = (t[333] & ~t[334]);
  assign t[256] = (t[335] & ~t[336]);
  assign t[257] = (t[337] & ~t[338]);
  assign t[258] = (t[339] & ~t[340]);
  assign t[259] = t[341] ^ x[2];
  assign t[25] = ~(t[143] | t[32]);
  assign t[260] = t[342] ^ x[1];
  assign t[261] = t[343] ^ x[6];
  assign t[262] = t[344] ^ x[5];
  assign t[263] = t[345] ^ x[9];
  assign t[264] = t[346] ^ x[8];
  assign t[265] = t[347] ^ x[12];
  assign t[266] = t[348] ^ x[11];
  assign t[267] = t[349] ^ x[15];
  assign t[268] = t[350] ^ x[14];
  assign t[269] = t[351] ^ x[18];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[352] ^ x[17];
  assign t[271] = t[353] ^ x[21];
  assign t[272] = t[354] ^ x[20];
  assign t[273] = t[355] ^ x[24];
  assign t[274] = t[356] ^ x[23];
  assign t[275] = t[357] ^ x[27];
  assign t[276] = t[358] ^ x[26];
  assign t[277] = t[359] ^ x[30];
  assign t[278] = t[360] ^ x[29];
  assign t[279] = t[361] ^ x[33];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[362] ^ x[32];
  assign t[281] = t[363] ^ x[36];
  assign t[282] = t[364] ^ x[35];
  assign t[283] = t[365] ^ x[39];
  assign t[284] = t[366] ^ x[38];
  assign t[285] = t[367] ^ x[42];
  assign t[286] = t[368] ^ x[41];
  assign t[287] = t[369] ^ x[45];
  assign t[288] = t[370] ^ x[44];
  assign t[289] = t[371] ^ x[48];
  assign t[28] = t[37] & t[38];
  assign t[290] = t[372] ^ x[47];
  assign t[291] = t[373] ^ x[51];
  assign t[292] = t[374] ^ x[50];
  assign t[293] = t[375] ^ x[54];
  assign t[294] = t[376] ^ x[53];
  assign t[295] = t[377] ^ x[57];
  assign t[296] = t[378] ^ x[56];
  assign t[297] = t[379] ^ x[60];
  assign t[298] = t[380] ^ x[59];
  assign t[299] = t[381] ^ x[63];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[62];
  assign t[301] = t[383] ^ x[66];
  assign t[302] = t[384] ^ x[65];
  assign t[303] = t[385] ^ x[69];
  assign t[304] = t[386] ^ x[68];
  assign t[305] = t[387] ^ x[72];
  assign t[306] = t[388] ^ x[71];
  assign t[307] = t[389] ^ x[75];
  assign t[308] = t[390] ^ x[74];
  assign t[309] = t[391] ^ x[78];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[392] ^ x[77];
  assign t[311] = t[393] ^ x[81];
  assign t[312] = t[394] ^ x[80];
  assign t[313] = t[395] ^ x[84];
  assign t[314] = t[396] ^ x[83];
  assign t[315] = t[397] ^ x[87];
  assign t[316] = t[398] ^ x[86];
  assign t[317] = t[399] ^ x[90];
  assign t[318] = t[400] ^ x[89];
  assign t[319] = t[401] ^ x[93];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[402] ^ x[92];
  assign t[321] = t[403] ^ x[96];
  assign t[322] = t[404] ^ x[95];
  assign t[323] = t[405] ^ x[99];
  assign t[324] = t[406] ^ x[98];
  assign t[325] = t[407] ^ x[102];
  assign t[326] = t[408] ^ x[101];
  assign t[327] = t[409] ^ x[105];
  assign t[328] = t[410] ^ x[104];
  assign t[329] = t[411] ^ x[108];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[412] ^ x[107];
  assign t[331] = t[413] ^ x[111];
  assign t[332] = t[414] ^ x[110];
  assign t[333] = t[415] ^ x[114];
  assign t[334] = t[416] ^ x[113];
  assign t[335] = t[417] ^ x[117];
  assign t[336] = t[418] ^ x[116];
  assign t[337] = t[419] ^ x[120];
  assign t[338] = t[420] ^ x[119];
  assign t[339] = t[421] ^ x[123];
  assign t[33] = ~(t[144] & t[145]);
  assign t[340] = t[422] ^ x[122];
  assign t[341] = (x[0]);
  assign t[342] = (x[0]);
  assign t[343] = (x[4]);
  assign t[344] = (x[4]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[146] & t[147]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[148] & t[47]);
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[49]);
  assign t[374] = (x[49]);
  assign t[375] = (x[52]);
  assign t[376] = (x[52]);
  assign t[377] = (x[55]);
  assign t[378] = (x[55]);
  assign t[379] = (x[58]);
  assign t[37] = t[48] ^ t[49];
  assign t[380] = (x[58]);
  assign t[381] = (x[61]);
  assign t[382] = (x[61]);
  assign t[383] = (x[64]);
  assign t[384] = (x[64]);
  assign t[385] = (x[67]);
  assign t[386] = (x[67]);
  assign t[387] = (x[70]);
  assign t[388] = (x[70]);
  assign t[389] = (x[73]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[73]);
  assign t[391] = (x[76]);
  assign t[392] = (x[76]);
  assign t[393] = (x[79]);
  assign t[394] = (x[79]);
  assign t[395] = (x[82]);
  assign t[396] = (x[82]);
  assign t[397] = (x[85]);
  assign t[398] = (x[85]);
  assign t[399] = (x[88]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[88]);
  assign t[401] = (x[91]);
  assign t[402] = (x[91]);
  assign t[403] = (x[94]);
  assign t[404] = (x[94]);
  assign t[405] = (x[97]);
  assign t[406] = (x[97]);
  assign t[407] = (x[100]);
  assign t[408] = (x[100]);
  assign t[409] = (x[103]);
  assign t[40] = t[48] & t[54];
  assign t[410] = (x[103]);
  assign t[411] = (x[106]);
  assign t[412] = (x[106]);
  assign t[413] = (x[109]);
  assign t[414] = (x[109]);
  assign t[415] = (x[112]);
  assign t[416] = (x[112]);
  assign t[417] = (x[115]);
  assign t[418] = (x[115]);
  assign t[419] = (x[118]);
  assign t[41] = t[52] & t[55];
  assign t[420] = (x[118]);
  assign t[421] = (x[121]);
  assign t[422] = (x[121]);
  assign t[42] = t[56] ^ t[57];
  assign t[43] = t[58] & t[59];
  assign t[44] = t[60] & t[61];
  assign t[45] = ~(t[149] | t[150]);
  assign t[46] = ~(t[151] | t[152]);
  assign t[47] = ~(t[153]);
  assign t[48] = t[62] ^ t[60];
  assign t[49] = t[63] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[13] ? t[154] : t[65];
  assign t[51] = t[13] ? t[155] : t[66];
  assign t[52] = t[62] ^ t[63];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[69] ^ t[50];
  assign t[55] = t[69] ^ t[70];
  assign t[56] = t[62] & t[71];
  assign t[57] = t[63] & t[72];
  assign t[58] = t[60] ^ t[64];
  assign t[59] = t[54] ^ t[67];
  assign t[5] = t[9] ? t[137] : x[3];
  assign t[60] = t[73] ^ t[74];
  assign t[61] = t[13] ? t[156] : t[75];
  assign t[62] = t[76] ^ t[77];
  assign t[63] = t[78] ^ t[79];
  assign t[64] = t[80] ^ t[81];
  assign t[65] = t[157] ^ t[158];
  assign t[66] = t[159] ^ t[160];
  assign t[67] = t[82] ^ t[70];
  assign t[68] = t[83] ^ t[51];
  assign t[69] = t[13] ? t[161] : t[84];
  assign t[6] = ~(t[10] ^ t[138]);
  assign t[70] = t[13] ? t[162] : t[85];
  assign t[71] = t[86] ^ t[53];
  assign t[72] = t[87] ^ t[88];
  assign t[73] = t[89] ^ t[90];
  assign t[74] = t[91] & t[92];
  assign t[75] = t[163] ^ t[138];
  assign t[76] = t[93] ^ t[94];
  assign t[77] = t[95] & t[96];
  assign t[78] = t[96] & t[97];
  assign t[79] = t[96] ^ t[98];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[92] & t[99];
  assign t[81] = t[92] ^ t[98];
  assign t[82] = t[13] ? t[164] : t[100];
  assign t[83] = t[13] ? t[165] : t[101];
  assign t[84] = t[166] ^ t[167];
  assign t[85] = t[168] ^ t[169];
  assign t[86] = t[61] ^ t[87];
  assign t[87] = t[102] ^ t[83];
  assign t[88] = t[70] ^ t[61];
  assign t[89] = t[103] ^ t[94];
  assign t[8] = ~(t[13]);
  assign t[90] = t[104] ^ t[71];
  assign t[91] = t[76] ^ t[98];
  assign t[92] = t[105] ^ t[73];
  assign t[93] = t[106] ^ t[107];
  assign t[94] = t[108] ^ t[109];
  assign t[95] = t[73] ^ t[98];
  assign t[96] = t[110] ^ t[76];
  assign t[97] = t[110] & t[73];
  assign t[98] = t[105] & t[110];
  assign t[99] = t[76] & t[105];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [120:0] x;
 output y;

 wire [414:0] t;
  assign t[0] = t[1] ? t[2] : t[135];
  assign t[100] = t[116] ^ t[57];
  assign t[101] = t[117] ^ t[118];
  assign t[102] = t[73] ^ t[64];
  assign t[103] = t[83] ^ t[82];
  assign t[104] = t[103] & t[119];
  assign t[105] = t[103] ^ t[64];
  assign t[106] = t[120] ^ t[121];
  assign t[107] = t[122] ^ t[78];
  assign t[108] = t[122] & t[78];
  assign t[109] = t[53] & t[123];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[13] ? t[171] : t[124];
  assign t[111] = t[172] ^ t[137];
  assign t[112] = t[125] ^ t[121];
  assign t[113] = t[126] & t[127];
  assign t[114] = t[55] & t[59];
  assign t[115] = t[128] ^ t[129];
  assign t[116] = t[53] ^ t[130];
  assign t[117] = t[131] ^ t[129];
  assign t[118] = t[58] & t[38];
  assign t[119] = t[73] & t[83];
  assign t[11] = ~(t[17]);
  assign t[120] = t[130] & t[50];
  assign t[121] = t[132] & t[96];
  assign t[122] = t[69] ^ t[72];
  assign t[123] = t[94] ^ t[133];
  assign t[124] = t[173] ^ t[174];
  assign t[125] = t[96] ^ t[133];
  assign t[126] = t[122] ^ t[58];
  assign t[127] = t[50] ^ t[96];
  assign t[128] = t[116] & t[57];
  assign t[129] = t[80] & t[75];
  assign t[12] = t[138] & t[18];
  assign t[130] = t[51] ^ t[134];
  assign t[131] = t[80] ^ t[75];
  assign t[132] = t[80] ^ t[55];
  assign t[133] = t[66] ^ t[72];
  assign t[134] = t[70] ^ t[50];
  assign t[135] = (t[175]);
  assign t[136] = (t[176]);
  assign t[137] = (t[177]);
  assign t[138] = (t[178]);
  assign t[139] = (t[179]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[180]);
  assign t[141] = (t[181]);
  assign t[142] = (t[182]);
  assign t[143] = (t[183]);
  assign t[144] = (t[184]);
  assign t[145] = (t[185]);
  assign t[146] = (t[186]);
  assign t[147] = (t[187]);
  assign t[148] = (t[188]);
  assign t[149] = (t[189]);
  assign t[14] = ~(t[138]);
  assign t[150] = (t[190]);
  assign t[151] = (t[191]);
  assign t[152] = (t[192]);
  assign t[153] = (t[193]);
  assign t[154] = (t[194]);
  assign t[155] = (t[195]);
  assign t[156] = (t[196]);
  assign t[157] = (t[197]);
  assign t[158] = (t[198]);
  assign t[159] = (t[199]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[200]);
  assign t[161] = (t[201]);
  assign t[162] = (t[202]);
  assign t[163] = (t[203]);
  assign t[164] = (t[204]);
  assign t[165] = (t[205]);
  assign t[166] = (t[206]);
  assign t[167] = (t[207]);
  assign t[168] = (t[208]);
  assign t[169] = (t[209]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (t[210]);
  assign t[171] = (t[211]);
  assign t[172] = (t[212]);
  assign t[173] = (t[213]);
  assign t[174] = (t[214]);
  assign t[175] = t[215] ^ x[2];
  assign t[176] = t[216] ^ x[6];
  assign t[177] = t[217] ^ x[9];
  assign t[178] = t[218] ^ x[12];
  assign t[179] = t[219] ^ x[15];
  assign t[17] = ~(t[138] & t[25]);
  assign t[180] = t[220] ^ x[18];
  assign t[181] = t[221] ^ x[21];
  assign t[182] = t[222] ^ x[24];
  assign t[183] = t[223] ^ x[27];
  assign t[184] = t[224] ^ x[30];
  assign t[185] = t[225] ^ x[33];
  assign t[186] = t[226] ^ x[36];
  assign t[187] = t[227] ^ x[39];
  assign t[188] = t[228] ^ x[42];
  assign t[189] = t[229] ^ x[45];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[230] ^ x[48];
  assign t[191] = t[231] ^ x[51];
  assign t[192] = t[232] ^ x[54];
  assign t[193] = t[233] ^ x[57];
  assign t[194] = t[234] ^ x[60];
  assign t[195] = t[235] ^ x[63];
  assign t[196] = t[236] ^ x[66];
  assign t[197] = t[237] ^ x[69];
  assign t[198] = t[238] ^ x[72];
  assign t[199] = t[239] ^ x[75];
  assign t[19] = ~(t[139]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[78];
  assign t[201] = t[241] ^ x[81];
  assign t[202] = t[242] ^ x[84];
  assign t[203] = t[243] ^ x[87];
  assign t[204] = t[244] ^ x[90];
  assign t[205] = t[245] ^ x[93];
  assign t[206] = t[246] ^ x[96];
  assign t[207] = t[247] ^ x[99];
  assign t[208] = t[248] ^ x[102];
  assign t[209] = t[249] ^ x[105];
  assign t[20] = ~(t[138]);
  assign t[210] = t[250] ^ x[108];
  assign t[211] = t[251] ^ x[111];
  assign t[212] = t[252] ^ x[114];
  assign t[213] = t[253] ^ x[117];
  assign t[214] = t[254] ^ x[120];
  assign t[215] = (t[255] & ~t[256]);
  assign t[216] = (t[257] & ~t[258]);
  assign t[217] = (t[259] & ~t[260]);
  assign t[218] = (t[261] & ~t[262]);
  assign t[219] = (t[263] & ~t[264]);
  assign t[21] = ~(t[140]);
  assign t[220] = (t[265] & ~t[266]);
  assign t[221] = (t[267] & ~t[268]);
  assign t[222] = (t[269] & ~t[270]);
  assign t[223] = (t[271] & ~t[272]);
  assign t[224] = (t[273] & ~t[274]);
  assign t[225] = (t[275] & ~t[276]);
  assign t[226] = (t[277] & ~t[278]);
  assign t[227] = (t[279] & ~t[280]);
  assign t[228] = (t[281] & ~t[282]);
  assign t[229] = (t[283] & ~t[284]);
  assign t[22] = ~(t[141]);
  assign t[230] = (t[285] & ~t[286]);
  assign t[231] = (t[287] & ~t[288]);
  assign t[232] = (t[289] & ~t[290]);
  assign t[233] = (t[291] & ~t[292]);
  assign t[234] = (t[293] & ~t[294]);
  assign t[235] = (t[295] & ~t[296]);
  assign t[236] = (t[297] & ~t[298]);
  assign t[237] = (t[299] & ~t[300]);
  assign t[238] = (t[301] & ~t[302]);
  assign t[239] = (t[303] & ~t[304]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[305] & ~t[306]);
  assign t[241] = (t[307] & ~t[308]);
  assign t[242] = (t[309] & ~t[310]);
  assign t[243] = (t[311] & ~t[312]);
  assign t[244] = (t[313] & ~t[314]);
  assign t[245] = (t[315] & ~t[316]);
  assign t[246] = (t[317] & ~t[318]);
  assign t[247] = (t[319] & ~t[320]);
  assign t[248] = (t[321] & ~t[322]);
  assign t[249] = (t[323] & ~t[324]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[325] & ~t[326]);
  assign t[251] = (t[327] & ~t[328]);
  assign t[252] = (t[329] & ~t[330]);
  assign t[253] = (t[331] & ~t[332]);
  assign t[254] = (t[333] & ~t[334]);
  assign t[255] = t[335] ^ x[2];
  assign t[256] = t[336] ^ x[1];
  assign t[257] = t[337] ^ x[6];
  assign t[258] = t[338] ^ x[5];
  assign t[259] = t[339] ^ x[9];
  assign t[25] = ~(t[142] | t[32]);
  assign t[260] = t[340] ^ x[8];
  assign t[261] = t[341] ^ x[12];
  assign t[262] = t[342] ^ x[11];
  assign t[263] = t[343] ^ x[15];
  assign t[264] = t[344] ^ x[14];
  assign t[265] = t[345] ^ x[18];
  assign t[266] = t[346] ^ x[17];
  assign t[267] = t[347] ^ x[21];
  assign t[268] = t[348] ^ x[20];
  assign t[269] = t[349] ^ x[24];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[350] ^ x[23];
  assign t[271] = t[351] ^ x[27];
  assign t[272] = t[352] ^ x[26];
  assign t[273] = t[353] ^ x[30];
  assign t[274] = t[354] ^ x[29];
  assign t[275] = t[355] ^ x[33];
  assign t[276] = t[356] ^ x[32];
  assign t[277] = t[357] ^ x[36];
  assign t[278] = t[358] ^ x[35];
  assign t[279] = t[359] ^ x[39];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[360] ^ x[38];
  assign t[281] = t[361] ^ x[42];
  assign t[282] = t[362] ^ x[41];
  assign t[283] = t[363] ^ x[45];
  assign t[284] = t[364] ^ x[44];
  assign t[285] = t[365] ^ x[48];
  assign t[286] = t[366] ^ x[47];
  assign t[287] = t[367] ^ x[51];
  assign t[288] = t[368] ^ x[50];
  assign t[289] = t[369] ^ x[54];
  assign t[28] = t[37] & t[38];
  assign t[290] = t[370] ^ x[53];
  assign t[291] = t[371] ^ x[57];
  assign t[292] = t[372] ^ x[56];
  assign t[293] = t[373] ^ x[60];
  assign t[294] = t[374] ^ x[59];
  assign t[295] = t[375] ^ x[63];
  assign t[296] = t[376] ^ x[62];
  assign t[297] = t[377] ^ x[66];
  assign t[298] = t[378] ^ x[65];
  assign t[299] = t[379] ^ x[69];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[380] ^ x[68];
  assign t[301] = t[381] ^ x[72];
  assign t[302] = t[382] ^ x[71];
  assign t[303] = t[383] ^ x[75];
  assign t[304] = t[384] ^ x[74];
  assign t[305] = t[385] ^ x[78];
  assign t[306] = t[386] ^ x[77];
  assign t[307] = t[387] ^ x[81];
  assign t[308] = t[388] ^ x[80];
  assign t[309] = t[389] ^ x[84];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[390] ^ x[83];
  assign t[311] = t[391] ^ x[87];
  assign t[312] = t[392] ^ x[86];
  assign t[313] = t[393] ^ x[90];
  assign t[314] = t[394] ^ x[89];
  assign t[315] = t[395] ^ x[93];
  assign t[316] = t[396] ^ x[92];
  assign t[317] = t[397] ^ x[96];
  assign t[318] = t[398] ^ x[95];
  assign t[319] = t[399] ^ x[99];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[400] ^ x[98];
  assign t[321] = t[401] ^ x[102];
  assign t[322] = t[402] ^ x[101];
  assign t[323] = t[403] ^ x[105];
  assign t[324] = t[404] ^ x[104];
  assign t[325] = t[405] ^ x[108];
  assign t[326] = t[406] ^ x[107];
  assign t[327] = t[407] ^ x[111];
  assign t[328] = t[408] ^ x[110];
  assign t[329] = t[409] ^ x[114];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[410] ^ x[113];
  assign t[331] = t[411] ^ x[117];
  assign t[332] = t[412] ^ x[116];
  assign t[333] = t[413] ^ x[120];
  assign t[334] = t[414] ^ x[119];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[4]);
  assign t[338] = (x[4]);
  assign t[339] = (x[7]);
  assign t[33] = ~(t[140] & t[143]);
  assign t[340] = (x[7]);
  assign t[341] = (x[10]);
  assign t[342] = (x[10]);
  assign t[343] = (x[13]);
  assign t[344] = (x[13]);
  assign t[345] = (x[16]);
  assign t[346] = (x[16]);
  assign t[347] = (x[19]);
  assign t[348] = (x[19]);
  assign t[349] = (x[22]);
  assign t[34] = ~(t[144] & t[145]);
  assign t[350] = (x[22]);
  assign t[351] = (x[25]);
  assign t[352] = (x[25]);
  assign t[353] = (x[28]);
  assign t[354] = (x[28]);
  assign t[355] = (x[31]);
  assign t[356] = (x[31]);
  assign t[357] = (x[34]);
  assign t[358] = (x[34]);
  assign t[359] = (x[37]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[37]);
  assign t[361] = (x[40]);
  assign t[362] = (x[40]);
  assign t[363] = (x[43]);
  assign t[364] = (x[43]);
  assign t[365] = (x[46]);
  assign t[366] = (x[46]);
  assign t[367] = (x[49]);
  assign t[368] = (x[49]);
  assign t[369] = (x[52]);
  assign t[36] = ~(t[146] & t[47]);
  assign t[370] = (x[52]);
  assign t[371] = (x[55]);
  assign t[372] = (x[55]);
  assign t[373] = (x[58]);
  assign t[374] = (x[58]);
  assign t[375] = (x[61]);
  assign t[376] = (x[61]);
  assign t[377] = (x[64]);
  assign t[378] = (x[64]);
  assign t[379] = (x[67]);
  assign t[37] = t[48] ^ t[49];
  assign t[380] = (x[67]);
  assign t[381] = (x[70]);
  assign t[382] = (x[70]);
  assign t[383] = (x[73]);
  assign t[384] = (x[73]);
  assign t[385] = (x[76]);
  assign t[386] = (x[76]);
  assign t[387] = (x[79]);
  assign t[388] = (x[79]);
  assign t[389] = (x[82]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[82]);
  assign t[391] = (x[85]);
  assign t[392] = (x[85]);
  assign t[393] = (x[88]);
  assign t[394] = (x[88]);
  assign t[395] = (x[91]);
  assign t[396] = (x[91]);
  assign t[397] = (x[94]);
  assign t[398] = (x[94]);
  assign t[399] = (x[97]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[97]);
  assign t[401] = (x[100]);
  assign t[402] = (x[100]);
  assign t[403] = (x[103]);
  assign t[404] = (x[103]);
  assign t[405] = (x[106]);
  assign t[406] = (x[106]);
  assign t[407] = (x[109]);
  assign t[408] = (x[109]);
  assign t[409] = (x[112]);
  assign t[40] = t[54] & t[55];
  assign t[410] = (x[112]);
  assign t[411] = (x[115]);
  assign t[412] = (x[115]);
  assign t[413] = (x[118]);
  assign t[414] = (x[118]);
  assign t[41] = t[56] & t[57];
  assign t[42] = t[37] & t[58];
  assign t[43] = t[54] & t[59];
  assign t[44] = t[60] ^ t[61];
  assign t[45] = ~(t[147] | t[148]);
  assign t[46] = ~(t[149] | t[150]);
  assign t[47] = ~(t[151]);
  assign t[48] = t[62] & t[63];
  assign t[49] = t[62] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[13] ? t[152] : t[65];
  assign t[51] = t[66] ^ t[67];
  assign t[52] = t[56] ^ t[68];
  assign t[53] = t[69] ^ t[70];
  assign t[54] = t[52] ^ t[71];
  assign t[55] = t[70] ^ t[72];
  assign t[56] = t[73] ^ t[74];
  assign t[57] = t[38] ^ t[75];
  assign t[58] = t[51] ^ t[76];
  assign t[59] = t[53] ^ t[77];
  assign t[5] = t[9] ? t[136] : x[3];
  assign t[60] = t[71] & t[78];
  assign t[61] = t[79] & t[80];
  assign t[62] = t[81] ^ t[73];
  assign t[63] = t[81] & t[82];
  assign t[64] = t[83] & t[81];
  assign t[65] = t[153] ^ t[154];
  assign t[66] = t[13] ? t[155] : t[84];
  assign t[67] = t[13] ? t[156] : t[85];
  assign t[68] = t[82] ^ t[86];
  assign t[69] = t[13] ? t[157] : t[87];
  assign t[6] = ~(t[10] ^ t[137]);
  assign t[70] = t[13] ? t[158] : t[88];
  assign t[71] = t[37] ^ t[89];
  assign t[72] = t[13] ? t[159] : t[90];
  assign t[73] = t[91] ^ t[92];
  assign t[74] = t[93] & t[62];
  assign t[75] = t[94] ^ t[77];
  assign t[76] = t[95] ^ t[50];
  assign t[77] = t[67] ^ t[72];
  assign t[78] = t[96] ^ t[51];
  assign t[79] = t[56] ^ t[37];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[69] ^ t[95];
  assign t[81] = t[97] ^ t[98];
  assign t[82] = t[99] ^ t[100];
  assign t[83] = t[101] ^ t[98];
  assign t[84] = t[160] ^ t[161];
  assign t[85] = t[162] ^ t[163];
  assign t[86] = t[102] & t[103];
  assign t[87] = t[164] ^ t[165];
  assign t[88] = t[166] ^ t[167];
  assign t[89] = t[104] ^ t[105];
  assign t[8] = ~(t[13]);
  assign t[90] = t[168] ^ t[169];
  assign t[91] = t[106] ^ t[107];
  assign t[92] = t[108] ^ t[109];
  assign t[93] = t[82] ^ t[64];
  assign t[94] = t[110] ^ t[95];
  assign t[95] = t[13] ? t[170] : t[111];
  assign t[96] = t[53] ^ t[94];
  assign t[97] = t[112] ^ t[113];
  assign t[98] = t[114] ^ t[109];
  assign t[99] = t[115] ^ t[92];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [120:0] x;
 output y;

 wire [414:0] t;
  assign t[0] = t[1] ? t[2] : t[135];
  assign t[100] = t[116] ^ t[57];
  assign t[101] = t[117] ^ t[118];
  assign t[102] = t[73] ^ t[64];
  assign t[103] = t[83] ^ t[82];
  assign t[104] = t[103] & t[119];
  assign t[105] = t[103] ^ t[64];
  assign t[106] = t[120] ^ t[121];
  assign t[107] = t[122] ^ t[78];
  assign t[108] = t[122] & t[78];
  assign t[109] = t[53] & t[123];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[13] ? t[171] : t[124];
  assign t[111] = t[172] ^ t[137];
  assign t[112] = t[125] ^ t[121];
  assign t[113] = t[126] & t[127];
  assign t[114] = t[55] & t[59];
  assign t[115] = t[128] ^ t[129];
  assign t[116] = t[53] ^ t[130];
  assign t[117] = t[131] ^ t[129];
  assign t[118] = t[58] & t[38];
  assign t[119] = t[73] & t[83];
  assign t[11] = ~(t[17]);
  assign t[120] = t[130] & t[50];
  assign t[121] = t[132] & t[96];
  assign t[122] = t[69] ^ t[72];
  assign t[123] = t[94] ^ t[133];
  assign t[124] = t[173] ^ t[174];
  assign t[125] = t[96] ^ t[133];
  assign t[126] = t[122] ^ t[58];
  assign t[127] = t[50] ^ t[96];
  assign t[128] = t[116] & t[57];
  assign t[129] = t[80] & t[75];
  assign t[12] = t[138] & t[18];
  assign t[130] = t[51] ^ t[134];
  assign t[131] = t[80] ^ t[75];
  assign t[132] = t[80] ^ t[55];
  assign t[133] = t[66] ^ t[72];
  assign t[134] = t[70] ^ t[50];
  assign t[135] = (t[175]);
  assign t[136] = (t[176]);
  assign t[137] = (t[177]);
  assign t[138] = (t[178]);
  assign t[139] = (t[179]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[180]);
  assign t[141] = (t[181]);
  assign t[142] = (t[182]);
  assign t[143] = (t[183]);
  assign t[144] = (t[184]);
  assign t[145] = (t[185]);
  assign t[146] = (t[186]);
  assign t[147] = (t[187]);
  assign t[148] = (t[188]);
  assign t[149] = (t[189]);
  assign t[14] = ~(t[138]);
  assign t[150] = (t[190]);
  assign t[151] = (t[191]);
  assign t[152] = (t[192]);
  assign t[153] = (t[193]);
  assign t[154] = (t[194]);
  assign t[155] = (t[195]);
  assign t[156] = (t[196]);
  assign t[157] = (t[197]);
  assign t[158] = (t[198]);
  assign t[159] = (t[199]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[200]);
  assign t[161] = (t[201]);
  assign t[162] = (t[202]);
  assign t[163] = (t[203]);
  assign t[164] = (t[204]);
  assign t[165] = (t[205]);
  assign t[166] = (t[206]);
  assign t[167] = (t[207]);
  assign t[168] = (t[208]);
  assign t[169] = (t[209]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (t[210]);
  assign t[171] = (t[211]);
  assign t[172] = (t[212]);
  assign t[173] = (t[213]);
  assign t[174] = (t[214]);
  assign t[175] = t[215] ^ x[2];
  assign t[176] = t[216] ^ x[6];
  assign t[177] = t[217] ^ x[9];
  assign t[178] = t[218] ^ x[12];
  assign t[179] = t[219] ^ x[15];
  assign t[17] = ~(t[138] & t[25]);
  assign t[180] = t[220] ^ x[18];
  assign t[181] = t[221] ^ x[21];
  assign t[182] = t[222] ^ x[24];
  assign t[183] = t[223] ^ x[27];
  assign t[184] = t[224] ^ x[30];
  assign t[185] = t[225] ^ x[33];
  assign t[186] = t[226] ^ x[36];
  assign t[187] = t[227] ^ x[39];
  assign t[188] = t[228] ^ x[42];
  assign t[189] = t[229] ^ x[45];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[230] ^ x[48];
  assign t[191] = t[231] ^ x[51];
  assign t[192] = t[232] ^ x[54];
  assign t[193] = t[233] ^ x[57];
  assign t[194] = t[234] ^ x[60];
  assign t[195] = t[235] ^ x[63];
  assign t[196] = t[236] ^ x[66];
  assign t[197] = t[237] ^ x[69];
  assign t[198] = t[238] ^ x[72];
  assign t[199] = t[239] ^ x[75];
  assign t[19] = ~(t[139]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[78];
  assign t[201] = t[241] ^ x[81];
  assign t[202] = t[242] ^ x[84];
  assign t[203] = t[243] ^ x[87];
  assign t[204] = t[244] ^ x[90];
  assign t[205] = t[245] ^ x[93];
  assign t[206] = t[246] ^ x[96];
  assign t[207] = t[247] ^ x[99];
  assign t[208] = t[248] ^ x[102];
  assign t[209] = t[249] ^ x[105];
  assign t[20] = ~(t[138]);
  assign t[210] = t[250] ^ x[108];
  assign t[211] = t[251] ^ x[111];
  assign t[212] = t[252] ^ x[114];
  assign t[213] = t[253] ^ x[117];
  assign t[214] = t[254] ^ x[120];
  assign t[215] = (t[255] & ~t[256]);
  assign t[216] = (t[257] & ~t[258]);
  assign t[217] = (t[259] & ~t[260]);
  assign t[218] = (t[261] & ~t[262]);
  assign t[219] = (t[263] & ~t[264]);
  assign t[21] = ~(t[140]);
  assign t[220] = (t[265] & ~t[266]);
  assign t[221] = (t[267] & ~t[268]);
  assign t[222] = (t[269] & ~t[270]);
  assign t[223] = (t[271] & ~t[272]);
  assign t[224] = (t[273] & ~t[274]);
  assign t[225] = (t[275] & ~t[276]);
  assign t[226] = (t[277] & ~t[278]);
  assign t[227] = (t[279] & ~t[280]);
  assign t[228] = (t[281] & ~t[282]);
  assign t[229] = (t[283] & ~t[284]);
  assign t[22] = ~(t[141]);
  assign t[230] = (t[285] & ~t[286]);
  assign t[231] = (t[287] & ~t[288]);
  assign t[232] = (t[289] & ~t[290]);
  assign t[233] = (t[291] & ~t[292]);
  assign t[234] = (t[293] & ~t[294]);
  assign t[235] = (t[295] & ~t[296]);
  assign t[236] = (t[297] & ~t[298]);
  assign t[237] = (t[299] & ~t[300]);
  assign t[238] = (t[301] & ~t[302]);
  assign t[239] = (t[303] & ~t[304]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[305] & ~t[306]);
  assign t[241] = (t[307] & ~t[308]);
  assign t[242] = (t[309] & ~t[310]);
  assign t[243] = (t[311] & ~t[312]);
  assign t[244] = (t[313] & ~t[314]);
  assign t[245] = (t[315] & ~t[316]);
  assign t[246] = (t[317] & ~t[318]);
  assign t[247] = (t[319] & ~t[320]);
  assign t[248] = (t[321] & ~t[322]);
  assign t[249] = (t[323] & ~t[324]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[325] & ~t[326]);
  assign t[251] = (t[327] & ~t[328]);
  assign t[252] = (t[329] & ~t[330]);
  assign t[253] = (t[331] & ~t[332]);
  assign t[254] = (t[333] & ~t[334]);
  assign t[255] = t[335] ^ x[2];
  assign t[256] = t[336] ^ x[1];
  assign t[257] = t[337] ^ x[6];
  assign t[258] = t[338] ^ x[5];
  assign t[259] = t[339] ^ x[9];
  assign t[25] = ~(t[142] | t[32]);
  assign t[260] = t[340] ^ x[8];
  assign t[261] = t[341] ^ x[12];
  assign t[262] = t[342] ^ x[11];
  assign t[263] = t[343] ^ x[15];
  assign t[264] = t[344] ^ x[14];
  assign t[265] = t[345] ^ x[18];
  assign t[266] = t[346] ^ x[17];
  assign t[267] = t[347] ^ x[21];
  assign t[268] = t[348] ^ x[20];
  assign t[269] = t[349] ^ x[24];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[350] ^ x[23];
  assign t[271] = t[351] ^ x[27];
  assign t[272] = t[352] ^ x[26];
  assign t[273] = t[353] ^ x[30];
  assign t[274] = t[354] ^ x[29];
  assign t[275] = t[355] ^ x[33];
  assign t[276] = t[356] ^ x[32];
  assign t[277] = t[357] ^ x[36];
  assign t[278] = t[358] ^ x[35];
  assign t[279] = t[359] ^ x[39];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[360] ^ x[38];
  assign t[281] = t[361] ^ x[42];
  assign t[282] = t[362] ^ x[41];
  assign t[283] = t[363] ^ x[45];
  assign t[284] = t[364] ^ x[44];
  assign t[285] = t[365] ^ x[48];
  assign t[286] = t[366] ^ x[47];
  assign t[287] = t[367] ^ x[51];
  assign t[288] = t[368] ^ x[50];
  assign t[289] = t[369] ^ x[54];
  assign t[28] = t[37] & t[38];
  assign t[290] = t[370] ^ x[53];
  assign t[291] = t[371] ^ x[57];
  assign t[292] = t[372] ^ x[56];
  assign t[293] = t[373] ^ x[60];
  assign t[294] = t[374] ^ x[59];
  assign t[295] = t[375] ^ x[63];
  assign t[296] = t[376] ^ x[62];
  assign t[297] = t[377] ^ x[66];
  assign t[298] = t[378] ^ x[65];
  assign t[299] = t[379] ^ x[69];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[380] ^ x[68];
  assign t[301] = t[381] ^ x[72];
  assign t[302] = t[382] ^ x[71];
  assign t[303] = t[383] ^ x[75];
  assign t[304] = t[384] ^ x[74];
  assign t[305] = t[385] ^ x[78];
  assign t[306] = t[386] ^ x[77];
  assign t[307] = t[387] ^ x[81];
  assign t[308] = t[388] ^ x[80];
  assign t[309] = t[389] ^ x[84];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[390] ^ x[83];
  assign t[311] = t[391] ^ x[87];
  assign t[312] = t[392] ^ x[86];
  assign t[313] = t[393] ^ x[90];
  assign t[314] = t[394] ^ x[89];
  assign t[315] = t[395] ^ x[93];
  assign t[316] = t[396] ^ x[92];
  assign t[317] = t[397] ^ x[96];
  assign t[318] = t[398] ^ x[95];
  assign t[319] = t[399] ^ x[99];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[400] ^ x[98];
  assign t[321] = t[401] ^ x[102];
  assign t[322] = t[402] ^ x[101];
  assign t[323] = t[403] ^ x[105];
  assign t[324] = t[404] ^ x[104];
  assign t[325] = t[405] ^ x[108];
  assign t[326] = t[406] ^ x[107];
  assign t[327] = t[407] ^ x[111];
  assign t[328] = t[408] ^ x[110];
  assign t[329] = t[409] ^ x[114];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[410] ^ x[113];
  assign t[331] = t[411] ^ x[117];
  assign t[332] = t[412] ^ x[116];
  assign t[333] = t[413] ^ x[120];
  assign t[334] = t[414] ^ x[119];
  assign t[335] = (x[0]);
  assign t[336] = (x[0]);
  assign t[337] = (x[4]);
  assign t[338] = (x[4]);
  assign t[339] = (x[7]);
  assign t[33] = ~(t[140] & t[143]);
  assign t[340] = (x[7]);
  assign t[341] = (x[10]);
  assign t[342] = (x[10]);
  assign t[343] = (x[13]);
  assign t[344] = (x[13]);
  assign t[345] = (x[16]);
  assign t[346] = (x[16]);
  assign t[347] = (x[19]);
  assign t[348] = (x[19]);
  assign t[349] = (x[22]);
  assign t[34] = ~(t[144] & t[145]);
  assign t[350] = (x[22]);
  assign t[351] = (x[25]);
  assign t[352] = (x[25]);
  assign t[353] = (x[28]);
  assign t[354] = (x[28]);
  assign t[355] = (x[31]);
  assign t[356] = (x[31]);
  assign t[357] = (x[34]);
  assign t[358] = (x[34]);
  assign t[359] = (x[37]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[37]);
  assign t[361] = (x[40]);
  assign t[362] = (x[40]);
  assign t[363] = (x[43]);
  assign t[364] = (x[43]);
  assign t[365] = (x[46]);
  assign t[366] = (x[46]);
  assign t[367] = (x[49]);
  assign t[368] = (x[49]);
  assign t[369] = (x[52]);
  assign t[36] = ~(t[146] & t[47]);
  assign t[370] = (x[52]);
  assign t[371] = (x[55]);
  assign t[372] = (x[55]);
  assign t[373] = (x[58]);
  assign t[374] = (x[58]);
  assign t[375] = (x[61]);
  assign t[376] = (x[61]);
  assign t[377] = (x[64]);
  assign t[378] = (x[64]);
  assign t[379] = (x[67]);
  assign t[37] = t[48] ^ t[49];
  assign t[380] = (x[67]);
  assign t[381] = (x[70]);
  assign t[382] = (x[70]);
  assign t[383] = (x[73]);
  assign t[384] = (x[73]);
  assign t[385] = (x[76]);
  assign t[386] = (x[76]);
  assign t[387] = (x[79]);
  assign t[388] = (x[79]);
  assign t[389] = (x[82]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[82]);
  assign t[391] = (x[85]);
  assign t[392] = (x[85]);
  assign t[393] = (x[88]);
  assign t[394] = (x[88]);
  assign t[395] = (x[91]);
  assign t[396] = (x[91]);
  assign t[397] = (x[94]);
  assign t[398] = (x[94]);
  assign t[399] = (x[97]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[97]);
  assign t[401] = (x[100]);
  assign t[402] = (x[100]);
  assign t[403] = (x[103]);
  assign t[404] = (x[103]);
  assign t[405] = (x[106]);
  assign t[406] = (x[106]);
  assign t[407] = (x[109]);
  assign t[408] = (x[109]);
  assign t[409] = (x[112]);
  assign t[40] = t[54] & t[55];
  assign t[410] = (x[112]);
  assign t[411] = (x[115]);
  assign t[412] = (x[115]);
  assign t[413] = (x[118]);
  assign t[414] = (x[118]);
  assign t[41] = t[56] & t[57];
  assign t[42] = t[37] & t[58];
  assign t[43] = t[54] & t[59];
  assign t[44] = t[60] ^ t[61];
  assign t[45] = ~(t[147] | t[148]);
  assign t[46] = ~(t[149] | t[150]);
  assign t[47] = ~(t[151]);
  assign t[48] = t[62] & t[63];
  assign t[49] = t[62] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[13] ? t[152] : t[65];
  assign t[51] = t[66] ^ t[67];
  assign t[52] = t[56] ^ t[68];
  assign t[53] = t[69] ^ t[70];
  assign t[54] = t[52] ^ t[71];
  assign t[55] = t[70] ^ t[72];
  assign t[56] = t[73] ^ t[74];
  assign t[57] = t[38] ^ t[75];
  assign t[58] = t[51] ^ t[76];
  assign t[59] = t[53] ^ t[77];
  assign t[5] = t[9] ? t[136] : x[3];
  assign t[60] = t[71] & t[78];
  assign t[61] = t[79] & t[80];
  assign t[62] = t[81] ^ t[73];
  assign t[63] = t[81] & t[82];
  assign t[64] = t[83] & t[81];
  assign t[65] = t[153] ^ t[154];
  assign t[66] = t[13] ? t[155] : t[84];
  assign t[67] = t[13] ? t[156] : t[85];
  assign t[68] = t[82] ^ t[86];
  assign t[69] = t[13] ? t[157] : t[87];
  assign t[6] = ~(t[10] ^ t[137]);
  assign t[70] = t[13] ? t[158] : t[88];
  assign t[71] = t[37] ^ t[89];
  assign t[72] = t[13] ? t[159] : t[90];
  assign t[73] = t[91] ^ t[92];
  assign t[74] = t[93] & t[62];
  assign t[75] = t[94] ^ t[77];
  assign t[76] = t[95] ^ t[50];
  assign t[77] = t[67] ^ t[72];
  assign t[78] = t[96] ^ t[51];
  assign t[79] = t[56] ^ t[37];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[69] ^ t[95];
  assign t[81] = t[97] ^ t[98];
  assign t[82] = t[99] ^ t[100];
  assign t[83] = t[101] ^ t[98];
  assign t[84] = t[160] ^ t[161];
  assign t[85] = t[162] ^ t[163];
  assign t[86] = t[102] & t[103];
  assign t[87] = t[164] ^ t[165];
  assign t[88] = t[166] ^ t[167];
  assign t[89] = t[104] ^ t[105];
  assign t[8] = ~(t[13]);
  assign t[90] = t[168] ^ t[169];
  assign t[91] = t[106] ^ t[107];
  assign t[92] = t[108] ^ t[109];
  assign t[93] = t[82] ^ t[64];
  assign t[94] = t[110] ^ t[95];
  assign t[95] = t[13] ? t[170] : t[111];
  assign t[96] = t[53] ^ t[94];
  assign t[97] = t[112] ^ t[113];
  assign t[98] = t[114] ^ t[109];
  assign t[99] = t[115] ^ t[92];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind236(x, y);
 input [120:0] x;
 output y;

 wire [423:0] t;
  assign t[0] = t[1] ? t[2] : t[144];
  assign t[100] = t[120] ^ t[78];
  assign t[101] = t[13] ? t[172] : t[121];
  assign t[102] = t[95] & t[122];
  assign t[103] = t[95] ^ t[116];
  assign t[104] = t[100] & t[123];
  assign t[105] = t[100] ^ t[116];
  assign t[106] = t[89] ^ t[66];
  assign t[107] = t[80] ^ t[124];
  assign t[108] = t[13] ? t[173] : t[125];
  assign t[109] = t[174] ^ t[175];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[176] ^ t[177];
  assign t[111] = t[178] ^ t[179];
  assign t[112] = t[126] ^ t[127];
  assign t[113] = t[106] ^ t[71];
  assign t[114] = t[106] & t[71];
  assign t[115] = t[69] & t[128];
  assign t[116] = t[120] & t[117];
  assign t[117] = t[129] ^ t[130];
  assign t[118] = t[131] ^ t[132];
  assign t[119] = t[83] ^ t[68];
  assign t[11] = ~(t[17]);
  assign t[120] = t[133] ^ t[130];
  assign t[121] = t[180] ^ t[181];
  assign t[122] = t[117] & t[78];
  assign t[123] = t[73] & t[120];
  assign t[124] = t[91] ^ t[77];
  assign t[125] = t[182] ^ t[183];
  assign t[126] = t[60] & t[77];
  assign t[127] = t[134] & t[76];
  assign t[128] = t[88] ^ t[135];
  assign t[129] = t[136] ^ t[137];
  assign t[12] = t[147] & t[18];
  assign t[130] = t[138] ^ t[115];
  assign t[131] = t[56] & t[119];
  assign t[132] = t[72] & t[68];
  assign t[133] = t[139] ^ t[140];
  assign t[134] = t[72] ^ t[49];
  assign t[135] = t[101] ^ t[66];
  assign t[136] = t[141] ^ t[127];
  assign t[137] = t[85] & t[142];
  assign t[138] = t[49] & t[52];
  assign t[139] = t[143] ^ t[132];
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = t[107] & t[83];
  assign t[141] = t[76] ^ t[135];
  assign t[142] = t[77] ^ t[76];
  assign t[143] = t[72] ^ t[68];
  assign t[144] = (t[184]);
  assign t[145] = (t[185]);
  assign t[146] = (t[186]);
  assign t[147] = (t[187]);
  assign t[148] = (t[188]);
  assign t[149] = (t[189]);
  assign t[14] = ~(t[147]);
  assign t[150] = (t[190]);
  assign t[151] = (t[191]);
  assign t[152] = (t[192]);
  assign t[153] = (t[193]);
  assign t[154] = (t[194]);
  assign t[155] = (t[195]);
  assign t[156] = (t[196]);
  assign t[157] = (t[197]);
  assign t[158] = (t[198]);
  assign t[159] = (t[199]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[200]);
  assign t[161] = (t[201]);
  assign t[162] = (t[202]);
  assign t[163] = (t[203]);
  assign t[164] = (t[204]);
  assign t[165] = (t[205]);
  assign t[166] = (t[206]);
  assign t[167] = (t[207]);
  assign t[168] = (t[208]);
  assign t[169] = (t[209]);
  assign t[16] = t[23] ^ t[24];
  assign t[170] = (t[210]);
  assign t[171] = (t[211]);
  assign t[172] = (t[212]);
  assign t[173] = (t[213]);
  assign t[174] = (t[214]);
  assign t[175] = (t[215]);
  assign t[176] = (t[216]);
  assign t[177] = (t[217]);
  assign t[178] = (t[218]);
  assign t[179] = (t[219]);
  assign t[17] = ~(t[147] & t[25]);
  assign t[180] = (t[220]);
  assign t[181] = (t[221]);
  assign t[182] = (t[222]);
  assign t[183] = (t[223]);
  assign t[184] = t[224] ^ x[2];
  assign t[185] = t[225] ^ x[6];
  assign t[186] = t[226] ^ x[9];
  assign t[187] = t[227] ^ x[12];
  assign t[188] = t[228] ^ x[15];
  assign t[189] = t[229] ^ x[18];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[230] ^ x[21];
  assign t[191] = t[231] ^ x[24];
  assign t[192] = t[232] ^ x[27];
  assign t[193] = t[233] ^ x[30];
  assign t[194] = t[234] ^ x[33];
  assign t[195] = t[235] ^ x[36];
  assign t[196] = t[236] ^ x[39];
  assign t[197] = t[237] ^ x[42];
  assign t[198] = t[238] ^ x[45];
  assign t[199] = t[239] ^ x[48];
  assign t[19] = ~(t[148]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[51];
  assign t[201] = t[241] ^ x[54];
  assign t[202] = t[242] ^ x[57];
  assign t[203] = t[243] ^ x[60];
  assign t[204] = t[244] ^ x[63];
  assign t[205] = t[245] ^ x[66];
  assign t[206] = t[246] ^ x[69];
  assign t[207] = t[247] ^ x[72];
  assign t[208] = t[248] ^ x[75];
  assign t[209] = t[249] ^ x[78];
  assign t[20] = ~(t[147]);
  assign t[210] = t[250] ^ x[81];
  assign t[211] = t[251] ^ x[84];
  assign t[212] = t[252] ^ x[87];
  assign t[213] = t[253] ^ x[90];
  assign t[214] = t[254] ^ x[93];
  assign t[215] = t[255] ^ x[96];
  assign t[216] = t[256] ^ x[99];
  assign t[217] = t[257] ^ x[102];
  assign t[218] = t[258] ^ x[105];
  assign t[219] = t[259] ^ x[108];
  assign t[21] = ~(t[149]);
  assign t[220] = t[260] ^ x[111];
  assign t[221] = t[261] ^ x[114];
  assign t[222] = t[262] ^ x[117];
  assign t[223] = t[263] ^ x[120];
  assign t[224] = (t[264] & ~t[265]);
  assign t[225] = (t[266] & ~t[267]);
  assign t[226] = (t[268] & ~t[269]);
  assign t[227] = (t[270] & ~t[271]);
  assign t[228] = (t[272] & ~t[273]);
  assign t[229] = (t[274] & ~t[275]);
  assign t[22] = ~(t[150]);
  assign t[230] = (t[276] & ~t[277]);
  assign t[231] = (t[278] & ~t[279]);
  assign t[232] = (t[280] & ~t[281]);
  assign t[233] = (t[282] & ~t[283]);
  assign t[234] = (t[284] & ~t[285]);
  assign t[235] = (t[286] & ~t[287]);
  assign t[236] = (t[288] & ~t[289]);
  assign t[237] = (t[290] & ~t[291]);
  assign t[238] = (t[292] & ~t[293]);
  assign t[239] = (t[294] & ~t[295]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[296] & ~t[297]);
  assign t[241] = (t[298] & ~t[299]);
  assign t[242] = (t[300] & ~t[301]);
  assign t[243] = (t[302] & ~t[303]);
  assign t[244] = (t[304] & ~t[305]);
  assign t[245] = (t[306] & ~t[307]);
  assign t[246] = (t[308] & ~t[309]);
  assign t[247] = (t[310] & ~t[311]);
  assign t[248] = (t[312] & ~t[313]);
  assign t[249] = (t[314] & ~t[315]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[316] & ~t[317]);
  assign t[251] = (t[318] & ~t[319]);
  assign t[252] = (t[320] & ~t[321]);
  assign t[253] = (t[322] & ~t[323]);
  assign t[254] = (t[324] & ~t[325]);
  assign t[255] = (t[326] & ~t[327]);
  assign t[256] = (t[328] & ~t[329]);
  assign t[257] = (t[330] & ~t[331]);
  assign t[258] = (t[332] & ~t[333]);
  assign t[259] = (t[334] & ~t[335]);
  assign t[25] = ~(t[151] | t[32]);
  assign t[260] = (t[336] & ~t[337]);
  assign t[261] = (t[338] & ~t[339]);
  assign t[262] = (t[340] & ~t[341]);
  assign t[263] = (t[342] & ~t[343]);
  assign t[264] = t[344] ^ x[2];
  assign t[265] = t[345] ^ x[1];
  assign t[266] = t[346] ^ x[6];
  assign t[267] = t[347] ^ x[5];
  assign t[268] = t[348] ^ x[9];
  assign t[269] = t[349] ^ x[8];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[350] ^ x[12];
  assign t[271] = t[351] ^ x[11];
  assign t[272] = t[352] ^ x[15];
  assign t[273] = t[353] ^ x[14];
  assign t[274] = t[354] ^ x[18];
  assign t[275] = t[355] ^ x[17];
  assign t[276] = t[356] ^ x[21];
  assign t[277] = t[357] ^ x[20];
  assign t[278] = t[358] ^ x[24];
  assign t[279] = t[359] ^ x[23];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[360] ^ x[27];
  assign t[281] = t[361] ^ x[26];
  assign t[282] = t[362] ^ x[30];
  assign t[283] = t[363] ^ x[29];
  assign t[284] = t[364] ^ x[33];
  assign t[285] = t[365] ^ x[32];
  assign t[286] = t[366] ^ x[36];
  assign t[287] = t[367] ^ x[35];
  assign t[288] = t[368] ^ x[39];
  assign t[289] = t[369] ^ x[38];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[370] ^ x[42];
  assign t[291] = t[371] ^ x[41];
  assign t[292] = t[372] ^ x[45];
  assign t[293] = t[373] ^ x[44];
  assign t[294] = t[374] ^ x[48];
  assign t[295] = t[375] ^ x[47];
  assign t[296] = t[376] ^ x[51];
  assign t[297] = t[377] ^ x[50];
  assign t[298] = t[378] ^ x[54];
  assign t[299] = t[379] ^ x[53];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[380] ^ x[57];
  assign t[301] = t[381] ^ x[56];
  assign t[302] = t[382] ^ x[60];
  assign t[303] = t[383] ^ x[59];
  assign t[304] = t[384] ^ x[63];
  assign t[305] = t[385] ^ x[62];
  assign t[306] = t[386] ^ x[66];
  assign t[307] = t[387] ^ x[65];
  assign t[308] = t[388] ^ x[69];
  assign t[309] = t[389] ^ x[68];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[390] ^ x[72];
  assign t[311] = t[391] ^ x[71];
  assign t[312] = t[392] ^ x[75];
  assign t[313] = t[393] ^ x[74];
  assign t[314] = t[394] ^ x[78];
  assign t[315] = t[395] ^ x[77];
  assign t[316] = t[396] ^ x[81];
  assign t[317] = t[397] ^ x[80];
  assign t[318] = t[398] ^ x[84];
  assign t[319] = t[399] ^ x[83];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[400] ^ x[87];
  assign t[321] = t[401] ^ x[86];
  assign t[322] = t[402] ^ x[90];
  assign t[323] = t[403] ^ x[89];
  assign t[324] = t[404] ^ x[93];
  assign t[325] = t[405] ^ x[92];
  assign t[326] = t[406] ^ x[96];
  assign t[327] = t[407] ^ x[95];
  assign t[328] = t[408] ^ x[99];
  assign t[329] = t[409] ^ x[98];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[410] ^ x[102];
  assign t[331] = t[411] ^ x[101];
  assign t[332] = t[412] ^ x[105];
  assign t[333] = t[413] ^ x[104];
  assign t[334] = t[414] ^ x[108];
  assign t[335] = t[415] ^ x[107];
  assign t[336] = t[416] ^ x[111];
  assign t[337] = t[417] ^ x[110];
  assign t[338] = t[418] ^ x[114];
  assign t[339] = t[419] ^ x[113];
  assign t[33] = ~(t[152] & t[153]);
  assign t[340] = t[420] ^ x[117];
  assign t[341] = t[421] ^ x[116];
  assign t[342] = t[422] ^ x[120];
  assign t[343] = t[423] ^ x[119];
  assign t[344] = (x[0]);
  assign t[345] = (x[0]);
  assign t[346] = (x[4]);
  assign t[347] = (x[4]);
  assign t[348] = (x[7]);
  assign t[349] = (x[7]);
  assign t[34] = ~(t[154] & t[149]);
  assign t[350] = (x[10]);
  assign t[351] = (x[10]);
  assign t[352] = (x[13]);
  assign t[353] = (x[13]);
  assign t[354] = (x[16]);
  assign t[355] = (x[16]);
  assign t[356] = (x[19]);
  assign t[357] = (x[19]);
  assign t[358] = (x[22]);
  assign t[359] = (x[22]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[25]);
  assign t[361] = (x[25]);
  assign t[362] = (x[28]);
  assign t[363] = (x[28]);
  assign t[364] = (x[31]);
  assign t[365] = (x[31]);
  assign t[366] = (x[34]);
  assign t[367] = (x[34]);
  assign t[368] = (x[37]);
  assign t[369] = (x[37]);
  assign t[36] = ~(t[155] & t[47]);
  assign t[370] = (x[40]);
  assign t[371] = (x[40]);
  assign t[372] = (x[43]);
  assign t[373] = (x[43]);
  assign t[374] = (x[46]);
  assign t[375] = (x[46]);
  assign t[376] = (x[49]);
  assign t[377] = (x[49]);
  assign t[378] = (x[52]);
  assign t[379] = (x[52]);
  assign t[37] = t[48] & t[49];
  assign t[380] = (x[55]);
  assign t[381] = (x[55]);
  assign t[382] = (x[58]);
  assign t[383] = (x[58]);
  assign t[384] = (x[61]);
  assign t[385] = (x[61]);
  assign t[386] = (x[64]);
  assign t[387] = (x[64]);
  assign t[388] = (x[67]);
  assign t[389] = (x[67]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[70]);
  assign t[391] = (x[70]);
  assign t[392] = (x[73]);
  assign t[393] = (x[73]);
  assign t[394] = (x[76]);
  assign t[395] = (x[76]);
  assign t[396] = (x[79]);
  assign t[397] = (x[79]);
  assign t[398] = (x[82]);
  assign t[399] = (x[82]);
  assign t[39] = t[48] & t[52];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[85]);
  assign t[401] = (x[85]);
  assign t[402] = (x[88]);
  assign t[403] = (x[88]);
  assign t[404] = (x[91]);
  assign t[405] = (x[91]);
  assign t[406] = (x[94]);
  assign t[407] = (x[94]);
  assign t[408] = (x[97]);
  assign t[409] = (x[97]);
  assign t[40] = t[53] ^ t[54];
  assign t[410] = (x[100]);
  assign t[411] = (x[100]);
  assign t[412] = (x[103]);
  assign t[413] = (x[103]);
  assign t[414] = (x[106]);
  assign t[415] = (x[106]);
  assign t[416] = (x[109]);
  assign t[417] = (x[109]);
  assign t[418] = (x[112]);
  assign t[419] = (x[112]);
  assign t[41] = t[55] & t[56];
  assign t[420] = (x[115]);
  assign t[421] = (x[115]);
  assign t[422] = (x[118]);
  assign t[423] = (x[118]);
  assign t[42] = t[57] ^ t[58];
  assign t[43] = t[59] & t[60];
  assign t[44] = t[61] ^ t[62];
  assign t[45] = ~(t[156] | t[157]);
  assign t[46] = ~(t[158] | t[159]);
  assign t[47] = ~(t[160]);
  assign t[48] = t[63] ^ t[64];
  assign t[49] = t[65] ^ t[66];
  assign t[4] = ~(t[8]);
  assign t[50] = t[67] & t[68];
  assign t[51] = t[63] & t[69];
  assign t[52] = t[69] ^ t[70];
  assign t[53] = t[64] & t[71];
  assign t[54] = t[67] & t[72];
  assign t[55] = t[73] ^ t[74];
  assign t[56] = t[69] ^ t[60];
  assign t[57] = t[75] & t[76];
  assign t[58] = t[59] & t[77];
  assign t[59] = t[78] ^ t[79];
  assign t[5] = t[9] ? t[145] : x[3];
  assign t[60] = t[80] ^ t[81];
  assign t[61] = t[82] & t[83];
  assign t[62] = t[84] & t[85];
  assign t[63] = t[55] ^ t[59];
  assign t[64] = t[82] ^ t[84];
  assign t[65] = t[13] ? t[161] : t[86];
  assign t[66] = t[13] ? t[162] : t[87];
  assign t[67] = t[55] ^ t[82];
  assign t[68] = t[88] ^ t[70];
  assign t[69] = t[89] ^ t[65];
  assign t[6] = ~(t[10] ^ t[146]);
  assign t[70] = t[90] ^ t[66];
  assign t[71] = t[76] ^ t[80];
  assign t[72] = t[89] ^ t[91];
  assign t[73] = t[92] ^ t[93];
  assign t[74] = t[94] & t[95];
  assign t[75] = t[59] ^ t[84];
  assign t[76] = t[69] ^ t[88];
  assign t[77] = t[13] ? t[163] : t[96];
  assign t[78] = t[97] ^ t[98];
  assign t[79] = t[99] & t[100];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[101] ^ t[90];
  assign t[81] = t[65] ^ t[77];
  assign t[82] = t[102] ^ t[103];
  assign t[83] = t[77] ^ t[80];
  assign t[84] = t[104] ^ t[105];
  assign t[85] = t[106] ^ t[107];
  assign t[86] = t[164] ^ t[165];
  assign t[87] = t[166] ^ t[146];
  assign t[88] = t[108] ^ t[91];
  assign t[89] = t[13] ? t[167] : t[109];
  assign t[8] = ~(t[13]);
  assign t[90] = t[13] ? t[168] : t[110];
  assign t[91] = t[13] ? t[169] : t[111];
  assign t[92] = t[112] ^ t[113];
  assign t[93] = t[114] ^ t[115];
  assign t[94] = t[78] ^ t[116];
  assign t[95] = t[117] ^ t[73];
  assign t[96] = t[170] ^ t[171];
  assign t[97] = t[118] ^ t[93];
  assign t[98] = t[56] ^ t[119];
  assign t[99] = t[73] ^ t[116];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [120:0] x;
 output y;

 wire [423:0] t;
  assign t[0] = t[1] ? t[2] : t[144];
  assign t[100] = t[120] ^ t[78];
  assign t[101] = t[13] ? t[172] : t[121];
  assign t[102] = t[95] & t[122];
  assign t[103] = t[95] ^ t[116];
  assign t[104] = t[100] & t[123];
  assign t[105] = t[100] ^ t[116];
  assign t[106] = t[89] ^ t[66];
  assign t[107] = t[80] ^ t[124];
  assign t[108] = t[13] ? t[173] : t[125];
  assign t[109] = t[174] ^ t[175];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[176] ^ t[177];
  assign t[111] = t[178] ^ t[179];
  assign t[112] = t[126] ^ t[127];
  assign t[113] = t[106] ^ t[71];
  assign t[114] = t[106] & t[71];
  assign t[115] = t[69] & t[128];
  assign t[116] = t[120] & t[117];
  assign t[117] = t[129] ^ t[130];
  assign t[118] = t[131] ^ t[132];
  assign t[119] = t[83] ^ t[68];
  assign t[11] = ~(t[17]);
  assign t[120] = t[133] ^ t[130];
  assign t[121] = t[180] ^ t[181];
  assign t[122] = t[117] & t[78];
  assign t[123] = t[73] & t[120];
  assign t[124] = t[91] ^ t[77];
  assign t[125] = t[182] ^ t[183];
  assign t[126] = t[60] & t[77];
  assign t[127] = t[134] & t[76];
  assign t[128] = t[88] ^ t[135];
  assign t[129] = t[136] ^ t[137];
  assign t[12] = t[147] & t[18];
  assign t[130] = t[138] ^ t[115];
  assign t[131] = t[56] & t[119];
  assign t[132] = t[72] & t[68];
  assign t[133] = t[139] ^ t[140];
  assign t[134] = t[72] ^ t[49];
  assign t[135] = t[101] ^ t[66];
  assign t[136] = t[141] ^ t[127];
  assign t[137] = t[85] & t[142];
  assign t[138] = t[49] & t[52];
  assign t[139] = t[143] ^ t[132];
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = t[107] & t[83];
  assign t[141] = t[76] ^ t[135];
  assign t[142] = t[77] ^ t[76];
  assign t[143] = t[72] ^ t[68];
  assign t[144] = (t[184]);
  assign t[145] = (t[185]);
  assign t[146] = (t[186]);
  assign t[147] = (t[187]);
  assign t[148] = (t[188]);
  assign t[149] = (t[189]);
  assign t[14] = ~(t[147]);
  assign t[150] = (t[190]);
  assign t[151] = (t[191]);
  assign t[152] = (t[192]);
  assign t[153] = (t[193]);
  assign t[154] = (t[194]);
  assign t[155] = (t[195]);
  assign t[156] = (t[196]);
  assign t[157] = (t[197]);
  assign t[158] = (t[198]);
  assign t[159] = (t[199]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[200]);
  assign t[161] = (t[201]);
  assign t[162] = (t[202]);
  assign t[163] = (t[203]);
  assign t[164] = (t[204]);
  assign t[165] = (t[205]);
  assign t[166] = (t[206]);
  assign t[167] = (t[207]);
  assign t[168] = (t[208]);
  assign t[169] = (t[209]);
  assign t[16] = t[23] ^ t[24];
  assign t[170] = (t[210]);
  assign t[171] = (t[211]);
  assign t[172] = (t[212]);
  assign t[173] = (t[213]);
  assign t[174] = (t[214]);
  assign t[175] = (t[215]);
  assign t[176] = (t[216]);
  assign t[177] = (t[217]);
  assign t[178] = (t[218]);
  assign t[179] = (t[219]);
  assign t[17] = ~(t[147] & t[25]);
  assign t[180] = (t[220]);
  assign t[181] = (t[221]);
  assign t[182] = (t[222]);
  assign t[183] = (t[223]);
  assign t[184] = t[224] ^ x[2];
  assign t[185] = t[225] ^ x[6];
  assign t[186] = t[226] ^ x[9];
  assign t[187] = t[227] ^ x[12];
  assign t[188] = t[228] ^ x[15];
  assign t[189] = t[229] ^ x[18];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[230] ^ x[21];
  assign t[191] = t[231] ^ x[24];
  assign t[192] = t[232] ^ x[27];
  assign t[193] = t[233] ^ x[30];
  assign t[194] = t[234] ^ x[33];
  assign t[195] = t[235] ^ x[36];
  assign t[196] = t[236] ^ x[39];
  assign t[197] = t[237] ^ x[42];
  assign t[198] = t[238] ^ x[45];
  assign t[199] = t[239] ^ x[48];
  assign t[19] = ~(t[148]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[51];
  assign t[201] = t[241] ^ x[54];
  assign t[202] = t[242] ^ x[57];
  assign t[203] = t[243] ^ x[60];
  assign t[204] = t[244] ^ x[63];
  assign t[205] = t[245] ^ x[66];
  assign t[206] = t[246] ^ x[69];
  assign t[207] = t[247] ^ x[72];
  assign t[208] = t[248] ^ x[75];
  assign t[209] = t[249] ^ x[78];
  assign t[20] = ~(t[147]);
  assign t[210] = t[250] ^ x[81];
  assign t[211] = t[251] ^ x[84];
  assign t[212] = t[252] ^ x[87];
  assign t[213] = t[253] ^ x[90];
  assign t[214] = t[254] ^ x[93];
  assign t[215] = t[255] ^ x[96];
  assign t[216] = t[256] ^ x[99];
  assign t[217] = t[257] ^ x[102];
  assign t[218] = t[258] ^ x[105];
  assign t[219] = t[259] ^ x[108];
  assign t[21] = ~(t[149]);
  assign t[220] = t[260] ^ x[111];
  assign t[221] = t[261] ^ x[114];
  assign t[222] = t[262] ^ x[117];
  assign t[223] = t[263] ^ x[120];
  assign t[224] = (t[264] & ~t[265]);
  assign t[225] = (t[266] & ~t[267]);
  assign t[226] = (t[268] & ~t[269]);
  assign t[227] = (t[270] & ~t[271]);
  assign t[228] = (t[272] & ~t[273]);
  assign t[229] = (t[274] & ~t[275]);
  assign t[22] = ~(t[150]);
  assign t[230] = (t[276] & ~t[277]);
  assign t[231] = (t[278] & ~t[279]);
  assign t[232] = (t[280] & ~t[281]);
  assign t[233] = (t[282] & ~t[283]);
  assign t[234] = (t[284] & ~t[285]);
  assign t[235] = (t[286] & ~t[287]);
  assign t[236] = (t[288] & ~t[289]);
  assign t[237] = (t[290] & ~t[291]);
  assign t[238] = (t[292] & ~t[293]);
  assign t[239] = (t[294] & ~t[295]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[296] & ~t[297]);
  assign t[241] = (t[298] & ~t[299]);
  assign t[242] = (t[300] & ~t[301]);
  assign t[243] = (t[302] & ~t[303]);
  assign t[244] = (t[304] & ~t[305]);
  assign t[245] = (t[306] & ~t[307]);
  assign t[246] = (t[308] & ~t[309]);
  assign t[247] = (t[310] & ~t[311]);
  assign t[248] = (t[312] & ~t[313]);
  assign t[249] = (t[314] & ~t[315]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[316] & ~t[317]);
  assign t[251] = (t[318] & ~t[319]);
  assign t[252] = (t[320] & ~t[321]);
  assign t[253] = (t[322] & ~t[323]);
  assign t[254] = (t[324] & ~t[325]);
  assign t[255] = (t[326] & ~t[327]);
  assign t[256] = (t[328] & ~t[329]);
  assign t[257] = (t[330] & ~t[331]);
  assign t[258] = (t[332] & ~t[333]);
  assign t[259] = (t[334] & ~t[335]);
  assign t[25] = ~(t[151] | t[32]);
  assign t[260] = (t[336] & ~t[337]);
  assign t[261] = (t[338] & ~t[339]);
  assign t[262] = (t[340] & ~t[341]);
  assign t[263] = (t[342] & ~t[343]);
  assign t[264] = t[344] ^ x[2];
  assign t[265] = t[345] ^ x[1];
  assign t[266] = t[346] ^ x[6];
  assign t[267] = t[347] ^ x[5];
  assign t[268] = t[348] ^ x[9];
  assign t[269] = t[349] ^ x[8];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[350] ^ x[12];
  assign t[271] = t[351] ^ x[11];
  assign t[272] = t[352] ^ x[15];
  assign t[273] = t[353] ^ x[14];
  assign t[274] = t[354] ^ x[18];
  assign t[275] = t[355] ^ x[17];
  assign t[276] = t[356] ^ x[21];
  assign t[277] = t[357] ^ x[20];
  assign t[278] = t[358] ^ x[24];
  assign t[279] = t[359] ^ x[23];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[360] ^ x[27];
  assign t[281] = t[361] ^ x[26];
  assign t[282] = t[362] ^ x[30];
  assign t[283] = t[363] ^ x[29];
  assign t[284] = t[364] ^ x[33];
  assign t[285] = t[365] ^ x[32];
  assign t[286] = t[366] ^ x[36];
  assign t[287] = t[367] ^ x[35];
  assign t[288] = t[368] ^ x[39];
  assign t[289] = t[369] ^ x[38];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[370] ^ x[42];
  assign t[291] = t[371] ^ x[41];
  assign t[292] = t[372] ^ x[45];
  assign t[293] = t[373] ^ x[44];
  assign t[294] = t[374] ^ x[48];
  assign t[295] = t[375] ^ x[47];
  assign t[296] = t[376] ^ x[51];
  assign t[297] = t[377] ^ x[50];
  assign t[298] = t[378] ^ x[54];
  assign t[299] = t[379] ^ x[53];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[380] ^ x[57];
  assign t[301] = t[381] ^ x[56];
  assign t[302] = t[382] ^ x[60];
  assign t[303] = t[383] ^ x[59];
  assign t[304] = t[384] ^ x[63];
  assign t[305] = t[385] ^ x[62];
  assign t[306] = t[386] ^ x[66];
  assign t[307] = t[387] ^ x[65];
  assign t[308] = t[388] ^ x[69];
  assign t[309] = t[389] ^ x[68];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[390] ^ x[72];
  assign t[311] = t[391] ^ x[71];
  assign t[312] = t[392] ^ x[75];
  assign t[313] = t[393] ^ x[74];
  assign t[314] = t[394] ^ x[78];
  assign t[315] = t[395] ^ x[77];
  assign t[316] = t[396] ^ x[81];
  assign t[317] = t[397] ^ x[80];
  assign t[318] = t[398] ^ x[84];
  assign t[319] = t[399] ^ x[83];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[400] ^ x[87];
  assign t[321] = t[401] ^ x[86];
  assign t[322] = t[402] ^ x[90];
  assign t[323] = t[403] ^ x[89];
  assign t[324] = t[404] ^ x[93];
  assign t[325] = t[405] ^ x[92];
  assign t[326] = t[406] ^ x[96];
  assign t[327] = t[407] ^ x[95];
  assign t[328] = t[408] ^ x[99];
  assign t[329] = t[409] ^ x[98];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[410] ^ x[102];
  assign t[331] = t[411] ^ x[101];
  assign t[332] = t[412] ^ x[105];
  assign t[333] = t[413] ^ x[104];
  assign t[334] = t[414] ^ x[108];
  assign t[335] = t[415] ^ x[107];
  assign t[336] = t[416] ^ x[111];
  assign t[337] = t[417] ^ x[110];
  assign t[338] = t[418] ^ x[114];
  assign t[339] = t[419] ^ x[113];
  assign t[33] = ~(t[152] & t[153]);
  assign t[340] = t[420] ^ x[117];
  assign t[341] = t[421] ^ x[116];
  assign t[342] = t[422] ^ x[120];
  assign t[343] = t[423] ^ x[119];
  assign t[344] = (x[0]);
  assign t[345] = (x[0]);
  assign t[346] = (x[4]);
  assign t[347] = (x[4]);
  assign t[348] = (x[7]);
  assign t[349] = (x[7]);
  assign t[34] = ~(t[154] & t[149]);
  assign t[350] = (x[10]);
  assign t[351] = (x[10]);
  assign t[352] = (x[13]);
  assign t[353] = (x[13]);
  assign t[354] = (x[16]);
  assign t[355] = (x[16]);
  assign t[356] = (x[19]);
  assign t[357] = (x[19]);
  assign t[358] = (x[22]);
  assign t[359] = (x[22]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[25]);
  assign t[361] = (x[25]);
  assign t[362] = (x[28]);
  assign t[363] = (x[28]);
  assign t[364] = (x[31]);
  assign t[365] = (x[31]);
  assign t[366] = (x[34]);
  assign t[367] = (x[34]);
  assign t[368] = (x[37]);
  assign t[369] = (x[37]);
  assign t[36] = ~(t[155] & t[47]);
  assign t[370] = (x[40]);
  assign t[371] = (x[40]);
  assign t[372] = (x[43]);
  assign t[373] = (x[43]);
  assign t[374] = (x[46]);
  assign t[375] = (x[46]);
  assign t[376] = (x[49]);
  assign t[377] = (x[49]);
  assign t[378] = (x[52]);
  assign t[379] = (x[52]);
  assign t[37] = t[48] & t[49];
  assign t[380] = (x[55]);
  assign t[381] = (x[55]);
  assign t[382] = (x[58]);
  assign t[383] = (x[58]);
  assign t[384] = (x[61]);
  assign t[385] = (x[61]);
  assign t[386] = (x[64]);
  assign t[387] = (x[64]);
  assign t[388] = (x[67]);
  assign t[389] = (x[67]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[70]);
  assign t[391] = (x[70]);
  assign t[392] = (x[73]);
  assign t[393] = (x[73]);
  assign t[394] = (x[76]);
  assign t[395] = (x[76]);
  assign t[396] = (x[79]);
  assign t[397] = (x[79]);
  assign t[398] = (x[82]);
  assign t[399] = (x[82]);
  assign t[39] = t[48] & t[52];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[85]);
  assign t[401] = (x[85]);
  assign t[402] = (x[88]);
  assign t[403] = (x[88]);
  assign t[404] = (x[91]);
  assign t[405] = (x[91]);
  assign t[406] = (x[94]);
  assign t[407] = (x[94]);
  assign t[408] = (x[97]);
  assign t[409] = (x[97]);
  assign t[40] = t[53] ^ t[54];
  assign t[410] = (x[100]);
  assign t[411] = (x[100]);
  assign t[412] = (x[103]);
  assign t[413] = (x[103]);
  assign t[414] = (x[106]);
  assign t[415] = (x[106]);
  assign t[416] = (x[109]);
  assign t[417] = (x[109]);
  assign t[418] = (x[112]);
  assign t[419] = (x[112]);
  assign t[41] = t[55] & t[56];
  assign t[420] = (x[115]);
  assign t[421] = (x[115]);
  assign t[422] = (x[118]);
  assign t[423] = (x[118]);
  assign t[42] = t[57] ^ t[58];
  assign t[43] = t[59] & t[60];
  assign t[44] = t[61] ^ t[62];
  assign t[45] = ~(t[156] | t[157]);
  assign t[46] = ~(t[158] | t[159]);
  assign t[47] = ~(t[160]);
  assign t[48] = t[63] ^ t[64];
  assign t[49] = t[65] ^ t[66];
  assign t[4] = ~(t[8]);
  assign t[50] = t[67] & t[68];
  assign t[51] = t[63] & t[69];
  assign t[52] = t[69] ^ t[70];
  assign t[53] = t[64] & t[71];
  assign t[54] = t[67] & t[72];
  assign t[55] = t[73] ^ t[74];
  assign t[56] = t[69] ^ t[60];
  assign t[57] = t[75] & t[76];
  assign t[58] = t[59] & t[77];
  assign t[59] = t[78] ^ t[79];
  assign t[5] = t[9] ? t[145] : x[3];
  assign t[60] = t[80] ^ t[81];
  assign t[61] = t[82] & t[83];
  assign t[62] = t[84] & t[85];
  assign t[63] = t[55] ^ t[59];
  assign t[64] = t[82] ^ t[84];
  assign t[65] = t[13] ? t[161] : t[86];
  assign t[66] = t[13] ? t[162] : t[87];
  assign t[67] = t[55] ^ t[82];
  assign t[68] = t[88] ^ t[70];
  assign t[69] = t[89] ^ t[65];
  assign t[6] = ~(t[10] ^ t[146]);
  assign t[70] = t[90] ^ t[66];
  assign t[71] = t[76] ^ t[80];
  assign t[72] = t[89] ^ t[91];
  assign t[73] = t[92] ^ t[93];
  assign t[74] = t[94] & t[95];
  assign t[75] = t[59] ^ t[84];
  assign t[76] = t[69] ^ t[88];
  assign t[77] = t[13] ? t[163] : t[96];
  assign t[78] = t[97] ^ t[98];
  assign t[79] = t[99] & t[100];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[101] ^ t[90];
  assign t[81] = t[65] ^ t[77];
  assign t[82] = t[102] ^ t[103];
  assign t[83] = t[77] ^ t[80];
  assign t[84] = t[104] ^ t[105];
  assign t[85] = t[106] ^ t[107];
  assign t[86] = t[164] ^ t[165];
  assign t[87] = t[166] ^ t[146];
  assign t[88] = t[108] ^ t[91];
  assign t[89] = t[13] ? t[167] : t[109];
  assign t[8] = ~(t[13]);
  assign t[90] = t[13] ? t[168] : t[110];
  assign t[91] = t[13] ? t[169] : t[111];
  assign t[92] = t[112] ^ t[113];
  assign t[93] = t[114] ^ t[115];
  assign t[94] = t[78] ^ t[116];
  assign t[95] = t[117] ^ t[73];
  assign t[96] = t[170] ^ t[171];
  assign t[97] = t[118] ^ t[93];
  assign t[98] = t[56] ^ t[119];
  assign t[99] = t[73] ^ t[116];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [123:0] x;
 output y;

 wire [421:0] t;
  assign t[0] = t[1] ? t[2] : t[135];
  assign t[100] = t[76] ^ t[87];
  assign t[101] = t[89] ^ t[66];
  assign t[102] = t[114] ^ t[115];
  assign t[103] = t[116] ^ t[115];
  assign t[104] = t[168] ^ t[169];
  assign t[105] = t[170] ^ t[171];
  assign t[106] = t[13] ? t[172] : t[117];
  assign t[107] = t[173] ^ t[174];
  assign t[108] = t[118] ^ t[119];
  assign t[109] = t[49] ^ t[120];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[121] ^ t[122];
  assign t[111] = t[72] ^ t[123];
  assign t[112] = t[72] & t[123];
  assign t[113] = t[49] & t[124];
  assign t[114] = t[125] ^ t[126];
  assign t[115] = t[127] ^ t[113];
  assign t[116] = t[128] ^ t[129];
  assign t[117] = t[175] ^ t[137];
  assign t[118] = t[109] & t[62];
  assign t[119] = t[75] & t[81];
  assign t[11] = ~(t[17]);
  assign t[120] = t[69] ^ t[130];
  assign t[121] = t[120] & t[60];
  assign t[122] = t[58] & t[74];
  assign t[123] = t[74] ^ t[69];
  assign t[124] = t[93] ^ t[131];
  assign t[125] = t[132] ^ t[122];
  assign t[126] = t[55] & t[56];
  assign t[127] = t[51] & t[133];
  assign t[128] = t[134] ^ t[119];
  assign t[129] = t[73] & t[53];
  assign t[12] = t[138] & t[18];
  assign t[130] = t[64] ^ t[60];
  assign t[131] = t[88] ^ t[66];
  assign t[132] = t[74] ^ t[131];
  assign t[133] = t[49] ^ t[101];
  assign t[134] = t[75] ^ t[81];
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = ~(t[138]);
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = (t[194]);
  assign t[154] = (t[195]);
  assign t[155] = (t[196]);
  assign t[156] = (t[197]);
  assign t[157] = (t[198]);
  assign t[158] = (t[199]);
  assign t[159] = (t[200]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[201]);
  assign t[161] = (t[202]);
  assign t[162] = (t[203]);
  assign t[163] = (t[204]);
  assign t[164] = (t[205]);
  assign t[165] = (t[206]);
  assign t[166] = (t[207]);
  assign t[167] = (t[208]);
  assign t[168] = (t[209]);
  assign t[169] = (t[210]);
  assign t[16] = t[23] ^ t[24];
  assign t[170] = (t[211]);
  assign t[171] = (t[212]);
  assign t[172] = (t[213]);
  assign t[173] = (t[214]);
  assign t[174] = (t[215]);
  assign t[175] = (t[216]);
  assign t[176] = t[217] ^ x[2];
  assign t[177] = t[218] ^ x[6];
  assign t[178] = t[219] ^ x[9];
  assign t[179] = t[220] ^ x[12];
  assign t[17] = ~(t[138] & t[25]);
  assign t[180] = t[221] ^ x[15];
  assign t[181] = t[222] ^ x[18];
  assign t[182] = t[223] ^ x[21];
  assign t[183] = t[224] ^ x[24];
  assign t[184] = t[225] ^ x[27];
  assign t[185] = t[226] ^ x[30];
  assign t[186] = t[227] ^ x[33];
  assign t[187] = t[228] ^ x[36];
  assign t[188] = t[229] ^ x[39];
  assign t[189] = t[230] ^ x[42];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[231] ^ x[45];
  assign t[191] = t[232] ^ x[48];
  assign t[192] = t[233] ^ x[51];
  assign t[193] = t[234] ^ x[54];
  assign t[194] = t[235] ^ x[57];
  assign t[195] = t[236] ^ x[60];
  assign t[196] = t[237] ^ x[63];
  assign t[197] = t[238] ^ x[66];
  assign t[198] = t[239] ^ x[69];
  assign t[199] = t[240] ^ x[72];
  assign t[19] = ~(t[139]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[241] ^ x[75];
  assign t[201] = t[242] ^ x[78];
  assign t[202] = t[243] ^ x[81];
  assign t[203] = t[244] ^ x[84];
  assign t[204] = t[245] ^ x[87];
  assign t[205] = t[246] ^ x[90];
  assign t[206] = t[247] ^ x[93];
  assign t[207] = t[248] ^ x[96];
  assign t[208] = t[249] ^ x[99];
  assign t[209] = t[250] ^ x[102];
  assign t[20] = ~(t[138]);
  assign t[210] = t[251] ^ x[105];
  assign t[211] = t[252] ^ x[108];
  assign t[212] = t[253] ^ x[111];
  assign t[213] = t[254] ^ x[114];
  assign t[214] = t[255] ^ x[117];
  assign t[215] = t[256] ^ x[120];
  assign t[216] = t[257] ^ x[123];
  assign t[217] = (t[258] & ~t[259]);
  assign t[218] = (t[260] & ~t[261]);
  assign t[219] = (t[262] & ~t[263]);
  assign t[21] = ~(t[140]);
  assign t[220] = (t[264] & ~t[265]);
  assign t[221] = (t[266] & ~t[267]);
  assign t[222] = (t[268] & ~t[269]);
  assign t[223] = (t[270] & ~t[271]);
  assign t[224] = (t[272] & ~t[273]);
  assign t[225] = (t[274] & ~t[275]);
  assign t[226] = (t[276] & ~t[277]);
  assign t[227] = (t[278] & ~t[279]);
  assign t[228] = (t[280] & ~t[281]);
  assign t[229] = (t[282] & ~t[283]);
  assign t[22] = ~(t[141]);
  assign t[230] = (t[284] & ~t[285]);
  assign t[231] = (t[286] & ~t[287]);
  assign t[232] = (t[288] & ~t[289]);
  assign t[233] = (t[290] & ~t[291]);
  assign t[234] = (t[292] & ~t[293]);
  assign t[235] = (t[294] & ~t[295]);
  assign t[236] = (t[296] & ~t[297]);
  assign t[237] = (t[298] & ~t[299]);
  assign t[238] = (t[300] & ~t[301]);
  assign t[239] = (t[302] & ~t[303]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[304] & ~t[305]);
  assign t[241] = (t[306] & ~t[307]);
  assign t[242] = (t[308] & ~t[309]);
  assign t[243] = (t[310] & ~t[311]);
  assign t[244] = (t[312] & ~t[313]);
  assign t[245] = (t[314] & ~t[315]);
  assign t[246] = (t[316] & ~t[317]);
  assign t[247] = (t[318] & ~t[319]);
  assign t[248] = (t[320] & ~t[321]);
  assign t[249] = (t[322] & ~t[323]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[324] & ~t[325]);
  assign t[251] = (t[326] & ~t[327]);
  assign t[252] = (t[328] & ~t[329]);
  assign t[253] = (t[330] & ~t[331]);
  assign t[254] = (t[332] & ~t[333]);
  assign t[255] = (t[334] & ~t[335]);
  assign t[256] = (t[336] & ~t[337]);
  assign t[257] = (t[338] & ~t[339]);
  assign t[258] = t[340] ^ x[2];
  assign t[259] = t[341] ^ x[1];
  assign t[25] = ~(t[142] | t[32]);
  assign t[260] = t[342] ^ x[6];
  assign t[261] = t[343] ^ x[5];
  assign t[262] = t[344] ^ x[9];
  assign t[263] = t[345] ^ x[8];
  assign t[264] = t[346] ^ x[12];
  assign t[265] = t[347] ^ x[11];
  assign t[266] = t[348] ^ x[15];
  assign t[267] = t[349] ^ x[14];
  assign t[268] = t[350] ^ x[18];
  assign t[269] = t[351] ^ x[17];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[352] ^ x[21];
  assign t[271] = t[353] ^ x[20];
  assign t[272] = t[354] ^ x[24];
  assign t[273] = t[355] ^ x[23];
  assign t[274] = t[356] ^ x[27];
  assign t[275] = t[357] ^ x[26];
  assign t[276] = t[358] ^ x[30];
  assign t[277] = t[359] ^ x[29];
  assign t[278] = t[360] ^ x[33];
  assign t[279] = t[361] ^ x[32];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[362] ^ x[36];
  assign t[281] = t[363] ^ x[35];
  assign t[282] = t[364] ^ x[39];
  assign t[283] = t[365] ^ x[38];
  assign t[284] = t[366] ^ x[42];
  assign t[285] = t[367] ^ x[41];
  assign t[286] = t[368] ^ x[45];
  assign t[287] = t[369] ^ x[44];
  assign t[288] = t[370] ^ x[48];
  assign t[289] = t[371] ^ x[47];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[372] ^ x[51];
  assign t[291] = t[373] ^ x[50];
  assign t[292] = t[374] ^ x[54];
  assign t[293] = t[375] ^ x[53];
  assign t[294] = t[376] ^ x[57];
  assign t[295] = t[377] ^ x[56];
  assign t[296] = t[378] ^ x[60];
  assign t[297] = t[379] ^ x[59];
  assign t[298] = t[380] ^ x[63];
  assign t[299] = t[381] ^ x[62];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[66];
  assign t[301] = t[383] ^ x[65];
  assign t[302] = t[384] ^ x[69];
  assign t[303] = t[385] ^ x[68];
  assign t[304] = t[386] ^ x[72];
  assign t[305] = t[387] ^ x[71];
  assign t[306] = t[388] ^ x[75];
  assign t[307] = t[389] ^ x[74];
  assign t[308] = t[390] ^ x[78];
  assign t[309] = t[391] ^ x[77];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[392] ^ x[81];
  assign t[311] = t[393] ^ x[80];
  assign t[312] = t[394] ^ x[84];
  assign t[313] = t[395] ^ x[83];
  assign t[314] = t[396] ^ x[87];
  assign t[315] = t[397] ^ x[86];
  assign t[316] = t[398] ^ x[90];
  assign t[317] = t[399] ^ x[89];
  assign t[318] = t[400] ^ x[93];
  assign t[319] = t[401] ^ x[92];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[402] ^ x[96];
  assign t[321] = t[403] ^ x[95];
  assign t[322] = t[404] ^ x[99];
  assign t[323] = t[405] ^ x[98];
  assign t[324] = t[406] ^ x[102];
  assign t[325] = t[407] ^ x[101];
  assign t[326] = t[408] ^ x[105];
  assign t[327] = t[409] ^ x[104];
  assign t[328] = t[410] ^ x[108];
  assign t[329] = t[411] ^ x[107];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[412] ^ x[111];
  assign t[331] = t[413] ^ x[110];
  assign t[332] = t[414] ^ x[114];
  assign t[333] = t[415] ^ x[113];
  assign t[334] = t[416] ^ x[117];
  assign t[335] = t[417] ^ x[116];
  assign t[336] = t[418] ^ x[120];
  assign t[337] = t[419] ^ x[119];
  assign t[338] = t[420] ^ x[123];
  assign t[339] = t[421] ^ x[122];
  assign t[33] = ~(t[143] & t[144]);
  assign t[340] = (x[0]);
  assign t[341] = (x[0]);
  assign t[342] = (x[4]);
  assign t[343] = (x[4]);
  assign t[344] = (x[7]);
  assign t[345] = (x[7]);
  assign t[346] = (x[10]);
  assign t[347] = (x[10]);
  assign t[348] = (x[13]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[145] & t[146]);
  assign t[350] = (x[16]);
  assign t[351] = (x[16]);
  assign t[352] = (x[19]);
  assign t[353] = (x[19]);
  assign t[354] = (x[22]);
  assign t[355] = (x[22]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[28]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[31]);
  assign t[361] = (x[31]);
  assign t[362] = (x[34]);
  assign t[363] = (x[34]);
  assign t[364] = (x[37]);
  assign t[365] = (x[37]);
  assign t[366] = (x[40]);
  assign t[367] = (x[40]);
  assign t[368] = (x[43]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[147] & t[47]);
  assign t[370] = (x[46]);
  assign t[371] = (x[46]);
  assign t[372] = (x[49]);
  assign t[373] = (x[49]);
  assign t[374] = (x[52]);
  assign t[375] = (x[52]);
  assign t[376] = (x[55]);
  assign t[377] = (x[55]);
  assign t[378] = (x[58]);
  assign t[379] = (x[58]);
  assign t[37] = t[48] & t[49];
  assign t[380] = (x[61]);
  assign t[381] = (x[61]);
  assign t[382] = (x[64]);
  assign t[383] = (x[64]);
  assign t[384] = (x[67]);
  assign t[385] = (x[67]);
  assign t[386] = (x[70]);
  assign t[387] = (x[70]);
  assign t[388] = (x[73]);
  assign t[389] = (x[73]);
  assign t[38] = t[50] & t[51];
  assign t[390] = (x[76]);
  assign t[391] = (x[76]);
  assign t[392] = (x[79]);
  assign t[393] = (x[79]);
  assign t[394] = (x[82]);
  assign t[395] = (x[82]);
  assign t[396] = (x[85]);
  assign t[397] = (x[85]);
  assign t[398] = (x[88]);
  assign t[399] = (x[88]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[91]);
  assign t[401] = (x[91]);
  assign t[402] = (x[94]);
  assign t[403] = (x[94]);
  assign t[404] = (x[97]);
  assign t[405] = (x[97]);
  assign t[406] = (x[100]);
  assign t[407] = (x[100]);
  assign t[408] = (x[103]);
  assign t[409] = (x[103]);
  assign t[40] = t[54] & t[55];
  assign t[410] = (x[106]);
  assign t[411] = (x[106]);
  assign t[412] = (x[109]);
  assign t[413] = (x[109]);
  assign t[414] = (x[112]);
  assign t[415] = (x[112]);
  assign t[416] = (x[115]);
  assign t[417] = (x[115]);
  assign t[418] = (x[118]);
  assign t[419] = (x[118]);
  assign t[41] = t[54] & t[56];
  assign t[420] = (x[121]);
  assign t[421] = (x[121]);
  assign t[42] = t[57] & t[58];
  assign t[43] = t[59] & t[60];
  assign t[44] = t[61] & t[62];
  assign t[45] = ~(t[148] | t[149]);
  assign t[46] = ~(t[150] | t[151]);
  assign t[47] = ~(t[152]);
  assign t[48] = t[61] ^ t[59];
  assign t[49] = t[63] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[48] ^ t[65];
  assign t[51] = t[64] ^ t[66];
  assign t[52] = t[67] ^ t[68];
  assign t[53] = t[60] ^ t[69];
  assign t[54] = t[70] ^ t[71];
  assign t[55] = t[72] ^ t[73];
  assign t[56] = t[60] ^ t[74];
  assign t[57] = t[59] ^ t[54];
  assign t[58] = t[75] ^ t[51];
  assign t[59] = t[76] ^ t[77];
  assign t[5] = t[9] ? t[136] : x[3];
  assign t[60] = t[13] ? t[153] : t[78];
  assign t[61] = t[79] ^ t[80];
  assign t[62] = t[53] ^ t[81];
  assign t[63] = t[13] ? t[154] : t[82];
  assign t[64] = t[13] ? t[155] : t[83];
  assign t[65] = t[52] ^ t[54];
  assign t[66] = t[13] ? t[156] : t[84];
  assign t[67] = t[85] & t[86];
  assign t[68] = t[85] ^ t[87];
  assign t[69] = t[88] ^ t[89];
  assign t[6] = ~(t[10] ^ t[137]);
  assign t[70] = t[90] & t[91];
  assign t[71] = t[90] ^ t[87];
  assign t[72] = t[63] ^ t[66];
  assign t[73] = t[69] ^ t[92];
  assign t[74] = t[49] ^ t[93];
  assign t[75] = t[63] ^ t[94];
  assign t[76] = t[95] ^ t[96];
  assign t[77] = t[97] & t[90];
  assign t[78] = t[157] ^ t[158];
  assign t[79] = t[98] ^ t[99];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[100] & t[85];
  assign t[81] = t[93] ^ t[101];
  assign t[82] = t[159] ^ t[160];
  assign t[83] = t[161] ^ t[162];
  assign t[84] = t[163] ^ t[164];
  assign t[85] = t[102] ^ t[79];
  assign t[86] = t[102] & t[76];
  assign t[87] = t[103] & t[102];
  assign t[88] = t[13] ? t[165] : t[104];
  assign t[89] = t[13] ? t[166] : t[105];
  assign t[8] = ~(t[13]);
  assign t[90] = t[103] ^ t[76];
  assign t[91] = t[79] & t[103];
  assign t[92] = t[94] ^ t[60];
  assign t[93] = t[106] ^ t[94];
  assign t[94] = t[13] ? t[167] : t[107];
  assign t[95] = t[108] ^ t[99];
  assign t[96] = t[109] ^ t[62];
  assign t[97] = t[79] ^ t[87];
  assign t[98] = t[110] ^ t[111];
  assign t[99] = t[112] ^ t[113];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [123:0] x;
 output y;

 wire [421:0] t;
  assign t[0] = t[1] ? t[2] : t[135];
  assign t[100] = t[76] ^ t[87];
  assign t[101] = t[89] ^ t[66];
  assign t[102] = t[114] ^ t[115];
  assign t[103] = t[116] ^ t[115];
  assign t[104] = t[168] ^ t[169];
  assign t[105] = t[170] ^ t[171];
  assign t[106] = t[13] ? t[172] : t[117];
  assign t[107] = t[173] ^ t[174];
  assign t[108] = t[118] ^ t[119];
  assign t[109] = t[49] ^ t[120];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[121] ^ t[122];
  assign t[111] = t[72] ^ t[123];
  assign t[112] = t[72] & t[123];
  assign t[113] = t[49] & t[124];
  assign t[114] = t[125] ^ t[126];
  assign t[115] = t[127] ^ t[113];
  assign t[116] = t[128] ^ t[129];
  assign t[117] = t[175] ^ t[137];
  assign t[118] = t[109] & t[62];
  assign t[119] = t[75] & t[81];
  assign t[11] = ~(t[17]);
  assign t[120] = t[69] ^ t[130];
  assign t[121] = t[120] & t[60];
  assign t[122] = t[58] & t[74];
  assign t[123] = t[74] ^ t[69];
  assign t[124] = t[93] ^ t[131];
  assign t[125] = t[132] ^ t[122];
  assign t[126] = t[55] & t[56];
  assign t[127] = t[51] & t[133];
  assign t[128] = t[134] ^ t[119];
  assign t[129] = t[73] & t[53];
  assign t[12] = t[138] & t[18];
  assign t[130] = t[64] ^ t[60];
  assign t[131] = t[88] ^ t[66];
  assign t[132] = t[74] ^ t[131];
  assign t[133] = t[49] ^ t[101];
  assign t[134] = t[75] ^ t[81];
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = ~(t[138]);
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = (t[194]);
  assign t[154] = (t[195]);
  assign t[155] = (t[196]);
  assign t[156] = (t[197]);
  assign t[157] = (t[198]);
  assign t[158] = (t[199]);
  assign t[159] = (t[200]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[201]);
  assign t[161] = (t[202]);
  assign t[162] = (t[203]);
  assign t[163] = (t[204]);
  assign t[164] = (t[205]);
  assign t[165] = (t[206]);
  assign t[166] = (t[207]);
  assign t[167] = (t[208]);
  assign t[168] = (t[209]);
  assign t[169] = (t[210]);
  assign t[16] = t[23] ^ t[24];
  assign t[170] = (t[211]);
  assign t[171] = (t[212]);
  assign t[172] = (t[213]);
  assign t[173] = (t[214]);
  assign t[174] = (t[215]);
  assign t[175] = (t[216]);
  assign t[176] = t[217] ^ x[2];
  assign t[177] = t[218] ^ x[6];
  assign t[178] = t[219] ^ x[9];
  assign t[179] = t[220] ^ x[12];
  assign t[17] = ~(t[138] & t[25]);
  assign t[180] = t[221] ^ x[15];
  assign t[181] = t[222] ^ x[18];
  assign t[182] = t[223] ^ x[21];
  assign t[183] = t[224] ^ x[24];
  assign t[184] = t[225] ^ x[27];
  assign t[185] = t[226] ^ x[30];
  assign t[186] = t[227] ^ x[33];
  assign t[187] = t[228] ^ x[36];
  assign t[188] = t[229] ^ x[39];
  assign t[189] = t[230] ^ x[42];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[231] ^ x[45];
  assign t[191] = t[232] ^ x[48];
  assign t[192] = t[233] ^ x[51];
  assign t[193] = t[234] ^ x[54];
  assign t[194] = t[235] ^ x[57];
  assign t[195] = t[236] ^ x[60];
  assign t[196] = t[237] ^ x[63];
  assign t[197] = t[238] ^ x[66];
  assign t[198] = t[239] ^ x[69];
  assign t[199] = t[240] ^ x[72];
  assign t[19] = ~(t[139]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[241] ^ x[75];
  assign t[201] = t[242] ^ x[78];
  assign t[202] = t[243] ^ x[81];
  assign t[203] = t[244] ^ x[84];
  assign t[204] = t[245] ^ x[87];
  assign t[205] = t[246] ^ x[90];
  assign t[206] = t[247] ^ x[93];
  assign t[207] = t[248] ^ x[96];
  assign t[208] = t[249] ^ x[99];
  assign t[209] = t[250] ^ x[102];
  assign t[20] = ~(t[138]);
  assign t[210] = t[251] ^ x[105];
  assign t[211] = t[252] ^ x[108];
  assign t[212] = t[253] ^ x[111];
  assign t[213] = t[254] ^ x[114];
  assign t[214] = t[255] ^ x[117];
  assign t[215] = t[256] ^ x[120];
  assign t[216] = t[257] ^ x[123];
  assign t[217] = (t[258] & ~t[259]);
  assign t[218] = (t[260] & ~t[261]);
  assign t[219] = (t[262] & ~t[263]);
  assign t[21] = ~(t[140]);
  assign t[220] = (t[264] & ~t[265]);
  assign t[221] = (t[266] & ~t[267]);
  assign t[222] = (t[268] & ~t[269]);
  assign t[223] = (t[270] & ~t[271]);
  assign t[224] = (t[272] & ~t[273]);
  assign t[225] = (t[274] & ~t[275]);
  assign t[226] = (t[276] & ~t[277]);
  assign t[227] = (t[278] & ~t[279]);
  assign t[228] = (t[280] & ~t[281]);
  assign t[229] = (t[282] & ~t[283]);
  assign t[22] = ~(t[141]);
  assign t[230] = (t[284] & ~t[285]);
  assign t[231] = (t[286] & ~t[287]);
  assign t[232] = (t[288] & ~t[289]);
  assign t[233] = (t[290] & ~t[291]);
  assign t[234] = (t[292] & ~t[293]);
  assign t[235] = (t[294] & ~t[295]);
  assign t[236] = (t[296] & ~t[297]);
  assign t[237] = (t[298] & ~t[299]);
  assign t[238] = (t[300] & ~t[301]);
  assign t[239] = (t[302] & ~t[303]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[304] & ~t[305]);
  assign t[241] = (t[306] & ~t[307]);
  assign t[242] = (t[308] & ~t[309]);
  assign t[243] = (t[310] & ~t[311]);
  assign t[244] = (t[312] & ~t[313]);
  assign t[245] = (t[314] & ~t[315]);
  assign t[246] = (t[316] & ~t[317]);
  assign t[247] = (t[318] & ~t[319]);
  assign t[248] = (t[320] & ~t[321]);
  assign t[249] = (t[322] & ~t[323]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[324] & ~t[325]);
  assign t[251] = (t[326] & ~t[327]);
  assign t[252] = (t[328] & ~t[329]);
  assign t[253] = (t[330] & ~t[331]);
  assign t[254] = (t[332] & ~t[333]);
  assign t[255] = (t[334] & ~t[335]);
  assign t[256] = (t[336] & ~t[337]);
  assign t[257] = (t[338] & ~t[339]);
  assign t[258] = t[340] ^ x[2];
  assign t[259] = t[341] ^ x[1];
  assign t[25] = ~(t[142] | t[32]);
  assign t[260] = t[342] ^ x[6];
  assign t[261] = t[343] ^ x[5];
  assign t[262] = t[344] ^ x[9];
  assign t[263] = t[345] ^ x[8];
  assign t[264] = t[346] ^ x[12];
  assign t[265] = t[347] ^ x[11];
  assign t[266] = t[348] ^ x[15];
  assign t[267] = t[349] ^ x[14];
  assign t[268] = t[350] ^ x[18];
  assign t[269] = t[351] ^ x[17];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[352] ^ x[21];
  assign t[271] = t[353] ^ x[20];
  assign t[272] = t[354] ^ x[24];
  assign t[273] = t[355] ^ x[23];
  assign t[274] = t[356] ^ x[27];
  assign t[275] = t[357] ^ x[26];
  assign t[276] = t[358] ^ x[30];
  assign t[277] = t[359] ^ x[29];
  assign t[278] = t[360] ^ x[33];
  assign t[279] = t[361] ^ x[32];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[362] ^ x[36];
  assign t[281] = t[363] ^ x[35];
  assign t[282] = t[364] ^ x[39];
  assign t[283] = t[365] ^ x[38];
  assign t[284] = t[366] ^ x[42];
  assign t[285] = t[367] ^ x[41];
  assign t[286] = t[368] ^ x[45];
  assign t[287] = t[369] ^ x[44];
  assign t[288] = t[370] ^ x[48];
  assign t[289] = t[371] ^ x[47];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[372] ^ x[51];
  assign t[291] = t[373] ^ x[50];
  assign t[292] = t[374] ^ x[54];
  assign t[293] = t[375] ^ x[53];
  assign t[294] = t[376] ^ x[57];
  assign t[295] = t[377] ^ x[56];
  assign t[296] = t[378] ^ x[60];
  assign t[297] = t[379] ^ x[59];
  assign t[298] = t[380] ^ x[63];
  assign t[299] = t[381] ^ x[62];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[66];
  assign t[301] = t[383] ^ x[65];
  assign t[302] = t[384] ^ x[69];
  assign t[303] = t[385] ^ x[68];
  assign t[304] = t[386] ^ x[72];
  assign t[305] = t[387] ^ x[71];
  assign t[306] = t[388] ^ x[75];
  assign t[307] = t[389] ^ x[74];
  assign t[308] = t[390] ^ x[78];
  assign t[309] = t[391] ^ x[77];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[392] ^ x[81];
  assign t[311] = t[393] ^ x[80];
  assign t[312] = t[394] ^ x[84];
  assign t[313] = t[395] ^ x[83];
  assign t[314] = t[396] ^ x[87];
  assign t[315] = t[397] ^ x[86];
  assign t[316] = t[398] ^ x[90];
  assign t[317] = t[399] ^ x[89];
  assign t[318] = t[400] ^ x[93];
  assign t[319] = t[401] ^ x[92];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[402] ^ x[96];
  assign t[321] = t[403] ^ x[95];
  assign t[322] = t[404] ^ x[99];
  assign t[323] = t[405] ^ x[98];
  assign t[324] = t[406] ^ x[102];
  assign t[325] = t[407] ^ x[101];
  assign t[326] = t[408] ^ x[105];
  assign t[327] = t[409] ^ x[104];
  assign t[328] = t[410] ^ x[108];
  assign t[329] = t[411] ^ x[107];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[412] ^ x[111];
  assign t[331] = t[413] ^ x[110];
  assign t[332] = t[414] ^ x[114];
  assign t[333] = t[415] ^ x[113];
  assign t[334] = t[416] ^ x[117];
  assign t[335] = t[417] ^ x[116];
  assign t[336] = t[418] ^ x[120];
  assign t[337] = t[419] ^ x[119];
  assign t[338] = t[420] ^ x[123];
  assign t[339] = t[421] ^ x[122];
  assign t[33] = ~(t[143] & t[144]);
  assign t[340] = (x[0]);
  assign t[341] = (x[0]);
  assign t[342] = (x[4]);
  assign t[343] = (x[4]);
  assign t[344] = (x[7]);
  assign t[345] = (x[7]);
  assign t[346] = (x[10]);
  assign t[347] = (x[10]);
  assign t[348] = (x[13]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[145] & t[146]);
  assign t[350] = (x[16]);
  assign t[351] = (x[16]);
  assign t[352] = (x[19]);
  assign t[353] = (x[19]);
  assign t[354] = (x[22]);
  assign t[355] = (x[22]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[28]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[31]);
  assign t[361] = (x[31]);
  assign t[362] = (x[34]);
  assign t[363] = (x[34]);
  assign t[364] = (x[37]);
  assign t[365] = (x[37]);
  assign t[366] = (x[40]);
  assign t[367] = (x[40]);
  assign t[368] = (x[43]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[147] & t[47]);
  assign t[370] = (x[46]);
  assign t[371] = (x[46]);
  assign t[372] = (x[49]);
  assign t[373] = (x[49]);
  assign t[374] = (x[52]);
  assign t[375] = (x[52]);
  assign t[376] = (x[55]);
  assign t[377] = (x[55]);
  assign t[378] = (x[58]);
  assign t[379] = (x[58]);
  assign t[37] = t[48] & t[49];
  assign t[380] = (x[61]);
  assign t[381] = (x[61]);
  assign t[382] = (x[64]);
  assign t[383] = (x[64]);
  assign t[384] = (x[67]);
  assign t[385] = (x[67]);
  assign t[386] = (x[70]);
  assign t[387] = (x[70]);
  assign t[388] = (x[73]);
  assign t[389] = (x[73]);
  assign t[38] = t[50] & t[51];
  assign t[390] = (x[76]);
  assign t[391] = (x[76]);
  assign t[392] = (x[79]);
  assign t[393] = (x[79]);
  assign t[394] = (x[82]);
  assign t[395] = (x[82]);
  assign t[396] = (x[85]);
  assign t[397] = (x[85]);
  assign t[398] = (x[88]);
  assign t[399] = (x[88]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[91]);
  assign t[401] = (x[91]);
  assign t[402] = (x[94]);
  assign t[403] = (x[94]);
  assign t[404] = (x[97]);
  assign t[405] = (x[97]);
  assign t[406] = (x[100]);
  assign t[407] = (x[100]);
  assign t[408] = (x[103]);
  assign t[409] = (x[103]);
  assign t[40] = t[54] & t[55];
  assign t[410] = (x[106]);
  assign t[411] = (x[106]);
  assign t[412] = (x[109]);
  assign t[413] = (x[109]);
  assign t[414] = (x[112]);
  assign t[415] = (x[112]);
  assign t[416] = (x[115]);
  assign t[417] = (x[115]);
  assign t[418] = (x[118]);
  assign t[419] = (x[118]);
  assign t[41] = t[54] & t[56];
  assign t[420] = (x[121]);
  assign t[421] = (x[121]);
  assign t[42] = t[57] & t[58];
  assign t[43] = t[59] & t[60];
  assign t[44] = t[61] & t[62];
  assign t[45] = ~(t[148] | t[149]);
  assign t[46] = ~(t[150] | t[151]);
  assign t[47] = ~(t[152]);
  assign t[48] = t[61] ^ t[59];
  assign t[49] = t[63] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[48] ^ t[65];
  assign t[51] = t[64] ^ t[66];
  assign t[52] = t[67] ^ t[68];
  assign t[53] = t[60] ^ t[69];
  assign t[54] = t[70] ^ t[71];
  assign t[55] = t[72] ^ t[73];
  assign t[56] = t[60] ^ t[74];
  assign t[57] = t[59] ^ t[54];
  assign t[58] = t[75] ^ t[51];
  assign t[59] = t[76] ^ t[77];
  assign t[5] = t[9] ? t[136] : x[3];
  assign t[60] = t[13] ? t[153] : t[78];
  assign t[61] = t[79] ^ t[80];
  assign t[62] = t[53] ^ t[81];
  assign t[63] = t[13] ? t[154] : t[82];
  assign t[64] = t[13] ? t[155] : t[83];
  assign t[65] = t[52] ^ t[54];
  assign t[66] = t[13] ? t[156] : t[84];
  assign t[67] = t[85] & t[86];
  assign t[68] = t[85] ^ t[87];
  assign t[69] = t[88] ^ t[89];
  assign t[6] = ~(t[10] ^ t[137]);
  assign t[70] = t[90] & t[91];
  assign t[71] = t[90] ^ t[87];
  assign t[72] = t[63] ^ t[66];
  assign t[73] = t[69] ^ t[92];
  assign t[74] = t[49] ^ t[93];
  assign t[75] = t[63] ^ t[94];
  assign t[76] = t[95] ^ t[96];
  assign t[77] = t[97] & t[90];
  assign t[78] = t[157] ^ t[158];
  assign t[79] = t[98] ^ t[99];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[100] & t[85];
  assign t[81] = t[93] ^ t[101];
  assign t[82] = t[159] ^ t[160];
  assign t[83] = t[161] ^ t[162];
  assign t[84] = t[163] ^ t[164];
  assign t[85] = t[102] ^ t[79];
  assign t[86] = t[102] & t[76];
  assign t[87] = t[103] & t[102];
  assign t[88] = t[13] ? t[165] : t[104];
  assign t[89] = t[13] ? t[166] : t[105];
  assign t[8] = ~(t[13]);
  assign t[90] = t[103] ^ t[76];
  assign t[91] = t[79] & t[103];
  assign t[92] = t[94] ^ t[60];
  assign t[93] = t[106] ^ t[94];
  assign t[94] = t[13] ? t[167] : t[107];
  assign t[95] = t[108] ^ t[99];
  assign t[96] = t[109] ^ t[62];
  assign t[97] = t[79] ^ t[87];
  assign t[98] = t[110] ^ t[111];
  assign t[99] = t[112] ^ t[113];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [120:0] x;
 output y;

 wire [413:0] t;
  assign t[0] = t[1] ? t[2] : t[134];
  assign t[100] = t[78] ^ t[88];
  assign t[101] = t[166] ^ t[167];
  assign t[102] = t[168] ^ t[169];
  assign t[103] = t[170] ^ t[171];
  assign t[104] = t[114] ^ t[115];
  assign t[105] = t[116] ^ t[115];
  assign t[106] = t[172] ^ t[173];
  assign t[107] = t[117] ^ t[118];
  assign t[108] = t[74] ^ t[119];
  assign t[109] = t[74] & t[119];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[52] & t[120];
  assign t[111] = t[121] ^ t[122];
  assign t[112] = t[52] ^ t[123];
  assign t[113] = t[54] ^ t[51];
  assign t[114] = t[124] ^ t[125];
  assign t[115] = t[126] ^ t[110];
  assign t[116] = t[127] ^ t[128];
  assign t[117] = t[123] & t[70];
  assign t[118] = t[77] & t[58];
  assign t[119] = t[58] ^ t[71];
  assign t[11] = ~(t[17]);
  assign t[120] = t[65] ^ t[129];
  assign t[121] = t[112] & t[113];
  assign t[122] = t[94] & t[51];
  assign t[123] = t[71] ^ t[130];
  assign t[124] = t[131] ^ t[118];
  assign t[125] = t[56] & t[76];
  assign t[126] = t[36] & t[132];
  assign t[127] = t[133] ^ t[122];
  assign t[128] = t[75] & t[54];
  assign t[129] = t[90] ^ t[49];
  assign t[12] = t[137] & t[18];
  assign t[130] = t[48] ^ t[70];
  assign t[131] = t[58] ^ t[129];
  assign t[132] = t[52] ^ t[66];
  assign t[133] = t[94] ^ t[51];
  assign t[134] = (t[174]);
  assign t[135] = (t[175]);
  assign t[136] = (t[176]);
  assign t[137] = (t[177]);
  assign t[138] = (t[178]);
  assign t[139] = (t[179]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[180]);
  assign t[141] = (t[181]);
  assign t[142] = (t[182]);
  assign t[143] = (t[183]);
  assign t[144] = (t[184]);
  assign t[145] = (t[185]);
  assign t[146] = (t[186]);
  assign t[147] = (t[187]);
  assign t[148] = (t[188]);
  assign t[149] = (t[189]);
  assign t[14] = ~(t[137]);
  assign t[150] = (t[190]);
  assign t[151] = (t[191]);
  assign t[152] = (t[192]);
  assign t[153] = (t[193]);
  assign t[154] = (t[194]);
  assign t[155] = (t[195]);
  assign t[156] = (t[196]);
  assign t[157] = (t[197]);
  assign t[158] = (t[198]);
  assign t[159] = (t[199]);
  assign t[15] = t[138] & t[139];
  assign t[160] = (t[200]);
  assign t[161] = (t[201]);
  assign t[162] = (t[202]);
  assign t[163] = (t[203]);
  assign t[164] = (t[204]);
  assign t[165] = (t[205]);
  assign t[166] = (t[206]);
  assign t[167] = (t[207]);
  assign t[168] = (t[208]);
  assign t[169] = (t[209]);
  assign t[16] = t[21] ^ t[22];
  assign t[170] = (t[210]);
  assign t[171] = (t[211]);
  assign t[172] = (t[212]);
  assign t[173] = (t[213]);
  assign t[174] = t[214] ^ x[2];
  assign t[175] = t[215] ^ x[6];
  assign t[176] = t[216] ^ x[9];
  assign t[177] = t[217] ^ x[12];
  assign t[178] = t[218] ^ x[15];
  assign t[179] = t[219] ^ x[18];
  assign t[17] = ~(t[137] & t[23]);
  assign t[180] = t[220] ^ x[21];
  assign t[181] = t[221] ^ x[24];
  assign t[182] = t[222] ^ x[27];
  assign t[183] = t[223] ^ x[30];
  assign t[184] = t[224] ^ x[33];
  assign t[185] = t[225] ^ x[36];
  assign t[186] = t[226] ^ x[39];
  assign t[187] = t[227] ^ x[42];
  assign t[188] = t[228] ^ x[45];
  assign t[189] = t[229] ^ x[48];
  assign t[18] = t[24] & t[25];
  assign t[190] = t[230] ^ x[51];
  assign t[191] = t[231] ^ x[54];
  assign t[192] = t[232] ^ x[57];
  assign t[193] = t[233] ^ x[60];
  assign t[194] = t[234] ^ x[63];
  assign t[195] = t[235] ^ x[66];
  assign t[196] = t[236] ^ x[69];
  assign t[197] = t[237] ^ x[72];
  assign t[198] = t[238] ^ x[75];
  assign t[199] = t[239] ^ x[78];
  assign t[19] = ~(t[140]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[81];
  assign t[201] = t[241] ^ x[84];
  assign t[202] = t[242] ^ x[87];
  assign t[203] = t[243] ^ x[90];
  assign t[204] = t[244] ^ x[93];
  assign t[205] = t[245] ^ x[96];
  assign t[206] = t[246] ^ x[99];
  assign t[207] = t[247] ^ x[102];
  assign t[208] = t[248] ^ x[105];
  assign t[209] = t[249] ^ x[108];
  assign t[20] = ~(t[137]);
  assign t[210] = t[250] ^ x[111];
  assign t[211] = t[251] ^ x[114];
  assign t[212] = t[252] ^ x[117];
  assign t[213] = t[253] ^ x[120];
  assign t[214] = (t[254] & ~t[255]);
  assign t[215] = (t[256] & ~t[257]);
  assign t[216] = (t[258] & ~t[259]);
  assign t[217] = (t[260] & ~t[261]);
  assign t[218] = (t[262] & ~t[263]);
  assign t[219] = (t[264] & ~t[265]);
  assign t[21] = t[26] ^ t[27];
  assign t[220] = (t[266] & ~t[267]);
  assign t[221] = (t[268] & ~t[269]);
  assign t[222] = (t[270] & ~t[271]);
  assign t[223] = (t[272] & ~t[273]);
  assign t[224] = (t[274] & ~t[275]);
  assign t[225] = (t[276] & ~t[277]);
  assign t[226] = (t[278] & ~t[279]);
  assign t[227] = (t[280] & ~t[281]);
  assign t[228] = (t[282] & ~t[283]);
  assign t[229] = (t[284] & ~t[285]);
  assign t[22] = t[28] ^ t[29];
  assign t[230] = (t[286] & ~t[287]);
  assign t[231] = (t[288] & ~t[289]);
  assign t[232] = (t[290] & ~t[291]);
  assign t[233] = (t[292] & ~t[293]);
  assign t[234] = (t[294] & ~t[295]);
  assign t[235] = (t[296] & ~t[297]);
  assign t[236] = (t[298] & ~t[299]);
  assign t[237] = (t[300] & ~t[301]);
  assign t[238] = (t[302] & ~t[303]);
  assign t[239] = (t[304] & ~t[305]);
  assign t[23] = ~(t[141] | t[30]);
  assign t[240] = (t[306] & ~t[307]);
  assign t[241] = (t[308] & ~t[309]);
  assign t[242] = (t[310] & ~t[311]);
  assign t[243] = (t[312] & ~t[313]);
  assign t[244] = (t[314] & ~t[315]);
  assign t[245] = (t[316] & ~t[317]);
  assign t[246] = (t[318] & ~t[319]);
  assign t[247] = (t[320] & ~t[321]);
  assign t[248] = (t[322] & ~t[323]);
  assign t[249] = (t[324] & ~t[325]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[250] = (t[326] & ~t[327]);
  assign t[251] = (t[328] & ~t[329]);
  assign t[252] = (t[330] & ~t[331]);
  assign t[253] = (t[332] & ~t[333]);
  assign t[254] = t[334] ^ x[2];
  assign t[255] = t[335] ^ x[1];
  assign t[256] = t[336] ^ x[6];
  assign t[257] = t[337] ^ x[5];
  assign t[258] = t[338] ^ x[9];
  assign t[259] = t[339] ^ x[8];
  assign t[25] = ~(t[33] | t[34]);
  assign t[260] = t[340] ^ x[12];
  assign t[261] = t[341] ^ x[11];
  assign t[262] = t[342] ^ x[15];
  assign t[263] = t[343] ^ x[14];
  assign t[264] = t[344] ^ x[18];
  assign t[265] = t[345] ^ x[17];
  assign t[266] = t[346] ^ x[21];
  assign t[267] = t[347] ^ x[20];
  assign t[268] = t[348] ^ x[24];
  assign t[269] = t[349] ^ x[23];
  assign t[26] = t[35] & t[36];
  assign t[270] = t[350] ^ x[27];
  assign t[271] = t[351] ^ x[26];
  assign t[272] = t[352] ^ x[30];
  assign t[273] = t[353] ^ x[29];
  assign t[274] = t[354] ^ x[33];
  assign t[275] = t[355] ^ x[32];
  assign t[276] = t[356] ^ x[36];
  assign t[277] = t[357] ^ x[35];
  assign t[278] = t[358] ^ x[39];
  assign t[279] = t[359] ^ x[38];
  assign t[27] = t[37] ^ t[38];
  assign t[280] = t[360] ^ x[42];
  assign t[281] = t[361] ^ x[41];
  assign t[282] = t[362] ^ x[45];
  assign t[283] = t[363] ^ x[44];
  assign t[284] = t[364] ^ x[48];
  assign t[285] = t[365] ^ x[47];
  assign t[286] = t[366] ^ x[51];
  assign t[287] = t[367] ^ x[50];
  assign t[288] = t[368] ^ x[54];
  assign t[289] = t[369] ^ x[53];
  assign t[28] = t[39] ^ t[40];
  assign t[290] = t[370] ^ x[57];
  assign t[291] = t[371] ^ x[56];
  assign t[292] = t[372] ^ x[60];
  assign t[293] = t[373] ^ x[59];
  assign t[294] = t[374] ^ x[63];
  assign t[295] = t[375] ^ x[62];
  assign t[296] = t[376] ^ x[66];
  assign t[297] = t[377] ^ x[65];
  assign t[298] = t[378] ^ x[69];
  assign t[299] = t[379] ^ x[68];
  assign t[29] = t[41] ^ t[42];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[380] ^ x[72];
  assign t[301] = t[381] ^ x[71];
  assign t[302] = t[382] ^ x[75];
  assign t[303] = t[383] ^ x[74];
  assign t[304] = t[384] ^ x[78];
  assign t[305] = t[385] ^ x[77];
  assign t[306] = t[386] ^ x[81];
  assign t[307] = t[387] ^ x[80];
  assign t[308] = t[388] ^ x[84];
  assign t[309] = t[389] ^ x[83];
  assign t[30] = ~(t[43] & t[44]);
  assign t[310] = t[390] ^ x[87];
  assign t[311] = t[391] ^ x[86];
  assign t[312] = t[392] ^ x[90];
  assign t[313] = t[393] ^ x[89];
  assign t[314] = t[394] ^ x[93];
  assign t[315] = t[395] ^ x[92];
  assign t[316] = t[396] ^ x[96];
  assign t[317] = t[397] ^ x[95];
  assign t[318] = t[398] ^ x[99];
  assign t[319] = t[399] ^ x[98];
  assign t[31] = ~(t[142] & t[143]);
  assign t[320] = t[400] ^ x[102];
  assign t[321] = t[401] ^ x[101];
  assign t[322] = t[402] ^ x[105];
  assign t[323] = t[403] ^ x[104];
  assign t[324] = t[404] ^ x[108];
  assign t[325] = t[405] ^ x[107];
  assign t[326] = t[406] ^ x[111];
  assign t[327] = t[407] ^ x[110];
  assign t[328] = t[408] ^ x[114];
  assign t[329] = t[409] ^ x[113];
  assign t[32] = ~(t[138] & t[144]);
  assign t[330] = t[410] ^ x[117];
  assign t[331] = t[411] ^ x[116];
  assign t[332] = t[412] ^ x[120];
  assign t[333] = t[413] ^ x[119];
  assign t[334] = (x[0]);
  assign t[335] = (x[0]);
  assign t[336] = (x[4]);
  assign t[337] = (x[4]);
  assign t[338] = (x[7]);
  assign t[339] = (x[7]);
  assign t[33] = ~(t[23]);
  assign t[340] = (x[10]);
  assign t[341] = (x[10]);
  assign t[342] = (x[13]);
  assign t[343] = (x[13]);
  assign t[344] = (x[16]);
  assign t[345] = (x[16]);
  assign t[346] = (x[19]);
  assign t[347] = (x[19]);
  assign t[348] = (x[22]);
  assign t[349] = (x[22]);
  assign t[34] = ~(t[145] & t[45]);
  assign t[350] = (x[25]);
  assign t[351] = (x[25]);
  assign t[352] = (x[28]);
  assign t[353] = (x[28]);
  assign t[354] = (x[31]);
  assign t[355] = (x[31]);
  assign t[356] = (x[34]);
  assign t[357] = (x[34]);
  assign t[358] = (x[37]);
  assign t[359] = (x[37]);
  assign t[35] = t[46] ^ t[47];
  assign t[360] = (x[40]);
  assign t[361] = (x[40]);
  assign t[362] = (x[43]);
  assign t[363] = (x[43]);
  assign t[364] = (x[46]);
  assign t[365] = (x[46]);
  assign t[366] = (x[49]);
  assign t[367] = (x[49]);
  assign t[368] = (x[52]);
  assign t[369] = (x[52]);
  assign t[36] = t[48] ^ t[49];
  assign t[370] = (x[55]);
  assign t[371] = (x[55]);
  assign t[372] = (x[58]);
  assign t[373] = (x[58]);
  assign t[374] = (x[61]);
  assign t[375] = (x[61]);
  assign t[376] = (x[64]);
  assign t[377] = (x[64]);
  assign t[378] = (x[67]);
  assign t[379] = (x[67]);
  assign t[37] = t[50] & t[51];
  assign t[380] = (x[70]);
  assign t[381] = (x[70]);
  assign t[382] = (x[73]);
  assign t[383] = (x[73]);
  assign t[384] = (x[76]);
  assign t[385] = (x[76]);
  assign t[386] = (x[79]);
  assign t[387] = (x[79]);
  assign t[388] = (x[82]);
  assign t[389] = (x[82]);
  assign t[38] = t[46] & t[52];
  assign t[390] = (x[85]);
  assign t[391] = (x[85]);
  assign t[392] = (x[88]);
  assign t[393] = (x[88]);
  assign t[394] = (x[91]);
  assign t[395] = (x[91]);
  assign t[396] = (x[94]);
  assign t[397] = (x[94]);
  assign t[398] = (x[97]);
  assign t[399] = (x[97]);
  assign t[39] = t[53] & t[54];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[100]);
  assign t[401] = (x[100]);
  assign t[402] = (x[103]);
  assign t[403] = (x[103]);
  assign t[404] = (x[106]);
  assign t[405] = (x[106]);
  assign t[406] = (x[109]);
  assign t[407] = (x[109]);
  assign t[408] = (x[112]);
  assign t[409] = (x[112]);
  assign t[40] = t[55] & t[56];
  assign t[410] = (x[115]);
  assign t[411] = (x[115]);
  assign t[412] = (x[118]);
  assign t[413] = (x[118]);
  assign t[41] = t[57] & t[58];
  assign t[42] = t[59] ^ t[60];
  assign t[43] = ~(t[146] | t[147]);
  assign t[44] = ~(t[148] | t[149]);
  assign t[45] = ~(t[150]);
  assign t[46] = t[61] ^ t[62];
  assign t[47] = t[53] ^ t[55];
  assign t[48] = t[13] ? t[151] : t[63];
  assign t[49] = t[13] ? t[152] : t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[61] ^ t[53];
  assign t[51] = t[65] ^ t[66];
  assign t[52] = t[67] ^ t[48];
  assign t[53] = t[68] ^ t[69];
  assign t[54] = t[70] ^ t[71];
  assign t[55] = t[72] ^ t[73];
  assign t[56] = t[74] ^ t[75];
  assign t[57] = t[62] ^ t[55];
  assign t[58] = t[52] ^ t[65];
  assign t[59] = t[55] & t[76];
  assign t[5] = t[9] ? t[135] : x[3];
  assign t[60] = t[57] & t[77];
  assign t[61] = t[78] ^ t[79];
  assign t[62] = t[80] ^ t[81];
  assign t[63] = t[153] ^ t[136];
  assign t[64] = t[154] ^ t[155];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[84] ^ t[49];
  assign t[67] = t[13] ? t[156] : t[85];
  assign t[68] = t[86] & t[87];
  assign t[69] = t[86] ^ t[88];
  assign t[6] = ~(t[10] ^ t[136]);
  assign t[70] = t[13] ? t[157] : t[89];
  assign t[71] = t[90] ^ t[84];
  assign t[72] = t[91] & t[92];
  assign t[73] = t[91] ^ t[88];
  assign t[74] = t[67] ^ t[49];
  assign t[75] = t[71] ^ t[93];
  assign t[76] = t[70] ^ t[58];
  assign t[77] = t[94] ^ t[36];
  assign t[78] = t[95] ^ t[96];
  assign t[79] = t[97] & t[86];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[98] ^ t[99];
  assign t[81] = t[100] & t[91];
  assign t[82] = t[13] ? t[158] : t[101];
  assign t[83] = t[13] ? t[159] : t[102];
  assign t[84] = t[13] ? t[160] : t[103];
  assign t[85] = t[161] ^ t[162];
  assign t[86] = t[104] ^ t[78];
  assign t[87] = t[104] & t[80];
  assign t[88] = t[105] & t[104];
  assign t[89] = t[163] ^ t[164];
  assign t[8] = ~(t[13]);
  assign t[90] = t[13] ? t[165] : t[106];
  assign t[91] = t[105] ^ t[80];
  assign t[92] = t[78] & t[105];
  assign t[93] = t[83] ^ t[70];
  assign t[94] = t[67] ^ t[83];
  assign t[95] = t[107] ^ t[108];
  assign t[96] = t[109] ^ t[110];
  assign t[97] = t[80] ^ t[88];
  assign t[98] = t[111] ^ t[96];
  assign t[99] = t[112] ^ t[113];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind241(x, y);
 input [120:0] x;
 output y;

 wire [413:0] t;
  assign t[0] = t[1] ? t[2] : t[134];
  assign t[100] = t[78] ^ t[88];
  assign t[101] = t[166] ^ t[167];
  assign t[102] = t[168] ^ t[169];
  assign t[103] = t[170] ^ t[171];
  assign t[104] = t[114] ^ t[115];
  assign t[105] = t[116] ^ t[115];
  assign t[106] = t[172] ^ t[173];
  assign t[107] = t[117] ^ t[118];
  assign t[108] = t[74] ^ t[119];
  assign t[109] = t[74] & t[119];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[52] & t[120];
  assign t[111] = t[121] ^ t[122];
  assign t[112] = t[52] ^ t[123];
  assign t[113] = t[54] ^ t[51];
  assign t[114] = t[124] ^ t[125];
  assign t[115] = t[126] ^ t[110];
  assign t[116] = t[127] ^ t[128];
  assign t[117] = t[123] & t[70];
  assign t[118] = t[77] & t[58];
  assign t[119] = t[58] ^ t[71];
  assign t[11] = ~(t[17]);
  assign t[120] = t[65] ^ t[129];
  assign t[121] = t[112] & t[113];
  assign t[122] = t[94] & t[51];
  assign t[123] = t[71] ^ t[130];
  assign t[124] = t[131] ^ t[118];
  assign t[125] = t[56] & t[76];
  assign t[126] = t[36] & t[132];
  assign t[127] = t[133] ^ t[122];
  assign t[128] = t[75] & t[54];
  assign t[129] = t[90] ^ t[49];
  assign t[12] = t[137] & t[18];
  assign t[130] = t[48] ^ t[70];
  assign t[131] = t[58] ^ t[129];
  assign t[132] = t[52] ^ t[66];
  assign t[133] = t[94] ^ t[51];
  assign t[134] = (t[174]);
  assign t[135] = (t[175]);
  assign t[136] = (t[176]);
  assign t[137] = (t[177]);
  assign t[138] = (t[178]);
  assign t[139] = (t[179]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[180]);
  assign t[141] = (t[181]);
  assign t[142] = (t[182]);
  assign t[143] = (t[183]);
  assign t[144] = (t[184]);
  assign t[145] = (t[185]);
  assign t[146] = (t[186]);
  assign t[147] = (t[187]);
  assign t[148] = (t[188]);
  assign t[149] = (t[189]);
  assign t[14] = ~(t[137]);
  assign t[150] = (t[190]);
  assign t[151] = (t[191]);
  assign t[152] = (t[192]);
  assign t[153] = (t[193]);
  assign t[154] = (t[194]);
  assign t[155] = (t[195]);
  assign t[156] = (t[196]);
  assign t[157] = (t[197]);
  assign t[158] = (t[198]);
  assign t[159] = (t[199]);
  assign t[15] = t[138] & t[139];
  assign t[160] = (t[200]);
  assign t[161] = (t[201]);
  assign t[162] = (t[202]);
  assign t[163] = (t[203]);
  assign t[164] = (t[204]);
  assign t[165] = (t[205]);
  assign t[166] = (t[206]);
  assign t[167] = (t[207]);
  assign t[168] = (t[208]);
  assign t[169] = (t[209]);
  assign t[16] = t[21] ^ t[22];
  assign t[170] = (t[210]);
  assign t[171] = (t[211]);
  assign t[172] = (t[212]);
  assign t[173] = (t[213]);
  assign t[174] = t[214] ^ x[2];
  assign t[175] = t[215] ^ x[6];
  assign t[176] = t[216] ^ x[9];
  assign t[177] = t[217] ^ x[12];
  assign t[178] = t[218] ^ x[15];
  assign t[179] = t[219] ^ x[18];
  assign t[17] = ~(t[137] & t[23]);
  assign t[180] = t[220] ^ x[21];
  assign t[181] = t[221] ^ x[24];
  assign t[182] = t[222] ^ x[27];
  assign t[183] = t[223] ^ x[30];
  assign t[184] = t[224] ^ x[33];
  assign t[185] = t[225] ^ x[36];
  assign t[186] = t[226] ^ x[39];
  assign t[187] = t[227] ^ x[42];
  assign t[188] = t[228] ^ x[45];
  assign t[189] = t[229] ^ x[48];
  assign t[18] = t[24] & t[25];
  assign t[190] = t[230] ^ x[51];
  assign t[191] = t[231] ^ x[54];
  assign t[192] = t[232] ^ x[57];
  assign t[193] = t[233] ^ x[60];
  assign t[194] = t[234] ^ x[63];
  assign t[195] = t[235] ^ x[66];
  assign t[196] = t[236] ^ x[69];
  assign t[197] = t[237] ^ x[72];
  assign t[198] = t[238] ^ x[75];
  assign t[199] = t[239] ^ x[78];
  assign t[19] = ~(t[140]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[81];
  assign t[201] = t[241] ^ x[84];
  assign t[202] = t[242] ^ x[87];
  assign t[203] = t[243] ^ x[90];
  assign t[204] = t[244] ^ x[93];
  assign t[205] = t[245] ^ x[96];
  assign t[206] = t[246] ^ x[99];
  assign t[207] = t[247] ^ x[102];
  assign t[208] = t[248] ^ x[105];
  assign t[209] = t[249] ^ x[108];
  assign t[20] = ~(t[137]);
  assign t[210] = t[250] ^ x[111];
  assign t[211] = t[251] ^ x[114];
  assign t[212] = t[252] ^ x[117];
  assign t[213] = t[253] ^ x[120];
  assign t[214] = (t[254] & ~t[255]);
  assign t[215] = (t[256] & ~t[257]);
  assign t[216] = (t[258] & ~t[259]);
  assign t[217] = (t[260] & ~t[261]);
  assign t[218] = (t[262] & ~t[263]);
  assign t[219] = (t[264] & ~t[265]);
  assign t[21] = t[26] ^ t[27];
  assign t[220] = (t[266] & ~t[267]);
  assign t[221] = (t[268] & ~t[269]);
  assign t[222] = (t[270] & ~t[271]);
  assign t[223] = (t[272] & ~t[273]);
  assign t[224] = (t[274] & ~t[275]);
  assign t[225] = (t[276] & ~t[277]);
  assign t[226] = (t[278] & ~t[279]);
  assign t[227] = (t[280] & ~t[281]);
  assign t[228] = (t[282] & ~t[283]);
  assign t[229] = (t[284] & ~t[285]);
  assign t[22] = t[28] ^ t[29];
  assign t[230] = (t[286] & ~t[287]);
  assign t[231] = (t[288] & ~t[289]);
  assign t[232] = (t[290] & ~t[291]);
  assign t[233] = (t[292] & ~t[293]);
  assign t[234] = (t[294] & ~t[295]);
  assign t[235] = (t[296] & ~t[297]);
  assign t[236] = (t[298] & ~t[299]);
  assign t[237] = (t[300] & ~t[301]);
  assign t[238] = (t[302] & ~t[303]);
  assign t[239] = (t[304] & ~t[305]);
  assign t[23] = ~(t[141] | t[30]);
  assign t[240] = (t[306] & ~t[307]);
  assign t[241] = (t[308] & ~t[309]);
  assign t[242] = (t[310] & ~t[311]);
  assign t[243] = (t[312] & ~t[313]);
  assign t[244] = (t[314] & ~t[315]);
  assign t[245] = (t[316] & ~t[317]);
  assign t[246] = (t[318] & ~t[319]);
  assign t[247] = (t[320] & ~t[321]);
  assign t[248] = (t[322] & ~t[323]);
  assign t[249] = (t[324] & ~t[325]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[250] = (t[326] & ~t[327]);
  assign t[251] = (t[328] & ~t[329]);
  assign t[252] = (t[330] & ~t[331]);
  assign t[253] = (t[332] & ~t[333]);
  assign t[254] = t[334] ^ x[2];
  assign t[255] = t[335] ^ x[1];
  assign t[256] = t[336] ^ x[6];
  assign t[257] = t[337] ^ x[5];
  assign t[258] = t[338] ^ x[9];
  assign t[259] = t[339] ^ x[8];
  assign t[25] = ~(t[33] | t[34]);
  assign t[260] = t[340] ^ x[12];
  assign t[261] = t[341] ^ x[11];
  assign t[262] = t[342] ^ x[15];
  assign t[263] = t[343] ^ x[14];
  assign t[264] = t[344] ^ x[18];
  assign t[265] = t[345] ^ x[17];
  assign t[266] = t[346] ^ x[21];
  assign t[267] = t[347] ^ x[20];
  assign t[268] = t[348] ^ x[24];
  assign t[269] = t[349] ^ x[23];
  assign t[26] = t[35] & t[36];
  assign t[270] = t[350] ^ x[27];
  assign t[271] = t[351] ^ x[26];
  assign t[272] = t[352] ^ x[30];
  assign t[273] = t[353] ^ x[29];
  assign t[274] = t[354] ^ x[33];
  assign t[275] = t[355] ^ x[32];
  assign t[276] = t[356] ^ x[36];
  assign t[277] = t[357] ^ x[35];
  assign t[278] = t[358] ^ x[39];
  assign t[279] = t[359] ^ x[38];
  assign t[27] = t[37] ^ t[38];
  assign t[280] = t[360] ^ x[42];
  assign t[281] = t[361] ^ x[41];
  assign t[282] = t[362] ^ x[45];
  assign t[283] = t[363] ^ x[44];
  assign t[284] = t[364] ^ x[48];
  assign t[285] = t[365] ^ x[47];
  assign t[286] = t[366] ^ x[51];
  assign t[287] = t[367] ^ x[50];
  assign t[288] = t[368] ^ x[54];
  assign t[289] = t[369] ^ x[53];
  assign t[28] = t[39] ^ t[40];
  assign t[290] = t[370] ^ x[57];
  assign t[291] = t[371] ^ x[56];
  assign t[292] = t[372] ^ x[60];
  assign t[293] = t[373] ^ x[59];
  assign t[294] = t[374] ^ x[63];
  assign t[295] = t[375] ^ x[62];
  assign t[296] = t[376] ^ x[66];
  assign t[297] = t[377] ^ x[65];
  assign t[298] = t[378] ^ x[69];
  assign t[299] = t[379] ^ x[68];
  assign t[29] = t[41] ^ t[42];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[380] ^ x[72];
  assign t[301] = t[381] ^ x[71];
  assign t[302] = t[382] ^ x[75];
  assign t[303] = t[383] ^ x[74];
  assign t[304] = t[384] ^ x[78];
  assign t[305] = t[385] ^ x[77];
  assign t[306] = t[386] ^ x[81];
  assign t[307] = t[387] ^ x[80];
  assign t[308] = t[388] ^ x[84];
  assign t[309] = t[389] ^ x[83];
  assign t[30] = ~(t[43] & t[44]);
  assign t[310] = t[390] ^ x[87];
  assign t[311] = t[391] ^ x[86];
  assign t[312] = t[392] ^ x[90];
  assign t[313] = t[393] ^ x[89];
  assign t[314] = t[394] ^ x[93];
  assign t[315] = t[395] ^ x[92];
  assign t[316] = t[396] ^ x[96];
  assign t[317] = t[397] ^ x[95];
  assign t[318] = t[398] ^ x[99];
  assign t[319] = t[399] ^ x[98];
  assign t[31] = ~(t[142] & t[143]);
  assign t[320] = t[400] ^ x[102];
  assign t[321] = t[401] ^ x[101];
  assign t[322] = t[402] ^ x[105];
  assign t[323] = t[403] ^ x[104];
  assign t[324] = t[404] ^ x[108];
  assign t[325] = t[405] ^ x[107];
  assign t[326] = t[406] ^ x[111];
  assign t[327] = t[407] ^ x[110];
  assign t[328] = t[408] ^ x[114];
  assign t[329] = t[409] ^ x[113];
  assign t[32] = ~(t[138] & t[144]);
  assign t[330] = t[410] ^ x[117];
  assign t[331] = t[411] ^ x[116];
  assign t[332] = t[412] ^ x[120];
  assign t[333] = t[413] ^ x[119];
  assign t[334] = (x[0]);
  assign t[335] = (x[0]);
  assign t[336] = (x[4]);
  assign t[337] = (x[4]);
  assign t[338] = (x[7]);
  assign t[339] = (x[7]);
  assign t[33] = ~(t[23]);
  assign t[340] = (x[10]);
  assign t[341] = (x[10]);
  assign t[342] = (x[13]);
  assign t[343] = (x[13]);
  assign t[344] = (x[16]);
  assign t[345] = (x[16]);
  assign t[346] = (x[19]);
  assign t[347] = (x[19]);
  assign t[348] = (x[22]);
  assign t[349] = (x[22]);
  assign t[34] = ~(t[145] & t[45]);
  assign t[350] = (x[25]);
  assign t[351] = (x[25]);
  assign t[352] = (x[28]);
  assign t[353] = (x[28]);
  assign t[354] = (x[31]);
  assign t[355] = (x[31]);
  assign t[356] = (x[34]);
  assign t[357] = (x[34]);
  assign t[358] = (x[37]);
  assign t[359] = (x[37]);
  assign t[35] = t[46] ^ t[47];
  assign t[360] = (x[40]);
  assign t[361] = (x[40]);
  assign t[362] = (x[43]);
  assign t[363] = (x[43]);
  assign t[364] = (x[46]);
  assign t[365] = (x[46]);
  assign t[366] = (x[49]);
  assign t[367] = (x[49]);
  assign t[368] = (x[52]);
  assign t[369] = (x[52]);
  assign t[36] = t[48] ^ t[49];
  assign t[370] = (x[55]);
  assign t[371] = (x[55]);
  assign t[372] = (x[58]);
  assign t[373] = (x[58]);
  assign t[374] = (x[61]);
  assign t[375] = (x[61]);
  assign t[376] = (x[64]);
  assign t[377] = (x[64]);
  assign t[378] = (x[67]);
  assign t[379] = (x[67]);
  assign t[37] = t[50] & t[51];
  assign t[380] = (x[70]);
  assign t[381] = (x[70]);
  assign t[382] = (x[73]);
  assign t[383] = (x[73]);
  assign t[384] = (x[76]);
  assign t[385] = (x[76]);
  assign t[386] = (x[79]);
  assign t[387] = (x[79]);
  assign t[388] = (x[82]);
  assign t[389] = (x[82]);
  assign t[38] = t[46] & t[52];
  assign t[390] = (x[85]);
  assign t[391] = (x[85]);
  assign t[392] = (x[88]);
  assign t[393] = (x[88]);
  assign t[394] = (x[91]);
  assign t[395] = (x[91]);
  assign t[396] = (x[94]);
  assign t[397] = (x[94]);
  assign t[398] = (x[97]);
  assign t[399] = (x[97]);
  assign t[39] = t[53] & t[54];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[100]);
  assign t[401] = (x[100]);
  assign t[402] = (x[103]);
  assign t[403] = (x[103]);
  assign t[404] = (x[106]);
  assign t[405] = (x[106]);
  assign t[406] = (x[109]);
  assign t[407] = (x[109]);
  assign t[408] = (x[112]);
  assign t[409] = (x[112]);
  assign t[40] = t[55] & t[56];
  assign t[410] = (x[115]);
  assign t[411] = (x[115]);
  assign t[412] = (x[118]);
  assign t[413] = (x[118]);
  assign t[41] = t[57] & t[58];
  assign t[42] = t[59] ^ t[60];
  assign t[43] = ~(t[146] | t[147]);
  assign t[44] = ~(t[148] | t[149]);
  assign t[45] = ~(t[150]);
  assign t[46] = t[61] ^ t[62];
  assign t[47] = t[53] ^ t[55];
  assign t[48] = t[13] ? t[151] : t[63];
  assign t[49] = t[13] ? t[152] : t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[61] ^ t[53];
  assign t[51] = t[65] ^ t[66];
  assign t[52] = t[67] ^ t[48];
  assign t[53] = t[68] ^ t[69];
  assign t[54] = t[70] ^ t[71];
  assign t[55] = t[72] ^ t[73];
  assign t[56] = t[74] ^ t[75];
  assign t[57] = t[62] ^ t[55];
  assign t[58] = t[52] ^ t[65];
  assign t[59] = t[55] & t[76];
  assign t[5] = t[9] ? t[135] : x[3];
  assign t[60] = t[57] & t[77];
  assign t[61] = t[78] ^ t[79];
  assign t[62] = t[80] ^ t[81];
  assign t[63] = t[153] ^ t[136];
  assign t[64] = t[154] ^ t[155];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[84] ^ t[49];
  assign t[67] = t[13] ? t[156] : t[85];
  assign t[68] = t[86] & t[87];
  assign t[69] = t[86] ^ t[88];
  assign t[6] = ~(t[10] ^ t[136]);
  assign t[70] = t[13] ? t[157] : t[89];
  assign t[71] = t[90] ^ t[84];
  assign t[72] = t[91] & t[92];
  assign t[73] = t[91] ^ t[88];
  assign t[74] = t[67] ^ t[49];
  assign t[75] = t[71] ^ t[93];
  assign t[76] = t[70] ^ t[58];
  assign t[77] = t[94] ^ t[36];
  assign t[78] = t[95] ^ t[96];
  assign t[79] = t[97] & t[86];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[98] ^ t[99];
  assign t[81] = t[100] & t[91];
  assign t[82] = t[13] ? t[158] : t[101];
  assign t[83] = t[13] ? t[159] : t[102];
  assign t[84] = t[13] ? t[160] : t[103];
  assign t[85] = t[161] ^ t[162];
  assign t[86] = t[104] ^ t[78];
  assign t[87] = t[104] & t[80];
  assign t[88] = t[105] & t[104];
  assign t[89] = t[163] ^ t[164];
  assign t[8] = ~(t[13]);
  assign t[90] = t[13] ? t[165] : t[106];
  assign t[91] = t[105] ^ t[80];
  assign t[92] = t[78] & t[105];
  assign t[93] = t[83] ^ t[70];
  assign t[94] = t[67] ^ t[83];
  assign t[95] = t[107] ^ t[108];
  assign t[96] = t[109] ^ t[110];
  assign t[97] = t[80] ^ t[88];
  assign t[98] = t[111] ^ t[96];
  assign t[99] = t[112] ^ t[113];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [120:0] x;
 output y;

 wire [412:0] t;
  assign t[0] = t[1] ? t[2] : t[133];
  assign t[100] = t[36] ^ t[50];
  assign t[101] = t[36] & t[50];
  assign t[102] = t[59] & t[58];
  assign t[103] = t[112] ^ t[87];
  assign t[104] = t[54] ^ t[113];
  assign t[105] = t[69] ^ t[80];
  assign t[106] = t[171] ^ t[172];
  assign t[107] = t[114] ^ t[115];
  assign t[108] = t[116] ^ t[102];
  assign t[109] = t[117] ^ t[118];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[71] & t[74];
  assign t[111] = t[119] & t[66];
  assign t[112] = t[120] ^ t[121];
  assign t[113] = t[122] ^ t[123];
  assign t[114] = t[124] ^ t[111];
  assign t[115] = t[125] & t[126];
  assign t[116] = t[127] & t[128];
  assign t[117] = t[129] ^ t[121];
  assign t[118] = t[130] & t[122];
  assign t[119] = t[52] ^ t[127];
  assign t[11] = ~(t[17]);
  assign t[120] = t[54] & t[113];
  assign t[121] = t[52] & t[123];
  assign t[122] = t[74] ^ t[67];
  assign t[123] = t[75] ^ t[131];
  assign t[124] = t[66] ^ t[76];
  assign t[125] = t[36] ^ t[130];
  assign t[126] = t[74] ^ t[66];
  assign t[127] = t[77] ^ t[49];
  assign t[128] = t[59] ^ t[131];
  assign t[129] = t[52] ^ t[123];
  assign t[12] = t[136] & t[18];
  assign t[130] = t[67] ^ t[132];
  assign t[131] = t[84] ^ t[49];
  assign t[132] = t[68] ^ t[74];
  assign t[133] = (t[173]);
  assign t[134] = (t[174]);
  assign t[135] = (t[175]);
  assign t[136] = (t[176]);
  assign t[137] = (t[177]);
  assign t[138] = (t[178]);
  assign t[139] = (t[179]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[180]);
  assign t[141] = (t[181]);
  assign t[142] = (t[182]);
  assign t[143] = (t[183]);
  assign t[144] = (t[184]);
  assign t[145] = (t[185]);
  assign t[146] = (t[186]);
  assign t[147] = (t[187]);
  assign t[148] = (t[188]);
  assign t[149] = (t[189]);
  assign t[14] = ~(t[136]);
  assign t[150] = (t[190]);
  assign t[151] = (t[191]);
  assign t[152] = (t[192]);
  assign t[153] = (t[193]);
  assign t[154] = (t[194]);
  assign t[155] = (t[195]);
  assign t[156] = (t[196]);
  assign t[157] = (t[197]);
  assign t[158] = (t[198]);
  assign t[159] = (t[199]);
  assign t[15] = t[137] & t[138];
  assign t[160] = (t[200]);
  assign t[161] = (t[201]);
  assign t[162] = (t[202]);
  assign t[163] = (t[203]);
  assign t[164] = (t[204]);
  assign t[165] = (t[205]);
  assign t[166] = (t[206]);
  assign t[167] = (t[207]);
  assign t[168] = (t[208]);
  assign t[169] = (t[209]);
  assign t[16] = ~(t[21] ^ t[22]);
  assign t[170] = (t[210]);
  assign t[171] = (t[211]);
  assign t[172] = (t[212]);
  assign t[173] = t[213] ^ x[2];
  assign t[174] = t[214] ^ x[6];
  assign t[175] = t[215] ^ x[9];
  assign t[176] = t[216] ^ x[12];
  assign t[177] = t[217] ^ x[15];
  assign t[178] = t[218] ^ x[18];
  assign t[179] = t[219] ^ x[21];
  assign t[17] = ~(t[136] & t[23]);
  assign t[180] = t[220] ^ x[24];
  assign t[181] = t[221] ^ x[27];
  assign t[182] = t[222] ^ x[30];
  assign t[183] = t[223] ^ x[33];
  assign t[184] = t[224] ^ x[36];
  assign t[185] = t[225] ^ x[39];
  assign t[186] = t[226] ^ x[42];
  assign t[187] = t[227] ^ x[45];
  assign t[188] = t[228] ^ x[48];
  assign t[189] = t[229] ^ x[51];
  assign t[18] = t[24] & t[25];
  assign t[190] = t[230] ^ x[54];
  assign t[191] = t[231] ^ x[57];
  assign t[192] = t[232] ^ x[60];
  assign t[193] = t[233] ^ x[63];
  assign t[194] = t[234] ^ x[66];
  assign t[195] = t[235] ^ x[69];
  assign t[196] = t[236] ^ x[72];
  assign t[197] = t[237] ^ x[75];
  assign t[198] = t[238] ^ x[78];
  assign t[199] = t[239] ^ x[81];
  assign t[19] = ~(t[139]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[84];
  assign t[201] = t[241] ^ x[87];
  assign t[202] = t[242] ^ x[90];
  assign t[203] = t[243] ^ x[93];
  assign t[204] = t[244] ^ x[96];
  assign t[205] = t[245] ^ x[99];
  assign t[206] = t[246] ^ x[102];
  assign t[207] = t[247] ^ x[105];
  assign t[208] = t[248] ^ x[108];
  assign t[209] = t[249] ^ x[111];
  assign t[20] = ~(t[136]);
  assign t[210] = t[250] ^ x[114];
  assign t[211] = t[251] ^ x[117];
  assign t[212] = t[252] ^ x[120];
  assign t[213] = (t[253] & ~t[254]);
  assign t[214] = (t[255] & ~t[256]);
  assign t[215] = (t[257] & ~t[258]);
  assign t[216] = (t[259] & ~t[260]);
  assign t[217] = (t[261] & ~t[262]);
  assign t[218] = (t[263] & ~t[264]);
  assign t[219] = (t[265] & ~t[266]);
  assign t[21] = t[26] ^ t[27];
  assign t[220] = (t[267] & ~t[268]);
  assign t[221] = (t[269] & ~t[270]);
  assign t[222] = (t[271] & ~t[272]);
  assign t[223] = (t[273] & ~t[274]);
  assign t[224] = (t[275] & ~t[276]);
  assign t[225] = (t[277] & ~t[278]);
  assign t[226] = (t[279] & ~t[280]);
  assign t[227] = (t[281] & ~t[282]);
  assign t[228] = (t[283] & ~t[284]);
  assign t[229] = (t[285] & ~t[286]);
  assign t[22] = t[28] ^ t[29];
  assign t[230] = (t[287] & ~t[288]);
  assign t[231] = (t[289] & ~t[290]);
  assign t[232] = (t[291] & ~t[292]);
  assign t[233] = (t[293] & ~t[294]);
  assign t[234] = (t[295] & ~t[296]);
  assign t[235] = (t[297] & ~t[298]);
  assign t[236] = (t[299] & ~t[300]);
  assign t[237] = (t[301] & ~t[302]);
  assign t[238] = (t[303] & ~t[304]);
  assign t[239] = (t[305] & ~t[306]);
  assign t[23] = ~(t[140] | t[30]);
  assign t[240] = (t[307] & ~t[308]);
  assign t[241] = (t[309] & ~t[310]);
  assign t[242] = (t[311] & ~t[312]);
  assign t[243] = (t[313] & ~t[314]);
  assign t[244] = (t[315] & ~t[316]);
  assign t[245] = (t[317] & ~t[318]);
  assign t[246] = (t[319] & ~t[320]);
  assign t[247] = (t[321] & ~t[322]);
  assign t[248] = (t[323] & ~t[324]);
  assign t[249] = (t[325] & ~t[326]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[250] = (t[327] & ~t[328]);
  assign t[251] = (t[329] & ~t[330]);
  assign t[252] = (t[331] & ~t[332]);
  assign t[253] = t[333] ^ x[2];
  assign t[254] = t[334] ^ x[1];
  assign t[255] = t[335] ^ x[6];
  assign t[256] = t[336] ^ x[5];
  assign t[257] = t[337] ^ x[9];
  assign t[258] = t[338] ^ x[8];
  assign t[259] = t[339] ^ x[12];
  assign t[25] = ~(t[33] | t[34]);
  assign t[260] = t[340] ^ x[11];
  assign t[261] = t[341] ^ x[15];
  assign t[262] = t[342] ^ x[14];
  assign t[263] = t[343] ^ x[18];
  assign t[264] = t[344] ^ x[17];
  assign t[265] = t[345] ^ x[21];
  assign t[266] = t[346] ^ x[20];
  assign t[267] = t[347] ^ x[24];
  assign t[268] = t[348] ^ x[23];
  assign t[269] = t[349] ^ x[27];
  assign t[26] = t[35] & t[36];
  assign t[270] = t[350] ^ x[26];
  assign t[271] = t[351] ^ x[30];
  assign t[272] = t[352] ^ x[29];
  assign t[273] = t[353] ^ x[33];
  assign t[274] = t[354] ^ x[32];
  assign t[275] = t[355] ^ x[36];
  assign t[276] = t[356] ^ x[35];
  assign t[277] = t[357] ^ x[39];
  assign t[278] = t[358] ^ x[38];
  assign t[279] = t[359] ^ x[42];
  assign t[27] = t[37] ^ t[38];
  assign t[280] = t[360] ^ x[41];
  assign t[281] = t[361] ^ x[45];
  assign t[282] = t[362] ^ x[44];
  assign t[283] = t[363] ^ x[48];
  assign t[284] = t[364] ^ x[47];
  assign t[285] = t[365] ^ x[51];
  assign t[286] = t[366] ^ x[50];
  assign t[287] = t[367] ^ x[54];
  assign t[288] = t[368] ^ x[53];
  assign t[289] = t[369] ^ x[57];
  assign t[28] = t[39] ^ t[40];
  assign t[290] = t[370] ^ x[56];
  assign t[291] = t[371] ^ x[60];
  assign t[292] = t[372] ^ x[59];
  assign t[293] = t[373] ^ x[63];
  assign t[294] = t[374] ^ x[62];
  assign t[295] = t[375] ^ x[66];
  assign t[296] = t[376] ^ x[65];
  assign t[297] = t[377] ^ x[69];
  assign t[298] = t[378] ^ x[68];
  assign t[299] = t[379] ^ x[72];
  assign t[29] = t[41] ^ t[42];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[380] ^ x[71];
  assign t[301] = t[381] ^ x[75];
  assign t[302] = t[382] ^ x[74];
  assign t[303] = t[383] ^ x[78];
  assign t[304] = t[384] ^ x[77];
  assign t[305] = t[385] ^ x[81];
  assign t[306] = t[386] ^ x[80];
  assign t[307] = t[387] ^ x[84];
  assign t[308] = t[388] ^ x[83];
  assign t[309] = t[389] ^ x[87];
  assign t[30] = ~(t[43] & t[44]);
  assign t[310] = t[390] ^ x[86];
  assign t[311] = t[391] ^ x[90];
  assign t[312] = t[392] ^ x[89];
  assign t[313] = t[393] ^ x[93];
  assign t[314] = t[394] ^ x[92];
  assign t[315] = t[395] ^ x[96];
  assign t[316] = t[396] ^ x[95];
  assign t[317] = t[397] ^ x[99];
  assign t[318] = t[398] ^ x[98];
  assign t[319] = t[399] ^ x[102];
  assign t[31] = ~(t[141] & t[137]);
  assign t[320] = t[400] ^ x[101];
  assign t[321] = t[401] ^ x[105];
  assign t[322] = t[402] ^ x[104];
  assign t[323] = t[403] ^ x[108];
  assign t[324] = t[404] ^ x[107];
  assign t[325] = t[405] ^ x[111];
  assign t[326] = t[406] ^ x[110];
  assign t[327] = t[407] ^ x[114];
  assign t[328] = t[408] ^ x[113];
  assign t[329] = t[409] ^ x[117];
  assign t[32] = ~(t[142] & t[143]);
  assign t[330] = t[410] ^ x[116];
  assign t[331] = t[411] ^ x[120];
  assign t[332] = t[412] ^ x[119];
  assign t[333] = (x[0]);
  assign t[334] = (x[0]);
  assign t[335] = (x[4]);
  assign t[336] = (x[4]);
  assign t[337] = (x[7]);
  assign t[338] = (x[7]);
  assign t[339] = (x[10]);
  assign t[33] = ~(t[23]);
  assign t[340] = (x[10]);
  assign t[341] = (x[13]);
  assign t[342] = (x[13]);
  assign t[343] = (x[16]);
  assign t[344] = (x[16]);
  assign t[345] = (x[19]);
  assign t[346] = (x[19]);
  assign t[347] = (x[22]);
  assign t[348] = (x[22]);
  assign t[349] = (x[25]);
  assign t[34] = ~(t[144] & t[45]);
  assign t[350] = (x[25]);
  assign t[351] = (x[28]);
  assign t[352] = (x[28]);
  assign t[353] = (x[31]);
  assign t[354] = (x[31]);
  assign t[355] = (x[34]);
  assign t[356] = (x[34]);
  assign t[357] = (x[37]);
  assign t[358] = (x[37]);
  assign t[359] = (x[40]);
  assign t[35] = t[46] ^ t[47];
  assign t[360] = (x[40]);
  assign t[361] = (x[43]);
  assign t[362] = (x[43]);
  assign t[363] = (x[46]);
  assign t[364] = (x[46]);
  assign t[365] = (x[49]);
  assign t[366] = (x[49]);
  assign t[367] = (x[52]);
  assign t[368] = (x[52]);
  assign t[369] = (x[55]);
  assign t[36] = t[48] ^ t[49];
  assign t[370] = (x[55]);
  assign t[371] = (x[58]);
  assign t[372] = (x[58]);
  assign t[373] = (x[61]);
  assign t[374] = (x[61]);
  assign t[375] = (x[64]);
  assign t[376] = (x[64]);
  assign t[377] = (x[67]);
  assign t[378] = (x[67]);
  assign t[379] = (x[70]);
  assign t[37] = t[35] & t[50];
  assign t[380] = (x[70]);
  assign t[381] = (x[73]);
  assign t[382] = (x[73]);
  assign t[383] = (x[76]);
  assign t[384] = (x[76]);
  assign t[385] = (x[79]);
  assign t[386] = (x[79]);
  assign t[387] = (x[82]);
  assign t[388] = (x[82]);
  assign t[389] = (x[85]);
  assign t[38] = t[51] & t[52];
  assign t[390] = (x[85]);
  assign t[391] = (x[88]);
  assign t[392] = (x[88]);
  assign t[393] = (x[91]);
  assign t[394] = (x[91]);
  assign t[395] = (x[94]);
  assign t[396] = (x[94]);
  assign t[397] = (x[97]);
  assign t[398] = (x[97]);
  assign t[399] = (x[100]);
  assign t[39] = t[53] & t[54];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[100]);
  assign t[401] = (x[103]);
  assign t[402] = (x[103]);
  assign t[403] = (x[106]);
  assign t[404] = (x[106]);
  assign t[405] = (x[109]);
  assign t[406] = (x[109]);
  assign t[407] = (x[112]);
  assign t[408] = (x[112]);
  assign t[409] = (x[115]);
  assign t[40] = t[55] ^ t[56];
  assign t[410] = (x[115]);
  assign t[411] = (x[118]);
  assign t[412] = (x[118]);
  assign t[41] = t[57] & t[58];
  assign t[42] = t[57] & t[59];
  assign t[43] = ~(t[145] | t[146]);
  assign t[44] = ~(t[147] | t[148]);
  assign t[45] = ~(t[149]);
  assign t[46] = t[60] ^ t[61];
  assign t[47] = t[62] ^ t[63];
  assign t[48] = t[13] ? t[150] : t[64];
  assign t[49] = t[13] ? t[151] : t[65];
  assign t[4] = ~(t[8]);
  assign t[50] = t[66] ^ t[67];
  assign t[51] = t[53] ^ t[46];
  assign t[52] = t[48] ^ t[68];
  assign t[53] = t[69] ^ t[70];
  assign t[54] = t[59] ^ t[71];
  assign t[55] = t[72] & t[66];
  assign t[56] = t[73] & t[74];
  assign t[57] = t[53] ^ t[73];
  assign t[58] = t[75] ^ t[76];
  assign t[59] = t[48] ^ t[77];
  assign t[5] = t[9] ? t[134] : x[3];
  assign t[60] = t[78] & t[79];
  assign t[61] = t[78] ^ t[80];
  assign t[62] = t[81] & t[82];
  assign t[63] = t[81] ^ t[80];
  assign t[64] = t[152] ^ t[153];
  assign t[65] = t[154] ^ t[155];
  assign t[66] = t[59] ^ t[75];
  assign t[67] = t[83] ^ t[84];
  assign t[68] = t[13] ? t[156] : t[85];
  assign t[69] = t[86] ^ t[87];
  assign t[6] = ~(t[10] ^ t[135]);
  assign t[70] = t[88] & t[78];
  assign t[71] = t[67] ^ t[89];
  assign t[72] = t[73] ^ t[47];
  assign t[73] = t[90] ^ t[91];
  assign t[74] = t[13] ? t[157] : t[92];
  assign t[75] = t[93] ^ t[68];
  assign t[76] = t[83] ^ t[49];
  assign t[77] = t[13] ? t[158] : t[94];
  assign t[78] = t[95] ^ t[69];
  assign t[79] = t[95] & t[90];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[96] & t[95];
  assign t[81] = t[96] ^ t[90];
  assign t[82] = t[69] & t[96];
  assign t[83] = t[13] ? t[159] : t[97];
  assign t[84] = t[13] ? t[160] : t[98];
  assign t[85] = t[161] ^ t[162];
  assign t[86] = t[99] ^ t[100];
  assign t[87] = t[101] ^ t[102];
  assign t[88] = t[90] ^ t[80];
  assign t[89] = t[77] ^ t[74];
  assign t[8] = ~(t[13]);
  assign t[90] = t[103] ^ t[104];
  assign t[91] = t[105] & t[81];
  assign t[92] = t[163] ^ t[164];
  assign t[93] = t[13] ? t[165] : t[106];
  assign t[94] = t[166] ^ t[167];
  assign t[95] = t[107] ^ t[108];
  assign t[96] = t[109] ^ t[108];
  assign t[97] = t[168] ^ t[169];
  assign t[98] = t[170] ^ t[135];
  assign t[99] = t[110] ^ t[111];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [120:0] x;
 output y;

 wire [412:0] t;
  assign t[0] = t[1] ? t[2] : t[133];
  assign t[100] = t[36] ^ t[50];
  assign t[101] = t[36] & t[50];
  assign t[102] = t[59] & t[58];
  assign t[103] = t[112] ^ t[87];
  assign t[104] = t[54] ^ t[113];
  assign t[105] = t[69] ^ t[80];
  assign t[106] = t[171] ^ t[172];
  assign t[107] = t[114] ^ t[115];
  assign t[108] = t[116] ^ t[102];
  assign t[109] = t[117] ^ t[118];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[71] & t[74];
  assign t[111] = t[119] & t[66];
  assign t[112] = t[120] ^ t[121];
  assign t[113] = t[122] ^ t[123];
  assign t[114] = t[124] ^ t[111];
  assign t[115] = t[125] & t[126];
  assign t[116] = t[127] & t[128];
  assign t[117] = t[129] ^ t[121];
  assign t[118] = t[130] & t[122];
  assign t[119] = t[52] ^ t[127];
  assign t[11] = ~(t[17]);
  assign t[120] = t[54] & t[113];
  assign t[121] = t[52] & t[123];
  assign t[122] = t[74] ^ t[67];
  assign t[123] = t[75] ^ t[131];
  assign t[124] = t[66] ^ t[76];
  assign t[125] = t[36] ^ t[130];
  assign t[126] = t[74] ^ t[66];
  assign t[127] = t[77] ^ t[49];
  assign t[128] = t[59] ^ t[131];
  assign t[129] = t[52] ^ t[123];
  assign t[12] = t[136] & t[18];
  assign t[130] = t[67] ^ t[132];
  assign t[131] = t[84] ^ t[49];
  assign t[132] = t[68] ^ t[74];
  assign t[133] = (t[173]);
  assign t[134] = (t[174]);
  assign t[135] = (t[175]);
  assign t[136] = (t[176]);
  assign t[137] = (t[177]);
  assign t[138] = (t[178]);
  assign t[139] = (t[179]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[180]);
  assign t[141] = (t[181]);
  assign t[142] = (t[182]);
  assign t[143] = (t[183]);
  assign t[144] = (t[184]);
  assign t[145] = (t[185]);
  assign t[146] = (t[186]);
  assign t[147] = (t[187]);
  assign t[148] = (t[188]);
  assign t[149] = (t[189]);
  assign t[14] = ~(t[136]);
  assign t[150] = (t[190]);
  assign t[151] = (t[191]);
  assign t[152] = (t[192]);
  assign t[153] = (t[193]);
  assign t[154] = (t[194]);
  assign t[155] = (t[195]);
  assign t[156] = (t[196]);
  assign t[157] = (t[197]);
  assign t[158] = (t[198]);
  assign t[159] = (t[199]);
  assign t[15] = t[137] & t[138];
  assign t[160] = (t[200]);
  assign t[161] = (t[201]);
  assign t[162] = (t[202]);
  assign t[163] = (t[203]);
  assign t[164] = (t[204]);
  assign t[165] = (t[205]);
  assign t[166] = (t[206]);
  assign t[167] = (t[207]);
  assign t[168] = (t[208]);
  assign t[169] = (t[209]);
  assign t[16] = ~(t[21] ^ t[22]);
  assign t[170] = (t[210]);
  assign t[171] = (t[211]);
  assign t[172] = (t[212]);
  assign t[173] = t[213] ^ x[2];
  assign t[174] = t[214] ^ x[6];
  assign t[175] = t[215] ^ x[9];
  assign t[176] = t[216] ^ x[12];
  assign t[177] = t[217] ^ x[15];
  assign t[178] = t[218] ^ x[18];
  assign t[179] = t[219] ^ x[21];
  assign t[17] = ~(t[136] & t[23]);
  assign t[180] = t[220] ^ x[24];
  assign t[181] = t[221] ^ x[27];
  assign t[182] = t[222] ^ x[30];
  assign t[183] = t[223] ^ x[33];
  assign t[184] = t[224] ^ x[36];
  assign t[185] = t[225] ^ x[39];
  assign t[186] = t[226] ^ x[42];
  assign t[187] = t[227] ^ x[45];
  assign t[188] = t[228] ^ x[48];
  assign t[189] = t[229] ^ x[51];
  assign t[18] = t[24] & t[25];
  assign t[190] = t[230] ^ x[54];
  assign t[191] = t[231] ^ x[57];
  assign t[192] = t[232] ^ x[60];
  assign t[193] = t[233] ^ x[63];
  assign t[194] = t[234] ^ x[66];
  assign t[195] = t[235] ^ x[69];
  assign t[196] = t[236] ^ x[72];
  assign t[197] = t[237] ^ x[75];
  assign t[198] = t[238] ^ x[78];
  assign t[199] = t[239] ^ x[81];
  assign t[19] = ~(t[139]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[240] ^ x[84];
  assign t[201] = t[241] ^ x[87];
  assign t[202] = t[242] ^ x[90];
  assign t[203] = t[243] ^ x[93];
  assign t[204] = t[244] ^ x[96];
  assign t[205] = t[245] ^ x[99];
  assign t[206] = t[246] ^ x[102];
  assign t[207] = t[247] ^ x[105];
  assign t[208] = t[248] ^ x[108];
  assign t[209] = t[249] ^ x[111];
  assign t[20] = ~(t[136]);
  assign t[210] = t[250] ^ x[114];
  assign t[211] = t[251] ^ x[117];
  assign t[212] = t[252] ^ x[120];
  assign t[213] = (t[253] & ~t[254]);
  assign t[214] = (t[255] & ~t[256]);
  assign t[215] = (t[257] & ~t[258]);
  assign t[216] = (t[259] & ~t[260]);
  assign t[217] = (t[261] & ~t[262]);
  assign t[218] = (t[263] & ~t[264]);
  assign t[219] = (t[265] & ~t[266]);
  assign t[21] = t[26] ^ t[27];
  assign t[220] = (t[267] & ~t[268]);
  assign t[221] = (t[269] & ~t[270]);
  assign t[222] = (t[271] & ~t[272]);
  assign t[223] = (t[273] & ~t[274]);
  assign t[224] = (t[275] & ~t[276]);
  assign t[225] = (t[277] & ~t[278]);
  assign t[226] = (t[279] & ~t[280]);
  assign t[227] = (t[281] & ~t[282]);
  assign t[228] = (t[283] & ~t[284]);
  assign t[229] = (t[285] & ~t[286]);
  assign t[22] = t[28] ^ t[29];
  assign t[230] = (t[287] & ~t[288]);
  assign t[231] = (t[289] & ~t[290]);
  assign t[232] = (t[291] & ~t[292]);
  assign t[233] = (t[293] & ~t[294]);
  assign t[234] = (t[295] & ~t[296]);
  assign t[235] = (t[297] & ~t[298]);
  assign t[236] = (t[299] & ~t[300]);
  assign t[237] = (t[301] & ~t[302]);
  assign t[238] = (t[303] & ~t[304]);
  assign t[239] = (t[305] & ~t[306]);
  assign t[23] = ~(t[140] | t[30]);
  assign t[240] = (t[307] & ~t[308]);
  assign t[241] = (t[309] & ~t[310]);
  assign t[242] = (t[311] & ~t[312]);
  assign t[243] = (t[313] & ~t[314]);
  assign t[244] = (t[315] & ~t[316]);
  assign t[245] = (t[317] & ~t[318]);
  assign t[246] = (t[319] & ~t[320]);
  assign t[247] = (t[321] & ~t[322]);
  assign t[248] = (t[323] & ~t[324]);
  assign t[249] = (t[325] & ~t[326]);
  assign t[24] = ~(t[31] | t[32]);
  assign t[250] = (t[327] & ~t[328]);
  assign t[251] = (t[329] & ~t[330]);
  assign t[252] = (t[331] & ~t[332]);
  assign t[253] = t[333] ^ x[2];
  assign t[254] = t[334] ^ x[1];
  assign t[255] = t[335] ^ x[6];
  assign t[256] = t[336] ^ x[5];
  assign t[257] = t[337] ^ x[9];
  assign t[258] = t[338] ^ x[8];
  assign t[259] = t[339] ^ x[12];
  assign t[25] = ~(t[33] | t[34]);
  assign t[260] = t[340] ^ x[11];
  assign t[261] = t[341] ^ x[15];
  assign t[262] = t[342] ^ x[14];
  assign t[263] = t[343] ^ x[18];
  assign t[264] = t[344] ^ x[17];
  assign t[265] = t[345] ^ x[21];
  assign t[266] = t[346] ^ x[20];
  assign t[267] = t[347] ^ x[24];
  assign t[268] = t[348] ^ x[23];
  assign t[269] = t[349] ^ x[27];
  assign t[26] = t[35] & t[36];
  assign t[270] = t[350] ^ x[26];
  assign t[271] = t[351] ^ x[30];
  assign t[272] = t[352] ^ x[29];
  assign t[273] = t[353] ^ x[33];
  assign t[274] = t[354] ^ x[32];
  assign t[275] = t[355] ^ x[36];
  assign t[276] = t[356] ^ x[35];
  assign t[277] = t[357] ^ x[39];
  assign t[278] = t[358] ^ x[38];
  assign t[279] = t[359] ^ x[42];
  assign t[27] = t[37] ^ t[38];
  assign t[280] = t[360] ^ x[41];
  assign t[281] = t[361] ^ x[45];
  assign t[282] = t[362] ^ x[44];
  assign t[283] = t[363] ^ x[48];
  assign t[284] = t[364] ^ x[47];
  assign t[285] = t[365] ^ x[51];
  assign t[286] = t[366] ^ x[50];
  assign t[287] = t[367] ^ x[54];
  assign t[288] = t[368] ^ x[53];
  assign t[289] = t[369] ^ x[57];
  assign t[28] = t[39] ^ t[40];
  assign t[290] = t[370] ^ x[56];
  assign t[291] = t[371] ^ x[60];
  assign t[292] = t[372] ^ x[59];
  assign t[293] = t[373] ^ x[63];
  assign t[294] = t[374] ^ x[62];
  assign t[295] = t[375] ^ x[66];
  assign t[296] = t[376] ^ x[65];
  assign t[297] = t[377] ^ x[69];
  assign t[298] = t[378] ^ x[68];
  assign t[299] = t[379] ^ x[72];
  assign t[29] = t[41] ^ t[42];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[380] ^ x[71];
  assign t[301] = t[381] ^ x[75];
  assign t[302] = t[382] ^ x[74];
  assign t[303] = t[383] ^ x[78];
  assign t[304] = t[384] ^ x[77];
  assign t[305] = t[385] ^ x[81];
  assign t[306] = t[386] ^ x[80];
  assign t[307] = t[387] ^ x[84];
  assign t[308] = t[388] ^ x[83];
  assign t[309] = t[389] ^ x[87];
  assign t[30] = ~(t[43] & t[44]);
  assign t[310] = t[390] ^ x[86];
  assign t[311] = t[391] ^ x[90];
  assign t[312] = t[392] ^ x[89];
  assign t[313] = t[393] ^ x[93];
  assign t[314] = t[394] ^ x[92];
  assign t[315] = t[395] ^ x[96];
  assign t[316] = t[396] ^ x[95];
  assign t[317] = t[397] ^ x[99];
  assign t[318] = t[398] ^ x[98];
  assign t[319] = t[399] ^ x[102];
  assign t[31] = ~(t[141] & t[137]);
  assign t[320] = t[400] ^ x[101];
  assign t[321] = t[401] ^ x[105];
  assign t[322] = t[402] ^ x[104];
  assign t[323] = t[403] ^ x[108];
  assign t[324] = t[404] ^ x[107];
  assign t[325] = t[405] ^ x[111];
  assign t[326] = t[406] ^ x[110];
  assign t[327] = t[407] ^ x[114];
  assign t[328] = t[408] ^ x[113];
  assign t[329] = t[409] ^ x[117];
  assign t[32] = ~(t[142] & t[143]);
  assign t[330] = t[410] ^ x[116];
  assign t[331] = t[411] ^ x[120];
  assign t[332] = t[412] ^ x[119];
  assign t[333] = (x[0]);
  assign t[334] = (x[0]);
  assign t[335] = (x[4]);
  assign t[336] = (x[4]);
  assign t[337] = (x[7]);
  assign t[338] = (x[7]);
  assign t[339] = (x[10]);
  assign t[33] = ~(t[23]);
  assign t[340] = (x[10]);
  assign t[341] = (x[13]);
  assign t[342] = (x[13]);
  assign t[343] = (x[16]);
  assign t[344] = (x[16]);
  assign t[345] = (x[19]);
  assign t[346] = (x[19]);
  assign t[347] = (x[22]);
  assign t[348] = (x[22]);
  assign t[349] = (x[25]);
  assign t[34] = ~(t[144] & t[45]);
  assign t[350] = (x[25]);
  assign t[351] = (x[28]);
  assign t[352] = (x[28]);
  assign t[353] = (x[31]);
  assign t[354] = (x[31]);
  assign t[355] = (x[34]);
  assign t[356] = (x[34]);
  assign t[357] = (x[37]);
  assign t[358] = (x[37]);
  assign t[359] = (x[40]);
  assign t[35] = t[46] ^ t[47];
  assign t[360] = (x[40]);
  assign t[361] = (x[43]);
  assign t[362] = (x[43]);
  assign t[363] = (x[46]);
  assign t[364] = (x[46]);
  assign t[365] = (x[49]);
  assign t[366] = (x[49]);
  assign t[367] = (x[52]);
  assign t[368] = (x[52]);
  assign t[369] = (x[55]);
  assign t[36] = t[48] ^ t[49];
  assign t[370] = (x[55]);
  assign t[371] = (x[58]);
  assign t[372] = (x[58]);
  assign t[373] = (x[61]);
  assign t[374] = (x[61]);
  assign t[375] = (x[64]);
  assign t[376] = (x[64]);
  assign t[377] = (x[67]);
  assign t[378] = (x[67]);
  assign t[379] = (x[70]);
  assign t[37] = t[35] & t[50];
  assign t[380] = (x[70]);
  assign t[381] = (x[73]);
  assign t[382] = (x[73]);
  assign t[383] = (x[76]);
  assign t[384] = (x[76]);
  assign t[385] = (x[79]);
  assign t[386] = (x[79]);
  assign t[387] = (x[82]);
  assign t[388] = (x[82]);
  assign t[389] = (x[85]);
  assign t[38] = t[51] & t[52];
  assign t[390] = (x[85]);
  assign t[391] = (x[88]);
  assign t[392] = (x[88]);
  assign t[393] = (x[91]);
  assign t[394] = (x[91]);
  assign t[395] = (x[94]);
  assign t[396] = (x[94]);
  assign t[397] = (x[97]);
  assign t[398] = (x[97]);
  assign t[399] = (x[100]);
  assign t[39] = t[53] & t[54];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[100]);
  assign t[401] = (x[103]);
  assign t[402] = (x[103]);
  assign t[403] = (x[106]);
  assign t[404] = (x[106]);
  assign t[405] = (x[109]);
  assign t[406] = (x[109]);
  assign t[407] = (x[112]);
  assign t[408] = (x[112]);
  assign t[409] = (x[115]);
  assign t[40] = t[55] ^ t[56];
  assign t[410] = (x[115]);
  assign t[411] = (x[118]);
  assign t[412] = (x[118]);
  assign t[41] = t[57] & t[58];
  assign t[42] = t[57] & t[59];
  assign t[43] = ~(t[145] | t[146]);
  assign t[44] = ~(t[147] | t[148]);
  assign t[45] = ~(t[149]);
  assign t[46] = t[60] ^ t[61];
  assign t[47] = t[62] ^ t[63];
  assign t[48] = t[13] ? t[150] : t[64];
  assign t[49] = t[13] ? t[151] : t[65];
  assign t[4] = ~(t[8]);
  assign t[50] = t[66] ^ t[67];
  assign t[51] = t[53] ^ t[46];
  assign t[52] = t[48] ^ t[68];
  assign t[53] = t[69] ^ t[70];
  assign t[54] = t[59] ^ t[71];
  assign t[55] = t[72] & t[66];
  assign t[56] = t[73] & t[74];
  assign t[57] = t[53] ^ t[73];
  assign t[58] = t[75] ^ t[76];
  assign t[59] = t[48] ^ t[77];
  assign t[5] = t[9] ? t[134] : x[3];
  assign t[60] = t[78] & t[79];
  assign t[61] = t[78] ^ t[80];
  assign t[62] = t[81] & t[82];
  assign t[63] = t[81] ^ t[80];
  assign t[64] = t[152] ^ t[153];
  assign t[65] = t[154] ^ t[155];
  assign t[66] = t[59] ^ t[75];
  assign t[67] = t[83] ^ t[84];
  assign t[68] = t[13] ? t[156] : t[85];
  assign t[69] = t[86] ^ t[87];
  assign t[6] = ~(t[10] ^ t[135]);
  assign t[70] = t[88] & t[78];
  assign t[71] = t[67] ^ t[89];
  assign t[72] = t[73] ^ t[47];
  assign t[73] = t[90] ^ t[91];
  assign t[74] = t[13] ? t[157] : t[92];
  assign t[75] = t[93] ^ t[68];
  assign t[76] = t[83] ^ t[49];
  assign t[77] = t[13] ? t[158] : t[94];
  assign t[78] = t[95] ^ t[69];
  assign t[79] = t[95] & t[90];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[96] & t[95];
  assign t[81] = t[96] ^ t[90];
  assign t[82] = t[69] & t[96];
  assign t[83] = t[13] ? t[159] : t[97];
  assign t[84] = t[13] ? t[160] : t[98];
  assign t[85] = t[161] ^ t[162];
  assign t[86] = t[99] ^ t[100];
  assign t[87] = t[101] ^ t[102];
  assign t[88] = t[90] ^ t[80];
  assign t[89] = t[77] ^ t[74];
  assign t[8] = ~(t[13]);
  assign t[90] = t[103] ^ t[104];
  assign t[91] = t[105] & t[81];
  assign t[92] = t[163] ^ t[164];
  assign t[93] = t[13] ? t[165] : t[106];
  assign t[94] = t[166] ^ t[167];
  assign t[95] = t[107] ^ t[108];
  assign t[96] = t[109] ^ t[108];
  assign t[97] = t[168] ^ t[169];
  assign t[98] = t[170] ^ t[135];
  assign t[99] = t[110] ^ t[111];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [123:0] x;
 output y;

 wire [421:0] t;
  assign t[0] = t[1] ? t[2] : t[135];
  assign t[100] = t[121] ^ t[122];
  assign t[101] = t[167] ^ t[137];
  assign t[102] = t[168] ^ t[169];
  assign t[103] = t[170] ^ t[171];
  assign t[104] = t[172] ^ t[173];
  assign t[105] = t[79] ^ t[64];
  assign t[106] = t[81] ^ t[80];
  assign t[107] = t[80] ^ t[64];
  assign t[108] = t[106] & t[123];
  assign t[109] = t[106] ^ t[64];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[174] ^ t[175];
  assign t[111] = t[124] ^ t[125];
  assign t[112] = t[51] & t[126];
  assign t[113] = t[55] & t[61];
  assign t[114] = t[53] & t[60];
  assign t[115] = t[127] ^ t[125];
  assign t[116] = t[53] ^ t[128];
  assign t[117] = t[126] ^ t[129];
  assign t[118] = t[130] ^ t[131];
  assign t[119] = t[50] ^ t[132];
  assign t[11] = ~(t[17]);
  assign t[120] = t[50] & t[132];
  assign t[121] = t[133] ^ t[131];
  assign t[122] = t[38] & t[74];
  assign t[123] = t[81] & t[79];
  assign t[124] = t[93] ^ t[129];
  assign t[125] = t[93] & t[129];
  assign t[126] = t[87] ^ t[67];
  assign t[127] = t[116] & t[117];
  assign t[128] = t[67] ^ t[134];
  assign t[129] = t[73] ^ t[77];
  assign t[12] = t[138] & t[18];
  assign t[130] = t[128] & t[87];
  assign t[131] = t[75] & t[57];
  assign t[132] = t[57] ^ t[67];
  assign t[133] = t[57] ^ t[76];
  assign t[134] = t[71] ^ t[87];
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = ~(t[138]);
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = (t[194]);
  assign t[154] = (t[195]);
  assign t[155] = (t[196]);
  assign t[156] = (t[197]);
  assign t[157] = (t[198]);
  assign t[158] = (t[199]);
  assign t[159] = (t[200]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[201]);
  assign t[161] = (t[202]);
  assign t[162] = (t[203]);
  assign t[163] = (t[204]);
  assign t[164] = (t[205]);
  assign t[165] = (t[206]);
  assign t[166] = (t[207]);
  assign t[167] = (t[208]);
  assign t[168] = (t[209]);
  assign t[169] = (t[210]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (t[211]);
  assign t[171] = (t[212]);
  assign t[172] = (t[213]);
  assign t[173] = (t[214]);
  assign t[174] = (t[215]);
  assign t[175] = (t[216]);
  assign t[176] = t[217] ^ x[2];
  assign t[177] = t[218] ^ x[6];
  assign t[178] = t[219] ^ x[9];
  assign t[179] = t[220] ^ x[12];
  assign t[17] = ~(t[138] & t[25]);
  assign t[180] = t[221] ^ x[15];
  assign t[181] = t[222] ^ x[18];
  assign t[182] = t[223] ^ x[21];
  assign t[183] = t[224] ^ x[24];
  assign t[184] = t[225] ^ x[27];
  assign t[185] = t[226] ^ x[30];
  assign t[186] = t[227] ^ x[33];
  assign t[187] = t[228] ^ x[36];
  assign t[188] = t[229] ^ x[39];
  assign t[189] = t[230] ^ x[42];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[231] ^ x[45];
  assign t[191] = t[232] ^ x[48];
  assign t[192] = t[233] ^ x[51];
  assign t[193] = t[234] ^ x[54];
  assign t[194] = t[235] ^ x[57];
  assign t[195] = t[236] ^ x[60];
  assign t[196] = t[237] ^ x[63];
  assign t[197] = t[238] ^ x[66];
  assign t[198] = t[239] ^ x[69];
  assign t[199] = t[240] ^ x[72];
  assign t[19] = ~(t[139]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[241] ^ x[75];
  assign t[201] = t[242] ^ x[78];
  assign t[202] = t[243] ^ x[81];
  assign t[203] = t[244] ^ x[84];
  assign t[204] = t[245] ^ x[87];
  assign t[205] = t[246] ^ x[90];
  assign t[206] = t[247] ^ x[93];
  assign t[207] = t[248] ^ x[96];
  assign t[208] = t[249] ^ x[99];
  assign t[209] = t[250] ^ x[102];
  assign t[20] = ~(t[138]);
  assign t[210] = t[251] ^ x[105];
  assign t[211] = t[252] ^ x[108];
  assign t[212] = t[253] ^ x[111];
  assign t[213] = t[254] ^ x[114];
  assign t[214] = t[255] ^ x[117];
  assign t[215] = t[256] ^ x[120];
  assign t[216] = t[257] ^ x[123];
  assign t[217] = (t[258] & ~t[259]);
  assign t[218] = (t[260] & ~t[261]);
  assign t[219] = (t[262] & ~t[263]);
  assign t[21] = ~(t[140]);
  assign t[220] = (t[264] & ~t[265]);
  assign t[221] = (t[266] & ~t[267]);
  assign t[222] = (t[268] & ~t[269]);
  assign t[223] = (t[270] & ~t[271]);
  assign t[224] = (t[272] & ~t[273]);
  assign t[225] = (t[274] & ~t[275]);
  assign t[226] = (t[276] & ~t[277]);
  assign t[227] = (t[278] & ~t[279]);
  assign t[228] = (t[280] & ~t[281]);
  assign t[229] = (t[282] & ~t[283]);
  assign t[22] = ~(t[141]);
  assign t[230] = (t[284] & ~t[285]);
  assign t[231] = (t[286] & ~t[287]);
  assign t[232] = (t[288] & ~t[289]);
  assign t[233] = (t[290] & ~t[291]);
  assign t[234] = (t[292] & ~t[293]);
  assign t[235] = (t[294] & ~t[295]);
  assign t[236] = (t[296] & ~t[297]);
  assign t[237] = (t[298] & ~t[299]);
  assign t[238] = (t[300] & ~t[301]);
  assign t[239] = (t[302] & ~t[303]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[304] & ~t[305]);
  assign t[241] = (t[306] & ~t[307]);
  assign t[242] = (t[308] & ~t[309]);
  assign t[243] = (t[310] & ~t[311]);
  assign t[244] = (t[312] & ~t[313]);
  assign t[245] = (t[314] & ~t[315]);
  assign t[246] = (t[316] & ~t[317]);
  assign t[247] = (t[318] & ~t[319]);
  assign t[248] = (t[320] & ~t[321]);
  assign t[249] = (t[322] & ~t[323]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[324] & ~t[325]);
  assign t[251] = (t[326] & ~t[327]);
  assign t[252] = (t[328] & ~t[329]);
  assign t[253] = (t[330] & ~t[331]);
  assign t[254] = (t[332] & ~t[333]);
  assign t[255] = (t[334] & ~t[335]);
  assign t[256] = (t[336] & ~t[337]);
  assign t[257] = (t[338] & ~t[339]);
  assign t[258] = t[340] ^ x[2];
  assign t[259] = t[341] ^ x[1];
  assign t[25] = ~(t[142] | t[32]);
  assign t[260] = t[342] ^ x[6];
  assign t[261] = t[343] ^ x[5];
  assign t[262] = t[344] ^ x[9];
  assign t[263] = t[345] ^ x[8];
  assign t[264] = t[346] ^ x[12];
  assign t[265] = t[347] ^ x[11];
  assign t[266] = t[348] ^ x[15];
  assign t[267] = t[349] ^ x[14];
  assign t[268] = t[350] ^ x[18];
  assign t[269] = t[351] ^ x[17];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[352] ^ x[21];
  assign t[271] = t[353] ^ x[20];
  assign t[272] = t[354] ^ x[24];
  assign t[273] = t[355] ^ x[23];
  assign t[274] = t[356] ^ x[27];
  assign t[275] = t[357] ^ x[26];
  assign t[276] = t[358] ^ x[30];
  assign t[277] = t[359] ^ x[29];
  assign t[278] = t[360] ^ x[33];
  assign t[279] = t[361] ^ x[32];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[362] ^ x[36];
  assign t[281] = t[363] ^ x[35];
  assign t[282] = t[364] ^ x[39];
  assign t[283] = t[365] ^ x[38];
  assign t[284] = t[366] ^ x[42];
  assign t[285] = t[367] ^ x[41];
  assign t[286] = t[368] ^ x[45];
  assign t[287] = t[369] ^ x[44];
  assign t[288] = t[370] ^ x[48];
  assign t[289] = t[371] ^ x[47];
  assign t[28] = t[37] & t[38];
  assign t[290] = t[372] ^ x[51];
  assign t[291] = t[373] ^ x[50];
  assign t[292] = t[374] ^ x[54];
  assign t[293] = t[375] ^ x[53];
  assign t[294] = t[376] ^ x[57];
  assign t[295] = t[377] ^ x[56];
  assign t[296] = t[378] ^ x[60];
  assign t[297] = t[379] ^ x[59];
  assign t[298] = t[380] ^ x[63];
  assign t[299] = t[381] ^ x[62];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[66];
  assign t[301] = t[383] ^ x[65];
  assign t[302] = t[384] ^ x[69];
  assign t[303] = t[385] ^ x[68];
  assign t[304] = t[386] ^ x[72];
  assign t[305] = t[387] ^ x[71];
  assign t[306] = t[388] ^ x[75];
  assign t[307] = t[389] ^ x[74];
  assign t[308] = t[390] ^ x[78];
  assign t[309] = t[391] ^ x[77];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[392] ^ x[81];
  assign t[311] = t[393] ^ x[80];
  assign t[312] = t[394] ^ x[84];
  assign t[313] = t[395] ^ x[83];
  assign t[314] = t[396] ^ x[87];
  assign t[315] = t[397] ^ x[86];
  assign t[316] = t[398] ^ x[90];
  assign t[317] = t[399] ^ x[89];
  assign t[318] = t[400] ^ x[93];
  assign t[319] = t[401] ^ x[92];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[402] ^ x[96];
  assign t[321] = t[403] ^ x[95];
  assign t[322] = t[404] ^ x[99];
  assign t[323] = t[405] ^ x[98];
  assign t[324] = t[406] ^ x[102];
  assign t[325] = t[407] ^ x[101];
  assign t[326] = t[408] ^ x[105];
  assign t[327] = t[409] ^ x[104];
  assign t[328] = t[410] ^ x[108];
  assign t[329] = t[411] ^ x[107];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[412] ^ x[111];
  assign t[331] = t[413] ^ x[110];
  assign t[332] = t[414] ^ x[114];
  assign t[333] = t[415] ^ x[113];
  assign t[334] = t[416] ^ x[117];
  assign t[335] = t[417] ^ x[116];
  assign t[336] = t[418] ^ x[120];
  assign t[337] = t[419] ^ x[119];
  assign t[338] = t[420] ^ x[123];
  assign t[339] = t[421] ^ x[122];
  assign t[33] = ~(t[143] & t[144]);
  assign t[340] = (x[0]);
  assign t[341] = (x[0]);
  assign t[342] = (x[4]);
  assign t[343] = (x[4]);
  assign t[344] = (x[7]);
  assign t[345] = (x[7]);
  assign t[346] = (x[10]);
  assign t[347] = (x[10]);
  assign t[348] = (x[13]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[145] & t[146]);
  assign t[350] = (x[16]);
  assign t[351] = (x[16]);
  assign t[352] = (x[19]);
  assign t[353] = (x[19]);
  assign t[354] = (x[22]);
  assign t[355] = (x[22]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[28]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[31]);
  assign t[361] = (x[31]);
  assign t[362] = (x[34]);
  assign t[363] = (x[34]);
  assign t[364] = (x[37]);
  assign t[365] = (x[37]);
  assign t[366] = (x[40]);
  assign t[367] = (x[40]);
  assign t[368] = (x[43]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[147] & t[47]);
  assign t[370] = (x[46]);
  assign t[371] = (x[46]);
  assign t[372] = (x[49]);
  assign t[373] = (x[49]);
  assign t[374] = (x[52]);
  assign t[375] = (x[52]);
  assign t[376] = (x[55]);
  assign t[377] = (x[55]);
  assign t[378] = (x[58]);
  assign t[379] = (x[58]);
  assign t[37] = t[48] ^ t[49];
  assign t[380] = (x[61]);
  assign t[381] = (x[61]);
  assign t[382] = (x[64]);
  assign t[383] = (x[64]);
  assign t[384] = (x[67]);
  assign t[385] = (x[67]);
  assign t[386] = (x[70]);
  assign t[387] = (x[70]);
  assign t[388] = (x[73]);
  assign t[389] = (x[73]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[76]);
  assign t[391] = (x[76]);
  assign t[392] = (x[79]);
  assign t[393] = (x[79]);
  assign t[394] = (x[82]);
  assign t[395] = (x[82]);
  assign t[396] = (x[85]);
  assign t[397] = (x[85]);
  assign t[398] = (x[88]);
  assign t[399] = (x[88]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[91]);
  assign t[401] = (x[91]);
  assign t[402] = (x[94]);
  assign t[403] = (x[94]);
  assign t[404] = (x[97]);
  assign t[405] = (x[97]);
  assign t[406] = (x[100]);
  assign t[407] = (x[100]);
  assign t[408] = (x[103]);
  assign t[409] = (x[103]);
  assign t[40] = t[54] & t[55];
  assign t[410] = (x[106]);
  assign t[411] = (x[106]);
  assign t[412] = (x[109]);
  assign t[413] = (x[109]);
  assign t[414] = (x[112]);
  assign t[415] = (x[112]);
  assign t[416] = (x[115]);
  assign t[417] = (x[115]);
  assign t[418] = (x[118]);
  assign t[419] = (x[118]);
  assign t[41] = t[56] & t[57];
  assign t[420] = (x[121]);
  assign t[421] = (x[121]);
  assign t[42] = t[58] ^ t[59];
  assign t[43] = t[52] & t[60];
  assign t[44] = t[54] & t[61];
  assign t[45] = ~(t[148] | t[149]);
  assign t[46] = ~(t[150] | t[151]);
  assign t[47] = ~(t[152]);
  assign t[48] = t[62] & t[63];
  assign t[49] = t[62] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[65] ^ t[66];
  assign t[51] = t[67] ^ t[68];
  assign t[52] = t[69] ^ t[70];
  assign t[53] = t[65] ^ t[71];
  assign t[54] = t[52] ^ t[72];
  assign t[55] = t[71] ^ t[66];
  assign t[56] = t[70] ^ t[37];
  assign t[57] = t[53] ^ t[73];
  assign t[58] = t[37] & t[74];
  assign t[59] = t[56] & t[75];
  assign t[5] = t[9] ? t[136] : x[3];
  assign t[60] = t[73] ^ t[76];
  assign t[61] = t[53] ^ t[77];
  assign t[62] = t[78] ^ t[79];
  assign t[63] = t[80] & t[78];
  assign t[64] = t[78] & t[81];
  assign t[65] = t[13] ? t[153] : t[82];
  assign t[66] = t[13] ? t[154] : t[83];
  assign t[67] = t[84] ^ t[85];
  assign t[68] = t[86] ^ t[87];
  assign t[69] = t[80] ^ t[88];
  assign t[6] = ~(t[10] ^ t[137]);
  assign t[70] = t[79] ^ t[89];
  assign t[71] = t[13] ? t[155] : t[90];
  assign t[72] = t[91] ^ t[37];
  assign t[73] = t[92] ^ t[86];
  assign t[74] = t[87] ^ t[57];
  assign t[75] = t[93] ^ t[55];
  assign t[76] = t[84] ^ t[66];
  assign t[77] = t[85] ^ t[66];
  assign t[78] = t[94] ^ t[95];
  assign t[79] = t[96] ^ t[97];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[98] ^ t[99];
  assign t[81] = t[100] ^ t[95];
  assign t[82] = t[156] ^ t[157];
  assign t[83] = t[158] ^ t[159];
  assign t[84] = t[13] ? t[160] : t[101];
  assign t[85] = t[13] ? t[161] : t[102];
  assign t[86] = t[13] ? t[162] : t[103];
  assign t[87] = t[13] ? t[163] : t[104];
  assign t[88] = t[105] & t[106];
  assign t[89] = t[107] & t[62];
  assign t[8] = ~(t[13]);
  assign t[90] = t[164] ^ t[165];
  assign t[91] = t[108] ^ t[109];
  assign t[92] = t[13] ? t[166] : t[110];
  assign t[93] = t[65] ^ t[86];
  assign t[94] = t[111] ^ t[112];
  assign t[95] = t[113] ^ t[114];
  assign t[96] = t[115] ^ t[99];
  assign t[97] = t[116] ^ t[117];
  assign t[98] = t[118] ^ t[119];
  assign t[99] = t[120] ^ t[114];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [123:0] x;
 output y;

 wire [421:0] t;
  assign t[0] = t[1] ? t[2] : t[135];
  assign t[100] = t[121] ^ t[122];
  assign t[101] = t[167] ^ t[137];
  assign t[102] = t[168] ^ t[169];
  assign t[103] = t[170] ^ t[171];
  assign t[104] = t[172] ^ t[173];
  assign t[105] = t[79] ^ t[64];
  assign t[106] = t[81] ^ t[80];
  assign t[107] = t[80] ^ t[64];
  assign t[108] = t[106] & t[123];
  assign t[109] = t[106] ^ t[64];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[174] ^ t[175];
  assign t[111] = t[124] ^ t[125];
  assign t[112] = t[51] & t[126];
  assign t[113] = t[55] & t[61];
  assign t[114] = t[53] & t[60];
  assign t[115] = t[127] ^ t[125];
  assign t[116] = t[53] ^ t[128];
  assign t[117] = t[126] ^ t[129];
  assign t[118] = t[130] ^ t[131];
  assign t[119] = t[50] ^ t[132];
  assign t[11] = ~(t[17]);
  assign t[120] = t[50] & t[132];
  assign t[121] = t[133] ^ t[131];
  assign t[122] = t[38] & t[74];
  assign t[123] = t[81] & t[79];
  assign t[124] = t[93] ^ t[129];
  assign t[125] = t[93] & t[129];
  assign t[126] = t[87] ^ t[67];
  assign t[127] = t[116] & t[117];
  assign t[128] = t[67] ^ t[134];
  assign t[129] = t[73] ^ t[77];
  assign t[12] = t[138] & t[18];
  assign t[130] = t[128] & t[87];
  assign t[131] = t[75] & t[57];
  assign t[132] = t[57] ^ t[67];
  assign t[133] = t[57] ^ t[76];
  assign t[134] = t[71] ^ t[87];
  assign t[135] = (t[176]);
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = ~(t[138]);
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = (t[194]);
  assign t[154] = (t[195]);
  assign t[155] = (t[196]);
  assign t[156] = (t[197]);
  assign t[157] = (t[198]);
  assign t[158] = (t[199]);
  assign t[159] = (t[200]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[201]);
  assign t[161] = (t[202]);
  assign t[162] = (t[203]);
  assign t[163] = (t[204]);
  assign t[164] = (t[205]);
  assign t[165] = (t[206]);
  assign t[166] = (t[207]);
  assign t[167] = (t[208]);
  assign t[168] = (t[209]);
  assign t[169] = (t[210]);
  assign t[16] = ~(t[23] ^ t[24]);
  assign t[170] = (t[211]);
  assign t[171] = (t[212]);
  assign t[172] = (t[213]);
  assign t[173] = (t[214]);
  assign t[174] = (t[215]);
  assign t[175] = (t[216]);
  assign t[176] = t[217] ^ x[2];
  assign t[177] = t[218] ^ x[6];
  assign t[178] = t[219] ^ x[9];
  assign t[179] = t[220] ^ x[12];
  assign t[17] = ~(t[138] & t[25]);
  assign t[180] = t[221] ^ x[15];
  assign t[181] = t[222] ^ x[18];
  assign t[182] = t[223] ^ x[21];
  assign t[183] = t[224] ^ x[24];
  assign t[184] = t[225] ^ x[27];
  assign t[185] = t[226] ^ x[30];
  assign t[186] = t[227] ^ x[33];
  assign t[187] = t[228] ^ x[36];
  assign t[188] = t[229] ^ x[39];
  assign t[189] = t[230] ^ x[42];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[231] ^ x[45];
  assign t[191] = t[232] ^ x[48];
  assign t[192] = t[233] ^ x[51];
  assign t[193] = t[234] ^ x[54];
  assign t[194] = t[235] ^ x[57];
  assign t[195] = t[236] ^ x[60];
  assign t[196] = t[237] ^ x[63];
  assign t[197] = t[238] ^ x[66];
  assign t[198] = t[239] ^ x[69];
  assign t[199] = t[240] ^ x[72];
  assign t[19] = ~(t[139]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[241] ^ x[75];
  assign t[201] = t[242] ^ x[78];
  assign t[202] = t[243] ^ x[81];
  assign t[203] = t[244] ^ x[84];
  assign t[204] = t[245] ^ x[87];
  assign t[205] = t[246] ^ x[90];
  assign t[206] = t[247] ^ x[93];
  assign t[207] = t[248] ^ x[96];
  assign t[208] = t[249] ^ x[99];
  assign t[209] = t[250] ^ x[102];
  assign t[20] = ~(t[138]);
  assign t[210] = t[251] ^ x[105];
  assign t[211] = t[252] ^ x[108];
  assign t[212] = t[253] ^ x[111];
  assign t[213] = t[254] ^ x[114];
  assign t[214] = t[255] ^ x[117];
  assign t[215] = t[256] ^ x[120];
  assign t[216] = t[257] ^ x[123];
  assign t[217] = (t[258] & ~t[259]);
  assign t[218] = (t[260] & ~t[261]);
  assign t[219] = (t[262] & ~t[263]);
  assign t[21] = ~(t[140]);
  assign t[220] = (t[264] & ~t[265]);
  assign t[221] = (t[266] & ~t[267]);
  assign t[222] = (t[268] & ~t[269]);
  assign t[223] = (t[270] & ~t[271]);
  assign t[224] = (t[272] & ~t[273]);
  assign t[225] = (t[274] & ~t[275]);
  assign t[226] = (t[276] & ~t[277]);
  assign t[227] = (t[278] & ~t[279]);
  assign t[228] = (t[280] & ~t[281]);
  assign t[229] = (t[282] & ~t[283]);
  assign t[22] = ~(t[141]);
  assign t[230] = (t[284] & ~t[285]);
  assign t[231] = (t[286] & ~t[287]);
  assign t[232] = (t[288] & ~t[289]);
  assign t[233] = (t[290] & ~t[291]);
  assign t[234] = (t[292] & ~t[293]);
  assign t[235] = (t[294] & ~t[295]);
  assign t[236] = (t[296] & ~t[297]);
  assign t[237] = (t[298] & ~t[299]);
  assign t[238] = (t[300] & ~t[301]);
  assign t[239] = (t[302] & ~t[303]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[304] & ~t[305]);
  assign t[241] = (t[306] & ~t[307]);
  assign t[242] = (t[308] & ~t[309]);
  assign t[243] = (t[310] & ~t[311]);
  assign t[244] = (t[312] & ~t[313]);
  assign t[245] = (t[314] & ~t[315]);
  assign t[246] = (t[316] & ~t[317]);
  assign t[247] = (t[318] & ~t[319]);
  assign t[248] = (t[320] & ~t[321]);
  assign t[249] = (t[322] & ~t[323]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[324] & ~t[325]);
  assign t[251] = (t[326] & ~t[327]);
  assign t[252] = (t[328] & ~t[329]);
  assign t[253] = (t[330] & ~t[331]);
  assign t[254] = (t[332] & ~t[333]);
  assign t[255] = (t[334] & ~t[335]);
  assign t[256] = (t[336] & ~t[337]);
  assign t[257] = (t[338] & ~t[339]);
  assign t[258] = t[340] ^ x[2];
  assign t[259] = t[341] ^ x[1];
  assign t[25] = ~(t[142] | t[32]);
  assign t[260] = t[342] ^ x[6];
  assign t[261] = t[343] ^ x[5];
  assign t[262] = t[344] ^ x[9];
  assign t[263] = t[345] ^ x[8];
  assign t[264] = t[346] ^ x[12];
  assign t[265] = t[347] ^ x[11];
  assign t[266] = t[348] ^ x[15];
  assign t[267] = t[349] ^ x[14];
  assign t[268] = t[350] ^ x[18];
  assign t[269] = t[351] ^ x[17];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[352] ^ x[21];
  assign t[271] = t[353] ^ x[20];
  assign t[272] = t[354] ^ x[24];
  assign t[273] = t[355] ^ x[23];
  assign t[274] = t[356] ^ x[27];
  assign t[275] = t[357] ^ x[26];
  assign t[276] = t[358] ^ x[30];
  assign t[277] = t[359] ^ x[29];
  assign t[278] = t[360] ^ x[33];
  assign t[279] = t[361] ^ x[32];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[362] ^ x[36];
  assign t[281] = t[363] ^ x[35];
  assign t[282] = t[364] ^ x[39];
  assign t[283] = t[365] ^ x[38];
  assign t[284] = t[366] ^ x[42];
  assign t[285] = t[367] ^ x[41];
  assign t[286] = t[368] ^ x[45];
  assign t[287] = t[369] ^ x[44];
  assign t[288] = t[370] ^ x[48];
  assign t[289] = t[371] ^ x[47];
  assign t[28] = t[37] & t[38];
  assign t[290] = t[372] ^ x[51];
  assign t[291] = t[373] ^ x[50];
  assign t[292] = t[374] ^ x[54];
  assign t[293] = t[375] ^ x[53];
  assign t[294] = t[376] ^ x[57];
  assign t[295] = t[377] ^ x[56];
  assign t[296] = t[378] ^ x[60];
  assign t[297] = t[379] ^ x[59];
  assign t[298] = t[380] ^ x[63];
  assign t[299] = t[381] ^ x[62];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[66];
  assign t[301] = t[383] ^ x[65];
  assign t[302] = t[384] ^ x[69];
  assign t[303] = t[385] ^ x[68];
  assign t[304] = t[386] ^ x[72];
  assign t[305] = t[387] ^ x[71];
  assign t[306] = t[388] ^ x[75];
  assign t[307] = t[389] ^ x[74];
  assign t[308] = t[390] ^ x[78];
  assign t[309] = t[391] ^ x[77];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[392] ^ x[81];
  assign t[311] = t[393] ^ x[80];
  assign t[312] = t[394] ^ x[84];
  assign t[313] = t[395] ^ x[83];
  assign t[314] = t[396] ^ x[87];
  assign t[315] = t[397] ^ x[86];
  assign t[316] = t[398] ^ x[90];
  assign t[317] = t[399] ^ x[89];
  assign t[318] = t[400] ^ x[93];
  assign t[319] = t[401] ^ x[92];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[402] ^ x[96];
  assign t[321] = t[403] ^ x[95];
  assign t[322] = t[404] ^ x[99];
  assign t[323] = t[405] ^ x[98];
  assign t[324] = t[406] ^ x[102];
  assign t[325] = t[407] ^ x[101];
  assign t[326] = t[408] ^ x[105];
  assign t[327] = t[409] ^ x[104];
  assign t[328] = t[410] ^ x[108];
  assign t[329] = t[411] ^ x[107];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[412] ^ x[111];
  assign t[331] = t[413] ^ x[110];
  assign t[332] = t[414] ^ x[114];
  assign t[333] = t[415] ^ x[113];
  assign t[334] = t[416] ^ x[117];
  assign t[335] = t[417] ^ x[116];
  assign t[336] = t[418] ^ x[120];
  assign t[337] = t[419] ^ x[119];
  assign t[338] = t[420] ^ x[123];
  assign t[339] = t[421] ^ x[122];
  assign t[33] = ~(t[143] & t[144]);
  assign t[340] = (x[0]);
  assign t[341] = (x[0]);
  assign t[342] = (x[4]);
  assign t[343] = (x[4]);
  assign t[344] = (x[7]);
  assign t[345] = (x[7]);
  assign t[346] = (x[10]);
  assign t[347] = (x[10]);
  assign t[348] = (x[13]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[145] & t[146]);
  assign t[350] = (x[16]);
  assign t[351] = (x[16]);
  assign t[352] = (x[19]);
  assign t[353] = (x[19]);
  assign t[354] = (x[22]);
  assign t[355] = (x[22]);
  assign t[356] = (x[25]);
  assign t[357] = (x[25]);
  assign t[358] = (x[28]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[31]);
  assign t[361] = (x[31]);
  assign t[362] = (x[34]);
  assign t[363] = (x[34]);
  assign t[364] = (x[37]);
  assign t[365] = (x[37]);
  assign t[366] = (x[40]);
  assign t[367] = (x[40]);
  assign t[368] = (x[43]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[147] & t[47]);
  assign t[370] = (x[46]);
  assign t[371] = (x[46]);
  assign t[372] = (x[49]);
  assign t[373] = (x[49]);
  assign t[374] = (x[52]);
  assign t[375] = (x[52]);
  assign t[376] = (x[55]);
  assign t[377] = (x[55]);
  assign t[378] = (x[58]);
  assign t[379] = (x[58]);
  assign t[37] = t[48] ^ t[49];
  assign t[380] = (x[61]);
  assign t[381] = (x[61]);
  assign t[382] = (x[64]);
  assign t[383] = (x[64]);
  assign t[384] = (x[67]);
  assign t[385] = (x[67]);
  assign t[386] = (x[70]);
  assign t[387] = (x[70]);
  assign t[388] = (x[73]);
  assign t[389] = (x[73]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[76]);
  assign t[391] = (x[76]);
  assign t[392] = (x[79]);
  assign t[393] = (x[79]);
  assign t[394] = (x[82]);
  assign t[395] = (x[82]);
  assign t[396] = (x[85]);
  assign t[397] = (x[85]);
  assign t[398] = (x[88]);
  assign t[399] = (x[88]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[91]);
  assign t[401] = (x[91]);
  assign t[402] = (x[94]);
  assign t[403] = (x[94]);
  assign t[404] = (x[97]);
  assign t[405] = (x[97]);
  assign t[406] = (x[100]);
  assign t[407] = (x[100]);
  assign t[408] = (x[103]);
  assign t[409] = (x[103]);
  assign t[40] = t[54] & t[55];
  assign t[410] = (x[106]);
  assign t[411] = (x[106]);
  assign t[412] = (x[109]);
  assign t[413] = (x[109]);
  assign t[414] = (x[112]);
  assign t[415] = (x[112]);
  assign t[416] = (x[115]);
  assign t[417] = (x[115]);
  assign t[418] = (x[118]);
  assign t[419] = (x[118]);
  assign t[41] = t[56] & t[57];
  assign t[420] = (x[121]);
  assign t[421] = (x[121]);
  assign t[42] = t[58] ^ t[59];
  assign t[43] = t[52] & t[60];
  assign t[44] = t[54] & t[61];
  assign t[45] = ~(t[148] | t[149]);
  assign t[46] = ~(t[150] | t[151]);
  assign t[47] = ~(t[152]);
  assign t[48] = t[62] & t[63];
  assign t[49] = t[62] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[65] ^ t[66];
  assign t[51] = t[67] ^ t[68];
  assign t[52] = t[69] ^ t[70];
  assign t[53] = t[65] ^ t[71];
  assign t[54] = t[52] ^ t[72];
  assign t[55] = t[71] ^ t[66];
  assign t[56] = t[70] ^ t[37];
  assign t[57] = t[53] ^ t[73];
  assign t[58] = t[37] & t[74];
  assign t[59] = t[56] & t[75];
  assign t[5] = t[9] ? t[136] : x[3];
  assign t[60] = t[73] ^ t[76];
  assign t[61] = t[53] ^ t[77];
  assign t[62] = t[78] ^ t[79];
  assign t[63] = t[80] & t[78];
  assign t[64] = t[78] & t[81];
  assign t[65] = t[13] ? t[153] : t[82];
  assign t[66] = t[13] ? t[154] : t[83];
  assign t[67] = t[84] ^ t[85];
  assign t[68] = t[86] ^ t[87];
  assign t[69] = t[80] ^ t[88];
  assign t[6] = ~(t[10] ^ t[137]);
  assign t[70] = t[79] ^ t[89];
  assign t[71] = t[13] ? t[155] : t[90];
  assign t[72] = t[91] ^ t[37];
  assign t[73] = t[92] ^ t[86];
  assign t[74] = t[87] ^ t[57];
  assign t[75] = t[93] ^ t[55];
  assign t[76] = t[84] ^ t[66];
  assign t[77] = t[85] ^ t[66];
  assign t[78] = t[94] ^ t[95];
  assign t[79] = t[96] ^ t[97];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[98] ^ t[99];
  assign t[81] = t[100] ^ t[95];
  assign t[82] = t[156] ^ t[157];
  assign t[83] = t[158] ^ t[159];
  assign t[84] = t[13] ? t[160] : t[101];
  assign t[85] = t[13] ? t[161] : t[102];
  assign t[86] = t[13] ? t[162] : t[103];
  assign t[87] = t[13] ? t[163] : t[104];
  assign t[88] = t[105] & t[106];
  assign t[89] = t[107] & t[62];
  assign t[8] = ~(t[13]);
  assign t[90] = t[164] ^ t[165];
  assign t[91] = t[108] ^ t[109];
  assign t[92] = t[13] ? t[166] : t[110];
  assign t[93] = t[65] ^ t[86];
  assign t[94] = t[111] ^ t[112];
  assign t[95] = t[113] ^ t[114];
  assign t[96] = t[115] ^ t[99];
  assign t[97] = t[116] ^ t[117];
  assign t[98] = t[118] ^ t[119];
  assign t[99] = t[120] ^ t[114];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind246(x, y);
 input [123:0] x;
 output y;

 wire [422:0] t;
  assign t[0] = t[1] ? t[2] : t[136];
  assign t[100] = t[116] & t[112];
  assign t[101] = t[74] & t[116];
  assign t[102] = t[167] ^ t[168];
  assign t[103] = t[169] ^ t[170];
  assign t[104] = t[171] ^ t[172];
  assign t[105] = t[173] ^ t[174];
  assign t[106] = t[83] ^ t[86];
  assign t[107] = t[175] ^ t[176];
  assign t[108] = t[117] ^ t[118];
  assign t[109] = t[88] ^ t[119];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[88] & t[119];
  assign t[111] = t[54] & t[59];
  assign t[112] = t[120] ^ t[121];
  assign t[113] = t[122] ^ t[123];
  assign t[114] = t[54] ^ t[124];
  assign t[115] = t[71] ^ t[53];
  assign t[116] = t[125] ^ t[121];
  assign t[117] = t[124] & t[86];
  assign t[118] = t[56] & t[126];
  assign t[119] = t[126] ^ t[87];
  assign t[11] = ~(t[17]);
  assign t[120] = t[127] ^ t[128];
  assign t[121] = t[129] ^ t[111];
  assign t[122] = t[114] & t[115];
  assign t[123] = t[70] & t[53];
  assign t[124] = t[87] ^ t[130];
  assign t[125] = t[131] ^ t[132];
  assign t[126] = t[54] ^ t[67];
  assign t[127] = t[133] ^ t[118];
  assign t[128] = t[72] & t[134];
  assign t[129] = t[38] & t[60];
  assign t[12] = t[139] & t[18];
  assign t[130] = t[50] ^ t[86];
  assign t[131] = t[135] ^ t[123];
  assign t[132] = t[89] & t[71];
  assign t[133] = t[126] ^ t[73];
  assign t[134] = t[86] ^ t[126];
  assign t[135] = t[70] ^ t[53];
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = ~(t[139]);
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = (t[194]);
  assign t[154] = (t[195]);
  assign t[155] = (t[196]);
  assign t[156] = (t[197]);
  assign t[157] = (t[198]);
  assign t[158] = (t[199]);
  assign t[159] = (t[200]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[201]);
  assign t[161] = (t[202]);
  assign t[162] = (t[203]);
  assign t[163] = (t[204]);
  assign t[164] = (t[205]);
  assign t[165] = (t[206]);
  assign t[166] = (t[207]);
  assign t[167] = (t[208]);
  assign t[168] = (t[209]);
  assign t[169] = (t[210]);
  assign t[16] = t[23] ^ t[24];
  assign t[170] = (t[211]);
  assign t[171] = (t[212]);
  assign t[172] = (t[213]);
  assign t[173] = (t[214]);
  assign t[174] = (t[215]);
  assign t[175] = (t[216]);
  assign t[176] = (t[217]);
  assign t[177] = t[218] ^ x[2];
  assign t[178] = t[219] ^ x[6];
  assign t[179] = t[220] ^ x[9];
  assign t[17] = ~(t[139] & t[25]);
  assign t[180] = t[221] ^ x[12];
  assign t[181] = t[222] ^ x[15];
  assign t[182] = t[223] ^ x[18];
  assign t[183] = t[224] ^ x[21];
  assign t[184] = t[225] ^ x[24];
  assign t[185] = t[226] ^ x[27];
  assign t[186] = t[227] ^ x[30];
  assign t[187] = t[228] ^ x[33];
  assign t[188] = t[229] ^ x[36];
  assign t[189] = t[230] ^ x[39];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[231] ^ x[42];
  assign t[191] = t[232] ^ x[45];
  assign t[192] = t[233] ^ x[48];
  assign t[193] = t[234] ^ x[51];
  assign t[194] = t[235] ^ x[54];
  assign t[195] = t[236] ^ x[57];
  assign t[196] = t[237] ^ x[60];
  assign t[197] = t[238] ^ x[63];
  assign t[198] = t[239] ^ x[66];
  assign t[199] = t[240] ^ x[69];
  assign t[19] = ~(t[140]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[241] ^ x[72];
  assign t[201] = t[242] ^ x[75];
  assign t[202] = t[243] ^ x[78];
  assign t[203] = t[244] ^ x[81];
  assign t[204] = t[245] ^ x[84];
  assign t[205] = t[246] ^ x[87];
  assign t[206] = t[247] ^ x[90];
  assign t[207] = t[248] ^ x[93];
  assign t[208] = t[249] ^ x[96];
  assign t[209] = t[250] ^ x[99];
  assign t[20] = ~(t[139]);
  assign t[210] = t[251] ^ x[102];
  assign t[211] = t[252] ^ x[105];
  assign t[212] = t[253] ^ x[108];
  assign t[213] = t[254] ^ x[111];
  assign t[214] = t[255] ^ x[114];
  assign t[215] = t[256] ^ x[117];
  assign t[216] = t[257] ^ x[120];
  assign t[217] = t[258] ^ x[123];
  assign t[218] = (t[259] & ~t[260]);
  assign t[219] = (t[261] & ~t[262]);
  assign t[21] = ~(t[141]);
  assign t[220] = (t[263] & ~t[264]);
  assign t[221] = (t[265] & ~t[266]);
  assign t[222] = (t[267] & ~t[268]);
  assign t[223] = (t[269] & ~t[270]);
  assign t[224] = (t[271] & ~t[272]);
  assign t[225] = (t[273] & ~t[274]);
  assign t[226] = (t[275] & ~t[276]);
  assign t[227] = (t[277] & ~t[278]);
  assign t[228] = (t[279] & ~t[280]);
  assign t[229] = (t[281] & ~t[282]);
  assign t[22] = ~(t[142]);
  assign t[230] = (t[283] & ~t[284]);
  assign t[231] = (t[285] & ~t[286]);
  assign t[232] = (t[287] & ~t[288]);
  assign t[233] = (t[289] & ~t[290]);
  assign t[234] = (t[291] & ~t[292]);
  assign t[235] = (t[293] & ~t[294]);
  assign t[236] = (t[295] & ~t[296]);
  assign t[237] = (t[297] & ~t[298]);
  assign t[238] = (t[299] & ~t[300]);
  assign t[239] = (t[301] & ~t[302]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[303] & ~t[304]);
  assign t[241] = (t[305] & ~t[306]);
  assign t[242] = (t[307] & ~t[308]);
  assign t[243] = (t[309] & ~t[310]);
  assign t[244] = (t[311] & ~t[312]);
  assign t[245] = (t[313] & ~t[314]);
  assign t[246] = (t[315] & ~t[316]);
  assign t[247] = (t[317] & ~t[318]);
  assign t[248] = (t[319] & ~t[320]);
  assign t[249] = (t[321] & ~t[322]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[323] & ~t[324]);
  assign t[251] = (t[325] & ~t[326]);
  assign t[252] = (t[327] & ~t[328]);
  assign t[253] = (t[329] & ~t[330]);
  assign t[254] = (t[331] & ~t[332]);
  assign t[255] = (t[333] & ~t[334]);
  assign t[256] = (t[335] & ~t[336]);
  assign t[257] = (t[337] & ~t[338]);
  assign t[258] = (t[339] & ~t[340]);
  assign t[259] = t[341] ^ x[2];
  assign t[25] = ~(t[143] | t[32]);
  assign t[260] = t[342] ^ x[1];
  assign t[261] = t[343] ^ x[6];
  assign t[262] = t[344] ^ x[5];
  assign t[263] = t[345] ^ x[9];
  assign t[264] = t[346] ^ x[8];
  assign t[265] = t[347] ^ x[12];
  assign t[266] = t[348] ^ x[11];
  assign t[267] = t[349] ^ x[15];
  assign t[268] = t[350] ^ x[14];
  assign t[269] = t[351] ^ x[18];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[352] ^ x[17];
  assign t[271] = t[353] ^ x[21];
  assign t[272] = t[354] ^ x[20];
  assign t[273] = t[355] ^ x[24];
  assign t[274] = t[356] ^ x[23];
  assign t[275] = t[357] ^ x[27];
  assign t[276] = t[358] ^ x[26];
  assign t[277] = t[359] ^ x[30];
  assign t[278] = t[360] ^ x[29];
  assign t[279] = t[361] ^ x[33];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[362] ^ x[32];
  assign t[281] = t[363] ^ x[36];
  assign t[282] = t[364] ^ x[35];
  assign t[283] = t[365] ^ x[39];
  assign t[284] = t[366] ^ x[38];
  assign t[285] = t[367] ^ x[42];
  assign t[286] = t[368] ^ x[41];
  assign t[287] = t[369] ^ x[45];
  assign t[288] = t[370] ^ x[44];
  assign t[289] = t[371] ^ x[48];
  assign t[28] = t[37] & t[38];
  assign t[290] = t[372] ^ x[47];
  assign t[291] = t[373] ^ x[51];
  assign t[292] = t[374] ^ x[50];
  assign t[293] = t[375] ^ x[54];
  assign t[294] = t[376] ^ x[53];
  assign t[295] = t[377] ^ x[57];
  assign t[296] = t[378] ^ x[56];
  assign t[297] = t[379] ^ x[60];
  assign t[298] = t[380] ^ x[59];
  assign t[299] = t[381] ^ x[63];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[62];
  assign t[301] = t[383] ^ x[66];
  assign t[302] = t[384] ^ x[65];
  assign t[303] = t[385] ^ x[69];
  assign t[304] = t[386] ^ x[68];
  assign t[305] = t[387] ^ x[72];
  assign t[306] = t[388] ^ x[71];
  assign t[307] = t[389] ^ x[75];
  assign t[308] = t[390] ^ x[74];
  assign t[309] = t[391] ^ x[78];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[392] ^ x[77];
  assign t[311] = t[393] ^ x[81];
  assign t[312] = t[394] ^ x[80];
  assign t[313] = t[395] ^ x[84];
  assign t[314] = t[396] ^ x[83];
  assign t[315] = t[397] ^ x[87];
  assign t[316] = t[398] ^ x[86];
  assign t[317] = t[399] ^ x[90];
  assign t[318] = t[400] ^ x[89];
  assign t[319] = t[401] ^ x[93];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[402] ^ x[92];
  assign t[321] = t[403] ^ x[96];
  assign t[322] = t[404] ^ x[95];
  assign t[323] = t[405] ^ x[99];
  assign t[324] = t[406] ^ x[98];
  assign t[325] = t[407] ^ x[102];
  assign t[326] = t[408] ^ x[101];
  assign t[327] = t[409] ^ x[105];
  assign t[328] = t[410] ^ x[104];
  assign t[329] = t[411] ^ x[108];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[412] ^ x[107];
  assign t[331] = t[413] ^ x[111];
  assign t[332] = t[414] ^ x[110];
  assign t[333] = t[415] ^ x[114];
  assign t[334] = t[416] ^ x[113];
  assign t[335] = t[417] ^ x[117];
  assign t[336] = t[418] ^ x[116];
  assign t[337] = t[419] ^ x[120];
  assign t[338] = t[420] ^ x[119];
  assign t[339] = t[421] ^ x[123];
  assign t[33] = ~(t[144] & t[145]);
  assign t[340] = t[422] ^ x[122];
  assign t[341] = (x[0]);
  assign t[342] = (x[0]);
  assign t[343] = (x[4]);
  assign t[344] = (x[4]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[146] & t[147]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[148] & t[47]);
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[49]);
  assign t[374] = (x[49]);
  assign t[375] = (x[52]);
  assign t[376] = (x[52]);
  assign t[377] = (x[55]);
  assign t[378] = (x[55]);
  assign t[379] = (x[58]);
  assign t[37] = t[48] ^ t[49];
  assign t[380] = (x[58]);
  assign t[381] = (x[61]);
  assign t[382] = (x[61]);
  assign t[383] = (x[64]);
  assign t[384] = (x[64]);
  assign t[385] = (x[67]);
  assign t[386] = (x[67]);
  assign t[387] = (x[70]);
  assign t[388] = (x[70]);
  assign t[389] = (x[73]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[73]);
  assign t[391] = (x[76]);
  assign t[392] = (x[76]);
  assign t[393] = (x[79]);
  assign t[394] = (x[79]);
  assign t[395] = (x[82]);
  assign t[396] = (x[82]);
  assign t[397] = (x[85]);
  assign t[398] = (x[85]);
  assign t[399] = (x[88]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[88]);
  assign t[401] = (x[91]);
  assign t[402] = (x[91]);
  assign t[403] = (x[94]);
  assign t[404] = (x[94]);
  assign t[405] = (x[97]);
  assign t[406] = (x[97]);
  assign t[407] = (x[100]);
  assign t[408] = (x[100]);
  assign t[409] = (x[103]);
  assign t[40] = t[48] & t[54];
  assign t[410] = (x[103]);
  assign t[411] = (x[106]);
  assign t[412] = (x[106]);
  assign t[413] = (x[109]);
  assign t[414] = (x[109]);
  assign t[415] = (x[112]);
  assign t[416] = (x[112]);
  assign t[417] = (x[115]);
  assign t[418] = (x[115]);
  assign t[419] = (x[118]);
  assign t[41] = t[55] & t[56];
  assign t[420] = (x[118]);
  assign t[421] = (x[121]);
  assign t[422] = (x[121]);
  assign t[42] = t[57] ^ t[58];
  assign t[43] = t[48] & t[59];
  assign t[44] = t[37] & t[60];
  assign t[45] = ~(t[149] | t[150]);
  assign t[46] = ~(t[151] | t[152]);
  assign t[47] = ~(t[153]);
  assign t[48] = t[61] ^ t[62];
  assign t[49] = t[63] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[13] ? t[154] : t[65];
  assign t[51] = t[13] ? t[155] : t[66];
  assign t[52] = t[61] ^ t[63];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[69] ^ t[50];
  assign t[55] = t[62] ^ t[64];
  assign t[56] = t[70] ^ t[38];
  assign t[57] = t[63] & t[71];
  assign t[58] = t[64] & t[72];
  assign t[59] = t[67] ^ t[73];
  assign t[5] = t[9] ? t[137] : x[3];
  assign t[60] = t[54] ^ t[68];
  assign t[61] = t[74] ^ t[75];
  assign t[62] = t[76] ^ t[77];
  assign t[63] = t[78] ^ t[79];
  assign t[64] = t[80] ^ t[81];
  assign t[65] = t[156] ^ t[157];
  assign t[66] = t[158] ^ t[159];
  assign t[67] = t[82] ^ t[83];
  assign t[68] = t[84] ^ t[51];
  assign t[69] = t[13] ? t[160] : t[85];
  assign t[6] = ~(t[10] ^ t[138]);
  assign t[70] = t[69] ^ t[83];
  assign t[71] = t[86] ^ t[87];
  assign t[72] = t[88] ^ t[89];
  assign t[73] = t[90] ^ t[51];
  assign t[74] = t[91] ^ t[92];
  assign t[75] = t[93] & t[94];
  assign t[76] = t[95] ^ t[96];
  assign t[77] = t[97] & t[98];
  assign t[78] = t[94] & t[99];
  assign t[79] = t[94] ^ t[100];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[98] & t[101];
  assign t[81] = t[98] ^ t[100];
  assign t[82] = t[13] ? t[161] : t[102];
  assign t[83] = t[13] ? t[162] : t[103];
  assign t[84] = t[13] ? t[163] : t[104];
  assign t[85] = t[164] ^ t[138];
  assign t[86] = t[13] ? t[165] : t[105];
  assign t[87] = t[90] ^ t[84];
  assign t[88] = t[69] ^ t[51];
  assign t[89] = t[87] ^ t[106];
  assign t[8] = ~(t[13]);
  assign t[90] = t[13] ? t[166] : t[107];
  assign t[91] = t[108] ^ t[109];
  assign t[92] = t[110] ^ t[111];
  assign t[93] = t[76] ^ t[100];
  assign t[94] = t[112] ^ t[74];
  assign t[95] = t[113] ^ t[92];
  assign t[96] = t[114] ^ t[115];
  assign t[97] = t[74] ^ t[100];
  assign t[98] = t[116] ^ t[76];
  assign t[99] = t[112] & t[76];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [123:0] x;
 output y;

 wire [422:0] t;
  assign t[0] = t[1] ? t[2] : t[136];
  assign t[100] = t[116] & t[112];
  assign t[101] = t[74] & t[116];
  assign t[102] = t[167] ^ t[168];
  assign t[103] = t[169] ^ t[170];
  assign t[104] = t[171] ^ t[172];
  assign t[105] = t[173] ^ t[174];
  assign t[106] = t[83] ^ t[86];
  assign t[107] = t[175] ^ t[176];
  assign t[108] = t[117] ^ t[118];
  assign t[109] = t[88] ^ t[119];
  assign t[10] = ~(t[15] ^ t[16]);
  assign t[110] = t[88] & t[119];
  assign t[111] = t[54] & t[59];
  assign t[112] = t[120] ^ t[121];
  assign t[113] = t[122] ^ t[123];
  assign t[114] = t[54] ^ t[124];
  assign t[115] = t[71] ^ t[53];
  assign t[116] = t[125] ^ t[121];
  assign t[117] = t[124] & t[86];
  assign t[118] = t[56] & t[126];
  assign t[119] = t[126] ^ t[87];
  assign t[11] = ~(t[17]);
  assign t[120] = t[127] ^ t[128];
  assign t[121] = t[129] ^ t[111];
  assign t[122] = t[114] & t[115];
  assign t[123] = t[70] & t[53];
  assign t[124] = t[87] ^ t[130];
  assign t[125] = t[131] ^ t[132];
  assign t[126] = t[54] ^ t[67];
  assign t[127] = t[133] ^ t[118];
  assign t[128] = t[72] & t[134];
  assign t[129] = t[38] & t[60];
  assign t[12] = t[139] & t[18];
  assign t[130] = t[50] ^ t[86];
  assign t[131] = t[135] ^ t[123];
  assign t[132] = t[89] & t[71];
  assign t[133] = t[126] ^ t[73];
  assign t[134] = t[86] ^ t[126];
  assign t[135] = t[70] ^ t[53];
  assign t[136] = (t[177]);
  assign t[137] = (t[178]);
  assign t[138] = (t[179]);
  assign t[139] = (t[180]);
  assign t[13] = ~(t[19] | t[20]);
  assign t[140] = (t[181]);
  assign t[141] = (t[182]);
  assign t[142] = (t[183]);
  assign t[143] = (t[184]);
  assign t[144] = (t[185]);
  assign t[145] = (t[186]);
  assign t[146] = (t[187]);
  assign t[147] = (t[188]);
  assign t[148] = (t[189]);
  assign t[149] = (t[190]);
  assign t[14] = ~(t[139]);
  assign t[150] = (t[191]);
  assign t[151] = (t[192]);
  assign t[152] = (t[193]);
  assign t[153] = (t[194]);
  assign t[154] = (t[195]);
  assign t[155] = (t[196]);
  assign t[156] = (t[197]);
  assign t[157] = (t[198]);
  assign t[158] = (t[199]);
  assign t[159] = (t[200]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[160] = (t[201]);
  assign t[161] = (t[202]);
  assign t[162] = (t[203]);
  assign t[163] = (t[204]);
  assign t[164] = (t[205]);
  assign t[165] = (t[206]);
  assign t[166] = (t[207]);
  assign t[167] = (t[208]);
  assign t[168] = (t[209]);
  assign t[169] = (t[210]);
  assign t[16] = t[23] ^ t[24];
  assign t[170] = (t[211]);
  assign t[171] = (t[212]);
  assign t[172] = (t[213]);
  assign t[173] = (t[214]);
  assign t[174] = (t[215]);
  assign t[175] = (t[216]);
  assign t[176] = (t[217]);
  assign t[177] = t[218] ^ x[2];
  assign t[178] = t[219] ^ x[6];
  assign t[179] = t[220] ^ x[9];
  assign t[17] = ~(t[139] & t[25]);
  assign t[180] = t[221] ^ x[12];
  assign t[181] = t[222] ^ x[15];
  assign t[182] = t[223] ^ x[18];
  assign t[183] = t[224] ^ x[21];
  assign t[184] = t[225] ^ x[24];
  assign t[185] = t[226] ^ x[27];
  assign t[186] = t[227] ^ x[30];
  assign t[187] = t[228] ^ x[33];
  assign t[188] = t[229] ^ x[36];
  assign t[189] = t[230] ^ x[39];
  assign t[18] = t[26] & t[27];
  assign t[190] = t[231] ^ x[42];
  assign t[191] = t[232] ^ x[45];
  assign t[192] = t[233] ^ x[48];
  assign t[193] = t[234] ^ x[51];
  assign t[194] = t[235] ^ x[54];
  assign t[195] = t[236] ^ x[57];
  assign t[196] = t[237] ^ x[60];
  assign t[197] = t[238] ^ x[63];
  assign t[198] = t[239] ^ x[66];
  assign t[199] = t[240] ^ x[69];
  assign t[19] = ~(t[140]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[241] ^ x[72];
  assign t[201] = t[242] ^ x[75];
  assign t[202] = t[243] ^ x[78];
  assign t[203] = t[244] ^ x[81];
  assign t[204] = t[245] ^ x[84];
  assign t[205] = t[246] ^ x[87];
  assign t[206] = t[247] ^ x[90];
  assign t[207] = t[248] ^ x[93];
  assign t[208] = t[249] ^ x[96];
  assign t[209] = t[250] ^ x[99];
  assign t[20] = ~(t[139]);
  assign t[210] = t[251] ^ x[102];
  assign t[211] = t[252] ^ x[105];
  assign t[212] = t[253] ^ x[108];
  assign t[213] = t[254] ^ x[111];
  assign t[214] = t[255] ^ x[114];
  assign t[215] = t[256] ^ x[117];
  assign t[216] = t[257] ^ x[120];
  assign t[217] = t[258] ^ x[123];
  assign t[218] = (t[259] & ~t[260]);
  assign t[219] = (t[261] & ~t[262]);
  assign t[21] = ~(t[141]);
  assign t[220] = (t[263] & ~t[264]);
  assign t[221] = (t[265] & ~t[266]);
  assign t[222] = (t[267] & ~t[268]);
  assign t[223] = (t[269] & ~t[270]);
  assign t[224] = (t[271] & ~t[272]);
  assign t[225] = (t[273] & ~t[274]);
  assign t[226] = (t[275] & ~t[276]);
  assign t[227] = (t[277] & ~t[278]);
  assign t[228] = (t[279] & ~t[280]);
  assign t[229] = (t[281] & ~t[282]);
  assign t[22] = ~(t[142]);
  assign t[230] = (t[283] & ~t[284]);
  assign t[231] = (t[285] & ~t[286]);
  assign t[232] = (t[287] & ~t[288]);
  assign t[233] = (t[289] & ~t[290]);
  assign t[234] = (t[291] & ~t[292]);
  assign t[235] = (t[293] & ~t[294]);
  assign t[236] = (t[295] & ~t[296]);
  assign t[237] = (t[297] & ~t[298]);
  assign t[238] = (t[299] & ~t[300]);
  assign t[239] = (t[301] & ~t[302]);
  assign t[23] = t[28] ^ t[29];
  assign t[240] = (t[303] & ~t[304]);
  assign t[241] = (t[305] & ~t[306]);
  assign t[242] = (t[307] & ~t[308]);
  assign t[243] = (t[309] & ~t[310]);
  assign t[244] = (t[311] & ~t[312]);
  assign t[245] = (t[313] & ~t[314]);
  assign t[246] = (t[315] & ~t[316]);
  assign t[247] = (t[317] & ~t[318]);
  assign t[248] = (t[319] & ~t[320]);
  assign t[249] = (t[321] & ~t[322]);
  assign t[24] = t[30] ^ t[31];
  assign t[250] = (t[323] & ~t[324]);
  assign t[251] = (t[325] & ~t[326]);
  assign t[252] = (t[327] & ~t[328]);
  assign t[253] = (t[329] & ~t[330]);
  assign t[254] = (t[331] & ~t[332]);
  assign t[255] = (t[333] & ~t[334]);
  assign t[256] = (t[335] & ~t[336]);
  assign t[257] = (t[337] & ~t[338]);
  assign t[258] = (t[339] & ~t[340]);
  assign t[259] = t[341] ^ x[2];
  assign t[25] = ~(t[143] | t[32]);
  assign t[260] = t[342] ^ x[1];
  assign t[261] = t[343] ^ x[6];
  assign t[262] = t[344] ^ x[5];
  assign t[263] = t[345] ^ x[9];
  assign t[264] = t[346] ^ x[8];
  assign t[265] = t[347] ^ x[12];
  assign t[266] = t[348] ^ x[11];
  assign t[267] = t[349] ^ x[15];
  assign t[268] = t[350] ^ x[14];
  assign t[269] = t[351] ^ x[18];
  assign t[26] = ~(t[33] | t[34]);
  assign t[270] = t[352] ^ x[17];
  assign t[271] = t[353] ^ x[21];
  assign t[272] = t[354] ^ x[20];
  assign t[273] = t[355] ^ x[24];
  assign t[274] = t[356] ^ x[23];
  assign t[275] = t[357] ^ x[27];
  assign t[276] = t[358] ^ x[26];
  assign t[277] = t[359] ^ x[30];
  assign t[278] = t[360] ^ x[29];
  assign t[279] = t[361] ^ x[33];
  assign t[27] = ~(t[35] | t[36]);
  assign t[280] = t[362] ^ x[32];
  assign t[281] = t[363] ^ x[36];
  assign t[282] = t[364] ^ x[35];
  assign t[283] = t[365] ^ x[39];
  assign t[284] = t[366] ^ x[38];
  assign t[285] = t[367] ^ x[42];
  assign t[286] = t[368] ^ x[41];
  assign t[287] = t[369] ^ x[45];
  assign t[288] = t[370] ^ x[44];
  assign t[289] = t[371] ^ x[48];
  assign t[28] = t[37] & t[38];
  assign t[290] = t[372] ^ x[47];
  assign t[291] = t[373] ^ x[51];
  assign t[292] = t[374] ^ x[50];
  assign t[293] = t[375] ^ x[54];
  assign t[294] = t[376] ^ x[53];
  assign t[295] = t[377] ^ x[57];
  assign t[296] = t[378] ^ x[56];
  assign t[297] = t[379] ^ x[60];
  assign t[298] = t[380] ^ x[59];
  assign t[299] = t[381] ^ x[63];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[6] : t[5];
  assign t[300] = t[382] ^ x[62];
  assign t[301] = t[383] ^ x[66];
  assign t[302] = t[384] ^ x[65];
  assign t[303] = t[385] ^ x[69];
  assign t[304] = t[386] ^ x[68];
  assign t[305] = t[387] ^ x[72];
  assign t[306] = t[388] ^ x[71];
  assign t[307] = t[389] ^ x[75];
  assign t[308] = t[390] ^ x[74];
  assign t[309] = t[391] ^ x[78];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[392] ^ x[77];
  assign t[311] = t[393] ^ x[81];
  assign t[312] = t[394] ^ x[80];
  assign t[313] = t[395] ^ x[84];
  assign t[314] = t[396] ^ x[83];
  assign t[315] = t[397] ^ x[87];
  assign t[316] = t[398] ^ x[86];
  assign t[317] = t[399] ^ x[90];
  assign t[318] = t[400] ^ x[89];
  assign t[319] = t[401] ^ x[93];
  assign t[31] = t[43] ^ t[44];
  assign t[320] = t[402] ^ x[92];
  assign t[321] = t[403] ^ x[96];
  assign t[322] = t[404] ^ x[95];
  assign t[323] = t[405] ^ x[99];
  assign t[324] = t[406] ^ x[98];
  assign t[325] = t[407] ^ x[102];
  assign t[326] = t[408] ^ x[101];
  assign t[327] = t[409] ^ x[105];
  assign t[328] = t[410] ^ x[104];
  assign t[329] = t[411] ^ x[108];
  assign t[32] = ~(t[45] & t[46]);
  assign t[330] = t[412] ^ x[107];
  assign t[331] = t[413] ^ x[111];
  assign t[332] = t[414] ^ x[110];
  assign t[333] = t[415] ^ x[114];
  assign t[334] = t[416] ^ x[113];
  assign t[335] = t[417] ^ x[117];
  assign t[336] = t[418] ^ x[116];
  assign t[337] = t[419] ^ x[120];
  assign t[338] = t[420] ^ x[119];
  assign t[339] = t[421] ^ x[123];
  assign t[33] = ~(t[144] & t[145]);
  assign t[340] = t[422] ^ x[122];
  assign t[341] = (x[0]);
  assign t[342] = (x[0]);
  assign t[343] = (x[4]);
  assign t[344] = (x[4]);
  assign t[345] = (x[7]);
  assign t[346] = (x[7]);
  assign t[347] = (x[10]);
  assign t[348] = (x[10]);
  assign t[349] = (x[13]);
  assign t[34] = ~(t[146] & t[147]);
  assign t[350] = (x[13]);
  assign t[351] = (x[16]);
  assign t[352] = (x[16]);
  assign t[353] = (x[19]);
  assign t[354] = (x[19]);
  assign t[355] = (x[22]);
  assign t[356] = (x[22]);
  assign t[357] = (x[25]);
  assign t[358] = (x[25]);
  assign t[359] = (x[28]);
  assign t[35] = ~(t[25]);
  assign t[360] = (x[28]);
  assign t[361] = (x[31]);
  assign t[362] = (x[31]);
  assign t[363] = (x[34]);
  assign t[364] = (x[34]);
  assign t[365] = (x[37]);
  assign t[366] = (x[37]);
  assign t[367] = (x[40]);
  assign t[368] = (x[40]);
  assign t[369] = (x[43]);
  assign t[36] = ~(t[148] & t[47]);
  assign t[370] = (x[43]);
  assign t[371] = (x[46]);
  assign t[372] = (x[46]);
  assign t[373] = (x[49]);
  assign t[374] = (x[49]);
  assign t[375] = (x[52]);
  assign t[376] = (x[52]);
  assign t[377] = (x[55]);
  assign t[378] = (x[55]);
  assign t[379] = (x[58]);
  assign t[37] = t[48] ^ t[49];
  assign t[380] = (x[58]);
  assign t[381] = (x[61]);
  assign t[382] = (x[61]);
  assign t[383] = (x[64]);
  assign t[384] = (x[64]);
  assign t[385] = (x[67]);
  assign t[386] = (x[67]);
  assign t[387] = (x[70]);
  assign t[388] = (x[70]);
  assign t[389] = (x[73]);
  assign t[38] = t[50] ^ t[51];
  assign t[390] = (x[73]);
  assign t[391] = (x[76]);
  assign t[392] = (x[76]);
  assign t[393] = (x[79]);
  assign t[394] = (x[79]);
  assign t[395] = (x[82]);
  assign t[396] = (x[82]);
  assign t[397] = (x[85]);
  assign t[398] = (x[85]);
  assign t[399] = (x[88]);
  assign t[39] = t[52] & t[53];
  assign t[3] = ~(t[7]);
  assign t[400] = (x[88]);
  assign t[401] = (x[91]);
  assign t[402] = (x[91]);
  assign t[403] = (x[94]);
  assign t[404] = (x[94]);
  assign t[405] = (x[97]);
  assign t[406] = (x[97]);
  assign t[407] = (x[100]);
  assign t[408] = (x[100]);
  assign t[409] = (x[103]);
  assign t[40] = t[48] & t[54];
  assign t[410] = (x[103]);
  assign t[411] = (x[106]);
  assign t[412] = (x[106]);
  assign t[413] = (x[109]);
  assign t[414] = (x[109]);
  assign t[415] = (x[112]);
  assign t[416] = (x[112]);
  assign t[417] = (x[115]);
  assign t[418] = (x[115]);
  assign t[419] = (x[118]);
  assign t[41] = t[55] & t[56];
  assign t[420] = (x[118]);
  assign t[421] = (x[121]);
  assign t[422] = (x[121]);
  assign t[42] = t[57] ^ t[58];
  assign t[43] = t[48] & t[59];
  assign t[44] = t[37] & t[60];
  assign t[45] = ~(t[149] | t[150]);
  assign t[46] = ~(t[151] | t[152]);
  assign t[47] = ~(t[153]);
  assign t[48] = t[61] ^ t[62];
  assign t[49] = t[63] ^ t[64];
  assign t[4] = ~(t[8]);
  assign t[50] = t[13] ? t[154] : t[65];
  assign t[51] = t[13] ? t[155] : t[66];
  assign t[52] = t[61] ^ t[63];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[69] ^ t[50];
  assign t[55] = t[62] ^ t[64];
  assign t[56] = t[70] ^ t[38];
  assign t[57] = t[63] & t[71];
  assign t[58] = t[64] & t[72];
  assign t[59] = t[67] ^ t[73];
  assign t[5] = t[9] ? t[137] : x[3];
  assign t[60] = t[54] ^ t[68];
  assign t[61] = t[74] ^ t[75];
  assign t[62] = t[76] ^ t[77];
  assign t[63] = t[78] ^ t[79];
  assign t[64] = t[80] ^ t[81];
  assign t[65] = t[156] ^ t[157];
  assign t[66] = t[158] ^ t[159];
  assign t[67] = t[82] ^ t[83];
  assign t[68] = t[84] ^ t[51];
  assign t[69] = t[13] ? t[160] : t[85];
  assign t[6] = ~(t[10] ^ t[138]);
  assign t[70] = t[69] ^ t[83];
  assign t[71] = t[86] ^ t[87];
  assign t[72] = t[88] ^ t[89];
  assign t[73] = t[90] ^ t[51];
  assign t[74] = t[91] ^ t[92];
  assign t[75] = t[93] & t[94];
  assign t[76] = t[95] ^ t[96];
  assign t[77] = t[97] & t[98];
  assign t[78] = t[94] & t[99];
  assign t[79] = t[94] ^ t[100];
  assign t[7] = ~(t[11] | t[12]);
  assign t[80] = t[98] & t[101];
  assign t[81] = t[98] ^ t[100];
  assign t[82] = t[13] ? t[161] : t[102];
  assign t[83] = t[13] ? t[162] : t[103];
  assign t[84] = t[13] ? t[163] : t[104];
  assign t[85] = t[164] ^ t[138];
  assign t[86] = t[13] ? t[165] : t[105];
  assign t[87] = t[90] ^ t[84];
  assign t[88] = t[69] ^ t[51];
  assign t[89] = t[87] ^ t[106];
  assign t[8] = ~(t[13]);
  assign t[90] = t[13] ? t[166] : t[107];
  assign t[91] = t[108] ^ t[109];
  assign t[92] = t[110] ^ t[111];
  assign t[93] = t[76] ^ t[100];
  assign t[94] = t[112] ^ t[74];
  assign t[95] = t[113] ^ t[92];
  assign t[96] = t[114] ^ t[115];
  assign t[97] = t[74] ^ t[100];
  assign t[98] = t[116] ^ t[76];
  assign t[99] = t[112] & t[76];
  assign t[9] = ~(t[14]);
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind251(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind255(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind256(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind257(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind258(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind259(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind260(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind261(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind262(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind263(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind264(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind265(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind266(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind267(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind268(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind269(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind270(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind271(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind272(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind273(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind274(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind275(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind276(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind277(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind278(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind279(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind280(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind281(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind282(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind283(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind284(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind285(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind286(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind287(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind288(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind289(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind290(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind291(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind292(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind293(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind294(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind295(x, y);
 input [48:0] x;
 output y;

 wire [139:0] t;
  assign t[0] = t[1] ? t[2] : t[28];
  assign t[100] = t[132] ^ x[39];
  assign t[101] = t[133] ^ x[38];
  assign t[102] = t[134] ^ x[42];
  assign t[103] = t[135] ^ x[41];
  assign t[104] = t[136] ^ x[45];
  assign t[105] = t[137] ^ x[44];
  assign t[106] = t[138] ^ x[48];
  assign t[107] = t[139] ^ x[47];
  assign t[108] = (x[0]);
  assign t[109] = (x[0]);
  assign t[10] = t[31] & t[14];
  assign t[110] = (x[3]);
  assign t[111] = (x[3]);
  assign t[112] = (x[7]);
  assign t[113] = (x[7]);
  assign t[114] = (x[10]);
  assign t[115] = (x[10]);
  assign t[116] = (x[13]);
  assign t[117] = (x[13]);
  assign t[118] = (x[16]);
  assign t[119] = (x[16]);
  assign t[11] = ~(t[15] | t[16]);
  assign t[120] = (x[19]);
  assign t[121] = (x[19]);
  assign t[122] = (x[22]);
  assign t[123] = (x[22]);
  assign t[124] = (x[25]);
  assign t[125] = (x[25]);
  assign t[126] = (x[28]);
  assign t[127] = (x[28]);
  assign t[128] = (x[31]);
  assign t[129] = (x[31]);
  assign t[12] = ~(t[31]);
  assign t[130] = (x[34]);
  assign t[131] = (x[34]);
  assign t[132] = (x[37]);
  assign t[133] = (x[37]);
  assign t[134] = (x[40]);
  assign t[135] = (x[40]);
  assign t[136] = (x[43]);
  assign t[137] = (x[43]);
  assign t[138] = (x[46]);
  assign t[139] = (x[46]);
  assign t[13] = ~(t[31] & t[17]);
  assign t[14] = t[18] & t[19];
  assign t[15] = ~(t[32]);
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[33] | t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[25] & t[26]);
  assign t[21] = ~(t[34] & t[35]);
  assign t[22] = ~(t[36] & t[37]);
  assign t[23] = ~(t[17]);
  assign t[24] = ~(t[38] & t[27]);
  assign t[25] = ~(t[39] | t[40]);
  assign t[26] = ~(t[41] | t[42]);
  assign t[27] = ~(t[43]);
  assign t[28] = (t[44]);
  assign t[29] = (t[45]);
  assign t[2] = t[4] ? t[29] : t[5];
  assign t[30] = (t[46]);
  assign t[31] = (t[47]);
  assign t[32] = (t[48]);
  assign t[33] = (t[49]);
  assign t[34] = (t[50]);
  assign t[35] = (t[51]);
  assign t[36] = (t[52]);
  assign t[37] = (t[53]);
  assign t[38] = (t[54]);
  assign t[39] = (t[55]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[56]);
  assign t[41] = (t[57]);
  assign t[42] = (t[58]);
  assign t[43] = (t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[5];
  assign t[46] = t[62] ^ x[9];
  assign t[47] = t[63] ^ x[12];
  assign t[48] = t[64] ^ x[15];
  assign t[49] = t[65] ^ x[18];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[24];
  assign t[52] = t[68] ^ x[27];
  assign t[53] = t[69] ^ x[30];
  assign t[54] = t[70] ^ x[33];
  assign t[55] = t[71] ^ x[36];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[42];
  assign t[58] = t[74] ^ x[45];
  assign t[59] = t[75] ^ x[48];
  assign t[5] = t[8] ? t[30] : x[6];
  assign t[60] = (t[76] & ~t[77]);
  assign t[61] = (t[78] & ~t[79]);
  assign t[62] = (t[80] & ~t[81]);
  assign t[63] = (t[82] & ~t[83]);
  assign t[64] = (t[84] & ~t[85]);
  assign t[65] = (t[86] & ~t[87]);
  assign t[66] = (t[88] & ~t[89]);
  assign t[67] = (t[90] & ~t[91]);
  assign t[68] = (t[92] & ~t[93]);
  assign t[69] = (t[94] & ~t[95]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = (t[96] & ~t[97]);
  assign t[71] = (t[98] & ~t[99]);
  assign t[72] = (t[100] & ~t[101]);
  assign t[73] = (t[102] & ~t[103]);
  assign t[74] = (t[104] & ~t[105]);
  assign t[75] = (t[106] & ~t[107]);
  assign t[76] = t[108] ^ x[2];
  assign t[77] = t[109] ^ x[1];
  assign t[78] = t[110] ^ x[5];
  assign t[79] = t[111] ^ x[4];
  assign t[7] = ~(t[11]);
  assign t[80] = t[112] ^ x[9];
  assign t[81] = t[113] ^ x[8];
  assign t[82] = t[114] ^ x[12];
  assign t[83] = t[115] ^ x[11];
  assign t[84] = t[116] ^ x[15];
  assign t[85] = t[117] ^ x[14];
  assign t[86] = t[118] ^ x[18];
  assign t[87] = t[119] ^ x[17];
  assign t[88] = t[120] ^ x[21];
  assign t[89] = t[121] ^ x[20];
  assign t[8] = ~(t[12]);
  assign t[90] = t[122] ^ x[24];
  assign t[91] = t[123] ^ x[23];
  assign t[92] = t[124] ^ x[27];
  assign t[93] = t[125] ^ x[26];
  assign t[94] = t[126] ^ x[30];
  assign t[95] = t[127] ^ x[29];
  assign t[96] = t[128] ^ x[33];
  assign t[97] = t[129] ^ x[32];
  assign t[98] = t[130] ^ x[36];
  assign t[99] = t[131] ^ x[35];
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind296(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind297(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind298(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind299(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind300(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind301(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind302(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind303(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind304(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind305(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind306(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind307(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind308(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind309(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind310(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind311(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind312(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind313(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind314(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind315(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind316(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind317(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind318(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind319(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind320(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind321(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind322(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind323(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind324(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind325(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind326(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind327(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind328(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind329(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind330(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind331(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind332(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind333(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind334(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind335(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind336(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind337(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind338(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind339(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind340(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind341(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind342(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind343(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[25] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[6];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[3];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[6];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[5];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[4]);
  assign t[98] = (x[4]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind344(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind345(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind346(x, y);
 input [66:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = (t[142] & ~t[143]);
  assign t[103] = (t[144] & ~t[145]);
  assign t[104] = (t[146] & ~t[147]);
  assign t[105] = (t[148] & ~t[149]);
  assign t[106] = t[150] ^ x[2];
  assign t[107] = t[151] ^ x[1];
  assign t[108] = t[152] ^ x[6];
  assign t[109] = t[153] ^ x[5];
  assign t[10] = t[42] & t[15];
  assign t[110] = t[154] ^ x[9];
  assign t[111] = t[155] ^ x[8];
  assign t[112] = t[156] ^ x[12];
  assign t[113] = t[157] ^ x[11];
  assign t[114] = t[158] ^ x[15];
  assign t[115] = t[159] ^ x[14];
  assign t[116] = t[160] ^ x[18];
  assign t[117] = t[161] ^ x[17];
  assign t[118] = t[162] ^ x[21];
  assign t[119] = t[163] ^ x[20];
  assign t[11] = ~(t[16]);
  assign t[120] = t[164] ^ x[24];
  assign t[121] = t[165] ^ x[23];
  assign t[122] = t[166] ^ x[27];
  assign t[123] = t[167] ^ x[26];
  assign t[124] = t[168] ^ x[30];
  assign t[125] = t[169] ^ x[29];
  assign t[126] = t[170] ^ x[33];
  assign t[127] = t[171] ^ x[32];
  assign t[128] = t[172] ^ x[36];
  assign t[129] = t[173] ^ x[35];
  assign t[12] = ~(t[42]);
  assign t[130] = t[174] ^ x[39];
  assign t[131] = t[175] ^ x[38];
  assign t[132] = t[176] ^ x[42];
  assign t[133] = t[177] ^ x[41];
  assign t[134] = t[178] ^ x[45];
  assign t[135] = t[179] ^ x[44];
  assign t[136] = t[180] ^ x[48];
  assign t[137] = t[181] ^ x[47];
  assign t[138] = t[182] ^ x[51];
  assign t[139] = t[183] ^ x[50];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[54];
  assign t[141] = t[185] ^ x[53];
  assign t[142] = t[186] ^ x[57];
  assign t[143] = t[187] ^ x[56];
  assign t[144] = t[188] ^ x[60];
  assign t[145] = t[189] ^ x[59];
  assign t[146] = t[190] ^ x[63];
  assign t[147] = t[191] ^ x[62];
  assign t[148] = t[192] ^ x[66];
  assign t[149] = t[193] ^ x[65];
  assign t[14] = t[18] ? t[43] : t[19];
  assign t[150] = (x[0]);
  assign t[151] = (x[0]);
  assign t[152] = (x[4]);
  assign t[153] = (x[4]);
  assign t[154] = (x[7]);
  assign t[155] = (x[7]);
  assign t[156] = (x[10]);
  assign t[157] = (x[10]);
  assign t[158] = (x[13]);
  assign t[159] = (x[13]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[16]);
  assign t[161] = (x[16]);
  assign t[162] = (x[19]);
  assign t[163] = (x[19]);
  assign t[164] = (x[22]);
  assign t[165] = (x[22]);
  assign t[166] = (x[25]);
  assign t[167] = (x[25]);
  assign t[168] = (x[28]);
  assign t[169] = (x[28]);
  assign t[16] = ~(t[42] & t[22]);
  assign t[170] = (x[31]);
  assign t[171] = (x[31]);
  assign t[172] = (x[34]);
  assign t[173] = (x[34]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[40]);
  assign t[177] = (x[40]);
  assign t[178] = (x[43]);
  assign t[179] = (x[43]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[46]);
  assign t[181] = (x[46]);
  assign t[182] = (x[49]);
  assign t[183] = (x[49]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[55]);
  assign t[187] = (x[55]);
  assign t[188] = (x[58]);
  assign t[189] = (x[58]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[61]);
  assign t[191] = (x[61]);
  assign t[192] = (x[64]);
  assign t[193] = (x[64]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[44] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[40] : t[5];
  assign t[30] = ~(t[51] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[42]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[41] ^ t[39];
  assign t[36] = ~(t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = (t[82]);
  assign t[61] = (t[83]);
  assign t[62] = t[84] ^ x[2];
  assign t[63] = t[85] ^ x[6];
  assign t[64] = t[86] ^ x[9];
  assign t[65] = t[87] ^ x[12];
  assign t[66] = t[88] ^ x[15];
  assign t[67] = t[89] ^ x[18];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[24];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[27];
  assign t[71] = t[93] ^ x[30];
  assign t[72] = t[94] ^ x[33];
  assign t[73] = t[95] ^ x[36];
  assign t[74] = t[96] ^ x[39];
  assign t[75] = t[97] ^ x[42];
  assign t[76] = t[98] ^ x[45];
  assign t[77] = t[99] ^ x[48];
  assign t[78] = t[100] ^ x[51];
  assign t[79] = t[101] ^ x[54];
  assign t[7] = ~(t[11]);
  assign t[80] = t[102] ^ x[57];
  assign t[81] = t[103] ^ x[60];
  assign t[82] = t[104] ^ x[63];
  assign t[83] = t[105] ^ x[66];
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind347(x, y);
 input [66:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = (t[142] & ~t[143]);
  assign t[103] = (t[144] & ~t[145]);
  assign t[104] = (t[146] & ~t[147]);
  assign t[105] = (t[148] & ~t[149]);
  assign t[106] = t[150] ^ x[2];
  assign t[107] = t[151] ^ x[1];
  assign t[108] = t[152] ^ x[6];
  assign t[109] = t[153] ^ x[5];
  assign t[10] = t[42] & t[15];
  assign t[110] = t[154] ^ x[9];
  assign t[111] = t[155] ^ x[8];
  assign t[112] = t[156] ^ x[12];
  assign t[113] = t[157] ^ x[11];
  assign t[114] = t[158] ^ x[15];
  assign t[115] = t[159] ^ x[14];
  assign t[116] = t[160] ^ x[18];
  assign t[117] = t[161] ^ x[17];
  assign t[118] = t[162] ^ x[21];
  assign t[119] = t[163] ^ x[20];
  assign t[11] = ~(t[16]);
  assign t[120] = t[164] ^ x[24];
  assign t[121] = t[165] ^ x[23];
  assign t[122] = t[166] ^ x[27];
  assign t[123] = t[167] ^ x[26];
  assign t[124] = t[168] ^ x[30];
  assign t[125] = t[169] ^ x[29];
  assign t[126] = t[170] ^ x[33];
  assign t[127] = t[171] ^ x[32];
  assign t[128] = t[172] ^ x[36];
  assign t[129] = t[173] ^ x[35];
  assign t[12] = ~(t[42]);
  assign t[130] = t[174] ^ x[39];
  assign t[131] = t[175] ^ x[38];
  assign t[132] = t[176] ^ x[42];
  assign t[133] = t[177] ^ x[41];
  assign t[134] = t[178] ^ x[45];
  assign t[135] = t[179] ^ x[44];
  assign t[136] = t[180] ^ x[48];
  assign t[137] = t[181] ^ x[47];
  assign t[138] = t[182] ^ x[51];
  assign t[139] = t[183] ^ x[50];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[54];
  assign t[141] = t[185] ^ x[53];
  assign t[142] = t[186] ^ x[57];
  assign t[143] = t[187] ^ x[56];
  assign t[144] = t[188] ^ x[60];
  assign t[145] = t[189] ^ x[59];
  assign t[146] = t[190] ^ x[63];
  assign t[147] = t[191] ^ x[62];
  assign t[148] = t[192] ^ x[66];
  assign t[149] = t[193] ^ x[65];
  assign t[14] = t[18] ? t[43] : t[19];
  assign t[150] = (x[0]);
  assign t[151] = (x[0]);
  assign t[152] = (x[4]);
  assign t[153] = (x[4]);
  assign t[154] = (x[7]);
  assign t[155] = (x[7]);
  assign t[156] = (x[10]);
  assign t[157] = (x[10]);
  assign t[158] = (x[13]);
  assign t[159] = (x[13]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[16]);
  assign t[161] = (x[16]);
  assign t[162] = (x[19]);
  assign t[163] = (x[19]);
  assign t[164] = (x[22]);
  assign t[165] = (x[22]);
  assign t[166] = (x[25]);
  assign t[167] = (x[25]);
  assign t[168] = (x[28]);
  assign t[169] = (x[28]);
  assign t[16] = ~(t[42] & t[22]);
  assign t[170] = (x[31]);
  assign t[171] = (x[31]);
  assign t[172] = (x[34]);
  assign t[173] = (x[34]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[40]);
  assign t[177] = (x[40]);
  assign t[178] = (x[43]);
  assign t[179] = (x[43]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[46]);
  assign t[181] = (x[46]);
  assign t[182] = (x[49]);
  assign t[183] = (x[49]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[55]);
  assign t[187] = (x[55]);
  assign t[188] = (x[58]);
  assign t[189] = (x[58]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[61]);
  assign t[191] = (x[61]);
  assign t[192] = (x[64]);
  assign t[193] = (x[64]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[44] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[40] : t[5];
  assign t[30] = ~(t[51] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[42]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[41] ^ t[39];
  assign t[36] = ~(t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = (t[82]);
  assign t[61] = (t[83]);
  assign t[62] = t[84] ^ x[2];
  assign t[63] = t[85] ^ x[6];
  assign t[64] = t[86] ^ x[9];
  assign t[65] = t[87] ^ x[12];
  assign t[66] = t[88] ^ x[15];
  assign t[67] = t[89] ^ x[18];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[24];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[27];
  assign t[71] = t[93] ^ x[30];
  assign t[72] = t[94] ^ x[33];
  assign t[73] = t[95] ^ x[36];
  assign t[74] = t[96] ^ x[39];
  assign t[75] = t[97] ^ x[42];
  assign t[76] = t[98] ^ x[45];
  assign t[77] = t[99] ^ x[48];
  assign t[78] = t[100] ^ x[51];
  assign t[79] = t[101] ^ x[54];
  assign t[7] = ~(t[11]);
  assign t[80] = t[102] ^ x[57];
  assign t[81] = t[103] ^ x[60];
  assign t[82] = t[104] ^ x[63];
  assign t[83] = t[105] ^ x[66];
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind348(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind349(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind350(x, y);
 input [66:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = (t[142] & ~t[143]);
  assign t[103] = (t[144] & ~t[145]);
  assign t[104] = (t[146] & ~t[147]);
  assign t[105] = (t[148] & ~t[149]);
  assign t[106] = t[150] ^ x[2];
  assign t[107] = t[151] ^ x[1];
  assign t[108] = t[152] ^ x[6];
  assign t[109] = t[153] ^ x[5];
  assign t[10] = t[42] & t[15];
  assign t[110] = t[154] ^ x[9];
  assign t[111] = t[155] ^ x[8];
  assign t[112] = t[156] ^ x[12];
  assign t[113] = t[157] ^ x[11];
  assign t[114] = t[158] ^ x[15];
  assign t[115] = t[159] ^ x[14];
  assign t[116] = t[160] ^ x[18];
  assign t[117] = t[161] ^ x[17];
  assign t[118] = t[162] ^ x[21];
  assign t[119] = t[163] ^ x[20];
  assign t[11] = ~(t[16]);
  assign t[120] = t[164] ^ x[24];
  assign t[121] = t[165] ^ x[23];
  assign t[122] = t[166] ^ x[27];
  assign t[123] = t[167] ^ x[26];
  assign t[124] = t[168] ^ x[30];
  assign t[125] = t[169] ^ x[29];
  assign t[126] = t[170] ^ x[33];
  assign t[127] = t[171] ^ x[32];
  assign t[128] = t[172] ^ x[36];
  assign t[129] = t[173] ^ x[35];
  assign t[12] = ~(t[42]);
  assign t[130] = t[174] ^ x[39];
  assign t[131] = t[175] ^ x[38];
  assign t[132] = t[176] ^ x[42];
  assign t[133] = t[177] ^ x[41];
  assign t[134] = t[178] ^ x[45];
  assign t[135] = t[179] ^ x[44];
  assign t[136] = t[180] ^ x[48];
  assign t[137] = t[181] ^ x[47];
  assign t[138] = t[182] ^ x[51];
  assign t[139] = t[183] ^ x[50];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[54];
  assign t[141] = t[185] ^ x[53];
  assign t[142] = t[186] ^ x[57];
  assign t[143] = t[187] ^ x[56];
  assign t[144] = t[188] ^ x[60];
  assign t[145] = t[189] ^ x[59];
  assign t[146] = t[190] ^ x[63];
  assign t[147] = t[191] ^ x[62];
  assign t[148] = t[192] ^ x[66];
  assign t[149] = t[193] ^ x[65];
  assign t[14] = t[18] ? t[43] : t[19];
  assign t[150] = (x[0]);
  assign t[151] = (x[0]);
  assign t[152] = (x[4]);
  assign t[153] = (x[4]);
  assign t[154] = (x[7]);
  assign t[155] = (x[7]);
  assign t[156] = (x[10]);
  assign t[157] = (x[10]);
  assign t[158] = (x[13]);
  assign t[159] = (x[13]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[16]);
  assign t[161] = (x[16]);
  assign t[162] = (x[19]);
  assign t[163] = (x[19]);
  assign t[164] = (x[22]);
  assign t[165] = (x[22]);
  assign t[166] = (x[25]);
  assign t[167] = (x[25]);
  assign t[168] = (x[28]);
  assign t[169] = (x[28]);
  assign t[16] = ~(t[42] & t[22]);
  assign t[170] = (x[31]);
  assign t[171] = (x[31]);
  assign t[172] = (x[34]);
  assign t[173] = (x[34]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[40]);
  assign t[177] = (x[40]);
  assign t[178] = (x[43]);
  assign t[179] = (x[43]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[46]);
  assign t[181] = (x[46]);
  assign t[182] = (x[49]);
  assign t[183] = (x[49]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[55]);
  assign t[187] = (x[55]);
  assign t[188] = (x[58]);
  assign t[189] = (x[58]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[61]);
  assign t[191] = (x[61]);
  assign t[192] = (x[64]);
  assign t[193] = (x[64]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[44] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[40] : t[5];
  assign t[30] = ~(t[51] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[42]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[41] ^ t[39];
  assign t[36] = ~(t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = (t[82]);
  assign t[61] = (t[83]);
  assign t[62] = t[84] ^ x[2];
  assign t[63] = t[85] ^ x[6];
  assign t[64] = t[86] ^ x[9];
  assign t[65] = t[87] ^ x[12];
  assign t[66] = t[88] ^ x[15];
  assign t[67] = t[89] ^ x[18];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[24];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[27];
  assign t[71] = t[93] ^ x[30];
  assign t[72] = t[94] ^ x[33];
  assign t[73] = t[95] ^ x[36];
  assign t[74] = t[96] ^ x[39];
  assign t[75] = t[97] ^ x[42];
  assign t[76] = t[98] ^ x[45];
  assign t[77] = t[99] ^ x[48];
  assign t[78] = t[100] ^ x[51];
  assign t[79] = t[101] ^ x[54];
  assign t[7] = ~(t[11]);
  assign t[80] = t[102] ^ x[57];
  assign t[81] = t[103] ^ x[60];
  assign t[82] = t[104] ^ x[63];
  assign t[83] = t[105] ^ x[66];
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind351(x, y);
 input [66:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = (t[142] & ~t[143]);
  assign t[103] = (t[144] & ~t[145]);
  assign t[104] = (t[146] & ~t[147]);
  assign t[105] = (t[148] & ~t[149]);
  assign t[106] = t[150] ^ x[2];
  assign t[107] = t[151] ^ x[1];
  assign t[108] = t[152] ^ x[6];
  assign t[109] = t[153] ^ x[5];
  assign t[10] = t[42] & t[15];
  assign t[110] = t[154] ^ x[9];
  assign t[111] = t[155] ^ x[8];
  assign t[112] = t[156] ^ x[12];
  assign t[113] = t[157] ^ x[11];
  assign t[114] = t[158] ^ x[15];
  assign t[115] = t[159] ^ x[14];
  assign t[116] = t[160] ^ x[18];
  assign t[117] = t[161] ^ x[17];
  assign t[118] = t[162] ^ x[21];
  assign t[119] = t[163] ^ x[20];
  assign t[11] = ~(t[16]);
  assign t[120] = t[164] ^ x[24];
  assign t[121] = t[165] ^ x[23];
  assign t[122] = t[166] ^ x[27];
  assign t[123] = t[167] ^ x[26];
  assign t[124] = t[168] ^ x[30];
  assign t[125] = t[169] ^ x[29];
  assign t[126] = t[170] ^ x[33];
  assign t[127] = t[171] ^ x[32];
  assign t[128] = t[172] ^ x[36];
  assign t[129] = t[173] ^ x[35];
  assign t[12] = ~(t[42]);
  assign t[130] = t[174] ^ x[39];
  assign t[131] = t[175] ^ x[38];
  assign t[132] = t[176] ^ x[42];
  assign t[133] = t[177] ^ x[41];
  assign t[134] = t[178] ^ x[45];
  assign t[135] = t[179] ^ x[44];
  assign t[136] = t[180] ^ x[48];
  assign t[137] = t[181] ^ x[47];
  assign t[138] = t[182] ^ x[51];
  assign t[139] = t[183] ^ x[50];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[54];
  assign t[141] = t[185] ^ x[53];
  assign t[142] = t[186] ^ x[57];
  assign t[143] = t[187] ^ x[56];
  assign t[144] = t[188] ^ x[60];
  assign t[145] = t[189] ^ x[59];
  assign t[146] = t[190] ^ x[63];
  assign t[147] = t[191] ^ x[62];
  assign t[148] = t[192] ^ x[66];
  assign t[149] = t[193] ^ x[65];
  assign t[14] = t[18] ? t[43] : t[19];
  assign t[150] = (x[0]);
  assign t[151] = (x[0]);
  assign t[152] = (x[4]);
  assign t[153] = (x[4]);
  assign t[154] = (x[7]);
  assign t[155] = (x[7]);
  assign t[156] = (x[10]);
  assign t[157] = (x[10]);
  assign t[158] = (x[13]);
  assign t[159] = (x[13]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[16]);
  assign t[161] = (x[16]);
  assign t[162] = (x[19]);
  assign t[163] = (x[19]);
  assign t[164] = (x[22]);
  assign t[165] = (x[22]);
  assign t[166] = (x[25]);
  assign t[167] = (x[25]);
  assign t[168] = (x[28]);
  assign t[169] = (x[28]);
  assign t[16] = ~(t[42] & t[22]);
  assign t[170] = (x[31]);
  assign t[171] = (x[31]);
  assign t[172] = (x[34]);
  assign t[173] = (x[34]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[40]);
  assign t[177] = (x[40]);
  assign t[178] = (x[43]);
  assign t[179] = (x[43]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[46]);
  assign t[181] = (x[46]);
  assign t[182] = (x[49]);
  assign t[183] = (x[49]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[55]);
  assign t[187] = (x[55]);
  assign t[188] = (x[58]);
  assign t[189] = (x[58]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[61]);
  assign t[191] = (x[61]);
  assign t[192] = (x[64]);
  assign t[193] = (x[64]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[44] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[40] : t[5];
  assign t[30] = ~(t[51] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[42]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[41] ^ t[39];
  assign t[36] = ~(t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = (t[82]);
  assign t[61] = (t[83]);
  assign t[62] = t[84] ^ x[2];
  assign t[63] = t[85] ^ x[6];
  assign t[64] = t[86] ^ x[9];
  assign t[65] = t[87] ^ x[12];
  assign t[66] = t[88] ^ x[15];
  assign t[67] = t[89] ^ x[18];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[24];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[27];
  assign t[71] = t[93] ^ x[30];
  assign t[72] = t[94] ^ x[33];
  assign t[73] = t[95] ^ x[36];
  assign t[74] = t[96] ^ x[39];
  assign t[75] = t[97] ^ x[42];
  assign t[76] = t[98] ^ x[45];
  assign t[77] = t[99] ^ x[48];
  assign t[78] = t[100] ^ x[51];
  assign t[79] = t[101] ^ x[54];
  assign t[7] = ~(t[11]);
  assign t[80] = t[102] ^ x[57];
  assign t[81] = t[103] ^ x[60];
  assign t[82] = t[104] ^ x[63];
  assign t[83] = t[105] ^ x[66];
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind352(x, y);
 input [66:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = (t[142] & ~t[143]);
  assign t[103] = (t[144] & ~t[145]);
  assign t[104] = (t[146] & ~t[147]);
  assign t[105] = (t[148] & ~t[149]);
  assign t[106] = t[150] ^ x[2];
  assign t[107] = t[151] ^ x[1];
  assign t[108] = t[152] ^ x[6];
  assign t[109] = t[153] ^ x[5];
  assign t[10] = t[42] & t[15];
  assign t[110] = t[154] ^ x[9];
  assign t[111] = t[155] ^ x[8];
  assign t[112] = t[156] ^ x[12];
  assign t[113] = t[157] ^ x[11];
  assign t[114] = t[158] ^ x[15];
  assign t[115] = t[159] ^ x[14];
  assign t[116] = t[160] ^ x[18];
  assign t[117] = t[161] ^ x[17];
  assign t[118] = t[162] ^ x[21];
  assign t[119] = t[163] ^ x[20];
  assign t[11] = ~(t[16]);
  assign t[120] = t[164] ^ x[24];
  assign t[121] = t[165] ^ x[23];
  assign t[122] = t[166] ^ x[27];
  assign t[123] = t[167] ^ x[26];
  assign t[124] = t[168] ^ x[30];
  assign t[125] = t[169] ^ x[29];
  assign t[126] = t[170] ^ x[33];
  assign t[127] = t[171] ^ x[32];
  assign t[128] = t[172] ^ x[36];
  assign t[129] = t[173] ^ x[35];
  assign t[12] = ~(t[42]);
  assign t[130] = t[174] ^ x[39];
  assign t[131] = t[175] ^ x[38];
  assign t[132] = t[176] ^ x[42];
  assign t[133] = t[177] ^ x[41];
  assign t[134] = t[178] ^ x[45];
  assign t[135] = t[179] ^ x[44];
  assign t[136] = t[180] ^ x[48];
  assign t[137] = t[181] ^ x[47];
  assign t[138] = t[182] ^ x[51];
  assign t[139] = t[183] ^ x[50];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[54];
  assign t[141] = t[185] ^ x[53];
  assign t[142] = t[186] ^ x[57];
  assign t[143] = t[187] ^ x[56];
  assign t[144] = t[188] ^ x[60];
  assign t[145] = t[189] ^ x[59];
  assign t[146] = t[190] ^ x[63];
  assign t[147] = t[191] ^ x[62];
  assign t[148] = t[192] ^ x[66];
  assign t[149] = t[193] ^ x[65];
  assign t[14] = t[18] ? t[43] : t[19];
  assign t[150] = (x[0]);
  assign t[151] = (x[0]);
  assign t[152] = (x[4]);
  assign t[153] = (x[4]);
  assign t[154] = (x[7]);
  assign t[155] = (x[7]);
  assign t[156] = (x[10]);
  assign t[157] = (x[10]);
  assign t[158] = (x[13]);
  assign t[159] = (x[13]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[16]);
  assign t[161] = (x[16]);
  assign t[162] = (x[19]);
  assign t[163] = (x[19]);
  assign t[164] = (x[22]);
  assign t[165] = (x[22]);
  assign t[166] = (x[25]);
  assign t[167] = (x[25]);
  assign t[168] = (x[28]);
  assign t[169] = (x[28]);
  assign t[16] = ~(t[42] & t[22]);
  assign t[170] = (x[31]);
  assign t[171] = (x[31]);
  assign t[172] = (x[34]);
  assign t[173] = (x[34]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[40]);
  assign t[177] = (x[40]);
  assign t[178] = (x[43]);
  assign t[179] = (x[43]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[46]);
  assign t[181] = (x[46]);
  assign t[182] = (x[49]);
  assign t[183] = (x[49]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[55]);
  assign t[187] = (x[55]);
  assign t[188] = (x[58]);
  assign t[189] = (x[58]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[61]);
  assign t[191] = (x[61]);
  assign t[192] = (x[64]);
  assign t[193] = (x[64]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[44] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[40] : t[5];
  assign t[30] = ~(t[51] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[42]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[41] ^ t[39];
  assign t[36] = ~(t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = (t[82]);
  assign t[61] = (t[83]);
  assign t[62] = t[84] ^ x[2];
  assign t[63] = t[85] ^ x[6];
  assign t[64] = t[86] ^ x[9];
  assign t[65] = t[87] ^ x[12];
  assign t[66] = t[88] ^ x[15];
  assign t[67] = t[89] ^ x[18];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[24];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[27];
  assign t[71] = t[93] ^ x[30];
  assign t[72] = t[94] ^ x[33];
  assign t[73] = t[95] ^ x[36];
  assign t[74] = t[96] ^ x[39];
  assign t[75] = t[97] ^ x[42];
  assign t[76] = t[98] ^ x[45];
  assign t[77] = t[99] ^ x[48];
  assign t[78] = t[100] ^ x[51];
  assign t[79] = t[101] ^ x[54];
  assign t[7] = ~(t[11]);
  assign t[80] = t[102] ^ x[57];
  assign t[81] = t[103] ^ x[60];
  assign t[82] = t[104] ^ x[63];
  assign t[83] = t[105] ^ x[66];
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind353(x, y);
 input [66:0] x;
 output y;

 wire [193:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[138] & ~t[139]);
  assign t[101] = (t[140] & ~t[141]);
  assign t[102] = (t[142] & ~t[143]);
  assign t[103] = (t[144] & ~t[145]);
  assign t[104] = (t[146] & ~t[147]);
  assign t[105] = (t[148] & ~t[149]);
  assign t[106] = t[150] ^ x[2];
  assign t[107] = t[151] ^ x[1];
  assign t[108] = t[152] ^ x[6];
  assign t[109] = t[153] ^ x[5];
  assign t[10] = t[42] & t[15];
  assign t[110] = t[154] ^ x[9];
  assign t[111] = t[155] ^ x[8];
  assign t[112] = t[156] ^ x[12];
  assign t[113] = t[157] ^ x[11];
  assign t[114] = t[158] ^ x[15];
  assign t[115] = t[159] ^ x[14];
  assign t[116] = t[160] ^ x[18];
  assign t[117] = t[161] ^ x[17];
  assign t[118] = t[162] ^ x[21];
  assign t[119] = t[163] ^ x[20];
  assign t[11] = ~(t[16]);
  assign t[120] = t[164] ^ x[24];
  assign t[121] = t[165] ^ x[23];
  assign t[122] = t[166] ^ x[27];
  assign t[123] = t[167] ^ x[26];
  assign t[124] = t[168] ^ x[30];
  assign t[125] = t[169] ^ x[29];
  assign t[126] = t[170] ^ x[33];
  assign t[127] = t[171] ^ x[32];
  assign t[128] = t[172] ^ x[36];
  assign t[129] = t[173] ^ x[35];
  assign t[12] = ~(t[42]);
  assign t[130] = t[174] ^ x[39];
  assign t[131] = t[175] ^ x[38];
  assign t[132] = t[176] ^ x[42];
  assign t[133] = t[177] ^ x[41];
  assign t[134] = t[178] ^ x[45];
  assign t[135] = t[179] ^ x[44];
  assign t[136] = t[180] ^ x[48];
  assign t[137] = t[181] ^ x[47];
  assign t[138] = t[182] ^ x[51];
  assign t[139] = t[183] ^ x[50];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[54];
  assign t[141] = t[185] ^ x[53];
  assign t[142] = t[186] ^ x[57];
  assign t[143] = t[187] ^ x[56];
  assign t[144] = t[188] ^ x[60];
  assign t[145] = t[189] ^ x[59];
  assign t[146] = t[190] ^ x[63];
  assign t[147] = t[191] ^ x[62];
  assign t[148] = t[192] ^ x[66];
  assign t[149] = t[193] ^ x[65];
  assign t[14] = t[18] ? t[43] : t[19];
  assign t[150] = (x[0]);
  assign t[151] = (x[0]);
  assign t[152] = (x[4]);
  assign t[153] = (x[4]);
  assign t[154] = (x[7]);
  assign t[155] = (x[7]);
  assign t[156] = (x[10]);
  assign t[157] = (x[10]);
  assign t[158] = (x[13]);
  assign t[159] = (x[13]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[16]);
  assign t[161] = (x[16]);
  assign t[162] = (x[19]);
  assign t[163] = (x[19]);
  assign t[164] = (x[22]);
  assign t[165] = (x[22]);
  assign t[166] = (x[25]);
  assign t[167] = (x[25]);
  assign t[168] = (x[28]);
  assign t[169] = (x[28]);
  assign t[16] = ~(t[42] & t[22]);
  assign t[170] = (x[31]);
  assign t[171] = (x[31]);
  assign t[172] = (x[34]);
  assign t[173] = (x[34]);
  assign t[174] = (x[37]);
  assign t[175] = (x[37]);
  assign t[176] = (x[40]);
  assign t[177] = (x[40]);
  assign t[178] = (x[43]);
  assign t[179] = (x[43]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[46]);
  assign t[181] = (x[46]);
  assign t[182] = (x[49]);
  assign t[183] = (x[49]);
  assign t[184] = (x[52]);
  assign t[185] = (x[52]);
  assign t[186] = (x[55]);
  assign t[187] = (x[55]);
  assign t[188] = (x[58]);
  assign t[189] = (x[58]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[61]);
  assign t[191] = (x[61]);
  assign t[192] = (x[64]);
  assign t[193] = (x[64]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[44] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[40] : t[5];
  assign t[30] = ~(t[51] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[42]);
  assign t[34] = t[53] ^ t[54];
  assign t[35] = t[41] ^ t[39];
  assign t[36] = ~(t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = ~(t[58] | t[59]);
  assign t[39] = t[60] ^ t[61];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = (t[82]);
  assign t[61] = (t[83]);
  assign t[62] = t[84] ^ x[2];
  assign t[63] = t[85] ^ x[6];
  assign t[64] = t[86] ^ x[9];
  assign t[65] = t[87] ^ x[12];
  assign t[66] = t[88] ^ x[15];
  assign t[67] = t[89] ^ x[18];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[24];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[27];
  assign t[71] = t[93] ^ x[30];
  assign t[72] = t[94] ^ x[33];
  assign t[73] = t[95] ^ x[36];
  assign t[74] = t[96] ^ x[39];
  assign t[75] = t[97] ^ x[42];
  assign t[76] = t[98] ^ x[45];
  assign t[77] = t[99] ^ x[48];
  assign t[78] = t[100] ^ x[51];
  assign t[79] = t[101] ^ x[54];
  assign t[7] = ~(t[11]);
  assign t[80] = t[102] ^ x[57];
  assign t[81] = t[103] ^ x[60];
  assign t[82] = t[104] ^ x[63];
  assign t[83] = t[105] ^ x[66];
  assign t[84] = (t[106] & ~t[107]);
  assign t[85] = (t[108] & ~t[109]);
  assign t[86] = (t[110] & ~t[111]);
  assign t[87] = (t[112] & ~t[113]);
  assign t[88] = (t[114] & ~t[115]);
  assign t[89] = (t[116] & ~t[117]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[118] & ~t[119]);
  assign t[91] = (t[120] & ~t[121]);
  assign t[92] = (t[122] & ~t[123]);
  assign t[93] = (t[124] & ~t[125]);
  assign t[94] = (t[126] & ~t[127]);
  assign t[95] = (t[128] & ~t[129]);
  assign t[96] = (t[130] & ~t[131]);
  assign t[97] = (t[132] & ~t[133]);
  assign t[98] = (t[134] & ~t[135]);
  assign t[99] = (t[136] & ~t[137]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind354(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind355(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind356(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind357(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind358(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind359(x, y);
 input [60:0] x;
 output y;

 wire [177:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = t[140] ^ x[6];
  assign t[101] = t[141] ^ x[5];
  assign t[102] = t[142] ^ x[9];
  assign t[103] = t[143] ^ x[8];
  assign t[104] = t[144] ^ x[12];
  assign t[105] = t[145] ^ x[11];
  assign t[106] = t[146] ^ x[15];
  assign t[107] = t[147] ^ x[14];
  assign t[108] = t[148] ^ x[18];
  assign t[109] = t[149] ^ x[17];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[150] ^ x[21];
  assign t[111] = t[151] ^ x[20];
  assign t[112] = t[152] ^ x[24];
  assign t[113] = t[153] ^ x[23];
  assign t[114] = t[154] ^ x[27];
  assign t[115] = t[155] ^ x[26];
  assign t[116] = t[156] ^ x[30];
  assign t[117] = t[157] ^ x[29];
  assign t[118] = t[158] ^ x[33];
  assign t[119] = t[159] ^ x[32];
  assign t[11] = ~(t[16]);
  assign t[120] = t[160] ^ x[36];
  assign t[121] = t[161] ^ x[35];
  assign t[122] = t[162] ^ x[39];
  assign t[123] = t[163] ^ x[38];
  assign t[124] = t[164] ^ x[42];
  assign t[125] = t[165] ^ x[41];
  assign t[126] = t[166] ^ x[45];
  assign t[127] = t[167] ^ x[44];
  assign t[128] = t[168] ^ x[48];
  assign t[129] = t[169] ^ x[47];
  assign t[12] = ~(t[40]);
  assign t[130] = t[170] ^ x[51];
  assign t[131] = t[171] ^ x[50];
  assign t[132] = t[172] ^ x[54];
  assign t[133] = t[173] ^ x[53];
  assign t[134] = t[174] ^ x[57];
  assign t[135] = t[175] ^ x[56];
  assign t[136] = t[176] ^ x[60];
  assign t[137] = t[177] ^ x[59];
  assign t[138] = (x[0]);
  assign t[139] = (x[0]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[4]);
  assign t[141] = (x[4]);
  assign t[142] = (x[7]);
  assign t[143] = (x[7]);
  assign t[144] = (x[10]);
  assign t[145] = (x[10]);
  assign t[146] = (x[13]);
  assign t[147] = (x[13]);
  assign t[148] = (x[16]);
  assign t[149] = (x[16]);
  assign t[14] = t[18] ? t[41] : t[19];
  assign t[150] = (x[19]);
  assign t[151] = (x[19]);
  assign t[152] = (x[22]);
  assign t[153] = (x[22]);
  assign t[154] = (x[25]);
  assign t[155] = (x[25]);
  assign t[156] = (x[28]);
  assign t[157] = (x[28]);
  assign t[158] = (x[31]);
  assign t[159] = (x[31]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[34]);
  assign t[161] = (x[34]);
  assign t[162] = (x[37]);
  assign t[163] = (x[37]);
  assign t[164] = (x[40]);
  assign t[165] = (x[40]);
  assign t[166] = (x[43]);
  assign t[167] = (x[43]);
  assign t[168] = (x[46]);
  assign t[169] = (x[46]);
  assign t[16] = ~(t[40] & t[22]);
  assign t[170] = (x[49]);
  assign t[171] = (x[49]);
  assign t[172] = (x[52]);
  assign t[173] = (x[52]);
  assign t[174] = (x[55]);
  assign t[175] = (x[55]);
  assign t[176] = (x[58]);
  assign t[177] = (x[58]);
  assign t[17] = ~(t[23]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[42] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[43] ^ t[34];
  assign t[26] = ~(t[44] ^ t[45]);
  assign t[27] = ~(t[46] & t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[38] : t[5];
  assign t[30] = ~(t[50] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[51]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[39] ^ t[52];
  assign t[35] = ~(t[53]);
  assign t[36] = ~(t[54] | t[55]);
  assign t[37] = ~(t[56] | t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = (t[76]);
  assign t[57] = (t[77]);
  assign t[58] = t[78] ^ x[2];
  assign t[59] = t[79] ^ x[6];
  assign t[5] = t[8] ? t[9] : x[3];
  assign t[60] = t[80] ^ x[9];
  assign t[61] = t[81] ^ x[12];
  assign t[62] = t[82] ^ x[15];
  assign t[63] = t[83] ^ x[18];
  assign t[64] = t[84] ^ x[21];
  assign t[65] = t[85] ^ x[24];
  assign t[66] = t[86] ^ x[27];
  assign t[67] = t[87] ^ x[30];
  assign t[68] = t[88] ^ x[33];
  assign t[69] = t[89] ^ x[36];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[39];
  assign t[71] = t[91] ^ x[42];
  assign t[72] = t[92] ^ x[45];
  assign t[73] = t[93] ^ x[48];
  assign t[74] = t[94] ^ x[51];
  assign t[75] = t[95] ^ x[54];
  assign t[76] = t[96] ^ x[57];
  assign t[77] = t[97] ^ x[60];
  assign t[78] = (t[98] & ~t[99]);
  assign t[79] = (t[100] & ~t[101]);
  assign t[7] = ~(t[11]);
  assign t[80] = (t[102] & ~t[103]);
  assign t[81] = (t[104] & ~t[105]);
  assign t[82] = (t[106] & ~t[107]);
  assign t[83] = (t[108] & ~t[109]);
  assign t[84] = (t[110] & ~t[111]);
  assign t[85] = (t[112] & ~t[113]);
  assign t[86] = (t[114] & ~t[115]);
  assign t[87] = (t[116] & ~t[117]);
  assign t[88] = (t[118] & ~t[119]);
  assign t[89] = (t[120] & ~t[121]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[122] & ~t[123]);
  assign t[91] = (t[124] & ~t[125]);
  assign t[92] = (t[126] & ~t[127]);
  assign t[93] = (t[128] & ~t[129]);
  assign t[94] = (t[130] & ~t[131]);
  assign t[95] = (t[132] & ~t[133]);
  assign t[96] = (t[134] & ~t[135]);
  assign t[97] = (t[136] & ~t[137]);
  assign t[98] = t[138] ^ x[2];
  assign t[99] = t[139] ^ x[1];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind360(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind361(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind362(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind363(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind364(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind365(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind366(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind367(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind368(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind369(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind370(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind371(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind372(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind373(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind374(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind375(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind376(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind377(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind378(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind379(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind380(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind381(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind382(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind383(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind384(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind385(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind386(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind387(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind388(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind389(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind390(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind391(x, y);
 input [42:0] x;
 output y;

 wire [122:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[7]);
  assign t[101] = (x[10]);
  assign t[102] = (x[10]);
  assign t[103] = (x[13]);
  assign t[104] = (x[13]);
  assign t[105] = (x[16]);
  assign t[106] = (x[16]);
  assign t[107] = (x[19]);
  assign t[108] = (x[19]);
  assign t[109] = (x[22]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[22]);
  assign t[111] = (x[25]);
  assign t[112] = (x[25]);
  assign t[113] = (x[28]);
  assign t[114] = (x[28]);
  assign t[115] = (x[31]);
  assign t[116] = (x[31]);
  assign t[117] = (x[34]);
  assign t[118] = (x[34]);
  assign t[119] = (x[37]);
  assign t[11] = ~(t[27]);
  assign t[120] = (x[37]);
  assign t[121] = (x[40]);
  assign t[122] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[27] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[28] | t[21]);
  assign t[17] = ~(t[29] & t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[33] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[35] | t[36]);
  assign t[24] = ~(t[37] | t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = t[53] ^ x[2];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[5];
  assign t[41] = t[55] ^ x[9];
  assign t[42] = t[56] ^ x[12];
  assign t[43] = t[57] ^ x[15];
  assign t[44] = t[58] ^ x[18];
  assign t[45] = t[59] ^ x[21];
  assign t[46] = t[60] ^ x[24];
  assign t[47] = t[61] ^ x[27];
  assign t[48] = t[62] ^ x[30];
  assign t[49] = t[63] ^ x[33];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[36];
  assign t[51] = t[65] ^ x[39];
  assign t[52] = t[66] ^ x[42];
  assign t[53] = (t[67] & ~t[68]);
  assign t[54] = (t[69] & ~t[70]);
  assign t[55] = (t[71] & ~t[72]);
  assign t[56] = (t[73] & ~t[74]);
  assign t[57] = (t[75] & ~t[76]);
  assign t[58] = (t[77] & ~t[78]);
  assign t[59] = (t[79] & ~t[80]);
  assign t[5] = t[8] ? t[26] : x[6];
  assign t[60] = (t[81] & ~t[82]);
  assign t[61] = (t[83] & ~t[84]);
  assign t[62] = (t[85] & ~t[86]);
  assign t[63] = (t[87] & ~t[88]);
  assign t[64] = (t[89] & ~t[90]);
  assign t[65] = (t[91] & ~t[92]);
  assign t[66] = (t[93] & ~t[94]);
  assign t[67] = t[95] ^ x[2];
  assign t[68] = t[96] ^ x[1];
  assign t[69] = t[97] ^ x[5];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[4];
  assign t[71] = t[99] ^ x[9];
  assign t[72] = t[100] ^ x[8];
  assign t[73] = t[101] ^ x[12];
  assign t[74] = t[102] ^ x[11];
  assign t[75] = t[103] ^ x[15];
  assign t[76] = t[104] ^ x[14];
  assign t[77] = t[105] ^ x[18];
  assign t[78] = t[106] ^ x[17];
  assign t[79] = t[107] ^ x[21];
  assign t[7] = ~(t[10]);
  assign t[80] = t[108] ^ x[20];
  assign t[81] = t[109] ^ x[24];
  assign t[82] = t[110] ^ x[23];
  assign t[83] = t[111] ^ x[27];
  assign t[84] = t[112] ^ x[26];
  assign t[85] = t[113] ^ x[30];
  assign t[86] = t[114] ^ x[29];
  assign t[87] = t[115] ^ x[33];
  assign t[88] = t[116] ^ x[32];
  assign t[89] = t[117] ^ x[36];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[35];
  assign t[91] = t[119] ^ x[39];
  assign t[92] = t[120] ^ x[38];
  assign t[93] = t[121] ^ x[42];
  assign t[94] = t[122] ^ x[41];
  assign t[95] = (x[0]);
  assign t[96] = (x[0]);
  assign t[97] = (x[3]);
  assign t[98] = (x[3]);
  assign t[99] = (x[7]);
  assign t[9] = t[27] & t[12];
  assign y = (t[0]);
endmodule

module R2ind392(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind393(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind394(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind395(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind396(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind397(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind398(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind399(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind400(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind401(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind402(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind403(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind404(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind405(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind406(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind407(x, y);
 input [42:0] x;
 output y;

 wire [120:0] t;
  assign t[0] = t[1] ? t[2] : t[23];
  assign t[100] = (x[10]);
  assign t[101] = (x[13]);
  assign t[102] = (x[13]);
  assign t[103] = (x[16]);
  assign t[104] = (x[16]);
  assign t[105] = (x[19]);
  assign t[106] = (x[19]);
  assign t[107] = (x[22]);
  assign t[108] = (x[22]);
  assign t[109] = (x[25]);
  assign t[10] = ~(t[26] | t[13]);
  assign t[110] = (x[25]);
  assign t[111] = (x[28]);
  assign t[112] = (x[28]);
  assign t[113] = (x[31]);
  assign t[114] = (x[31]);
  assign t[115] = (x[34]);
  assign t[116] = (x[34]);
  assign t[117] = (x[37]);
  assign t[118] = (x[37]);
  assign t[119] = (x[40]);
  assign t[11] = ~(t[25]);
  assign t[120] = (x[40]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[16] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = ~(t[20] | t[21]);
  assign t[16] = ~(t[27] | t[28]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[31] & t[32]);
  assign t[19] = ~(t[33] & t[34]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[10]);
  assign t[21] = ~(t[35] & t[22]);
  assign t[22] = ~(t[36]);
  assign t[23] = (t[37]);
  assign t[24] = (t[38]);
  assign t[25] = (t[39]);
  assign t[26] = (t[40]);
  assign t[27] = (t[41]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = t[4] ? t[24] : t[5];
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = t[51] ^ x[2];
  assign t[38] = t[52] ^ x[5];
  assign t[39] = t[53] ^ x[9];
  assign t[3] = ~(t[6]);
  assign t[40] = t[54] ^ x[12];
  assign t[41] = t[55] ^ x[15];
  assign t[42] = t[56] ^ x[18];
  assign t[43] = t[57] ^ x[21];
  assign t[44] = t[58] ^ x[24];
  assign t[45] = t[59] ^ x[27];
  assign t[46] = t[60] ^ x[30];
  assign t[47] = t[61] ^ x[33];
  assign t[48] = t[62] ^ x[36];
  assign t[49] = t[63] ^ x[39];
  assign t[4] = ~(t[7]);
  assign t[50] = t[64] ^ x[42];
  assign t[51] = (t[65] & ~t[66]);
  assign t[52] = (t[67] & ~t[68]);
  assign t[53] = (t[69] & ~t[70]);
  assign t[54] = (t[71] & ~t[72]);
  assign t[55] = (t[73] & ~t[74]);
  assign t[56] = (t[75] & ~t[76]);
  assign t[57] = (t[77] & ~t[78]);
  assign t[58] = (t[79] & ~t[80]);
  assign t[59] = (t[81] & ~t[82]);
  assign t[5] = t[8] ? t[24] : x[6];
  assign t[60] = (t[83] & ~t[84]);
  assign t[61] = (t[85] & ~t[86]);
  assign t[62] = (t[87] & ~t[88]);
  assign t[63] = (t[89] & ~t[90]);
  assign t[64] = (t[91] & ~t[92]);
  assign t[65] = t[93] ^ x[2];
  assign t[66] = t[94] ^ x[1];
  assign t[67] = t[95] ^ x[5];
  assign t[68] = t[96] ^ x[4];
  assign t[69] = t[97] ^ x[9];
  assign t[6] = ~(t[9]);
  assign t[70] = t[98] ^ x[8];
  assign t[71] = t[99] ^ x[12];
  assign t[72] = t[100] ^ x[11];
  assign t[73] = t[101] ^ x[15];
  assign t[74] = t[102] ^ x[14];
  assign t[75] = t[103] ^ x[18];
  assign t[76] = t[104] ^ x[17];
  assign t[77] = t[105] ^ x[21];
  assign t[78] = t[106] ^ x[20];
  assign t[79] = t[107] ^ x[24];
  assign t[7] = ~(t[25] & t[10]);
  assign t[80] = t[108] ^ x[23];
  assign t[81] = t[109] ^ x[27];
  assign t[82] = t[110] ^ x[26];
  assign t[83] = t[111] ^ x[30];
  assign t[84] = t[112] ^ x[29];
  assign t[85] = t[113] ^ x[33];
  assign t[86] = t[114] ^ x[32];
  assign t[87] = t[115] ^ x[36];
  assign t[88] = t[116] ^ x[35];
  assign t[89] = t[117] ^ x[39];
  assign t[8] = ~(t[11]);
  assign t[90] = t[118] ^ x[38];
  assign t[91] = t[119] ^ x[42];
  assign t[92] = t[120] ^ x[41];
  assign t[93] = (x[0]);
  assign t[94] = (x[0]);
  assign t[95] = (x[3]);
  assign t[96] = (x[3]);
  assign t[97] = (x[7]);
  assign t[98] = (x[7]);
  assign t[99] = (x[10]);
  assign t[9] = t[25] & t[12];
  assign y = (t[0]);
endmodule

module R2ind408(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind409(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind410(x, y);
 input [66:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[140] & ~t[141]);
  assign t[101] = (t[142] & ~t[143]);
  assign t[102] = (t[144] & ~t[145]);
  assign t[103] = (t[146] & ~t[147]);
  assign t[104] = t[148] ^ x[2];
  assign t[105] = t[149] ^ x[1];
  assign t[106] = t[150] ^ x[5];
  assign t[107] = t[151] ^ x[4];
  assign t[108] = t[152] ^ x[9];
  assign t[109] = t[153] ^ x[8];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[154] ^ x[12];
  assign t[111] = t[155] ^ x[11];
  assign t[112] = t[156] ^ x[15];
  assign t[113] = t[157] ^ x[14];
  assign t[114] = t[158] ^ x[18];
  assign t[115] = t[159] ^ x[17];
  assign t[116] = t[160] ^ x[21];
  assign t[117] = t[161] ^ x[20];
  assign t[118] = t[162] ^ x[24];
  assign t[119] = t[163] ^ x[23];
  assign t[11] = ~(t[42] | t[16]);
  assign t[120] = t[164] ^ x[27];
  assign t[121] = t[165] ^ x[26];
  assign t[122] = t[166] ^ x[30];
  assign t[123] = t[167] ^ x[29];
  assign t[124] = t[168] ^ x[33];
  assign t[125] = t[169] ^ x[32];
  assign t[126] = t[170] ^ x[36];
  assign t[127] = t[171] ^ x[35];
  assign t[128] = t[172] ^ x[39];
  assign t[129] = t[173] ^ x[38];
  assign t[12] = ~(t[40]);
  assign t[130] = t[174] ^ x[42];
  assign t[131] = t[175] ^ x[41];
  assign t[132] = t[176] ^ x[45];
  assign t[133] = t[177] ^ x[44];
  assign t[134] = t[178] ^ x[48];
  assign t[135] = t[179] ^ x[47];
  assign t[136] = t[180] ^ x[51];
  assign t[137] = t[181] ^ x[50];
  assign t[138] = t[182] ^ x[54];
  assign t[139] = t[183] ^ x[53];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[57];
  assign t[141] = t[185] ^ x[56];
  assign t[142] = t[186] ^ x[60];
  assign t[143] = t[187] ^ x[59];
  assign t[144] = t[188] ^ x[63];
  assign t[145] = t[189] ^ x[62];
  assign t[146] = t[190] ^ x[66];
  assign t[147] = t[191] ^ x[65];
  assign t[148] = (x[0]);
  assign t[149] = (x[0]);
  assign t[14] = t[18] ? t[39] : t[19];
  assign t[150] = (x[3]);
  assign t[151] = (x[3]);
  assign t[152] = (x[7]);
  assign t[153] = (x[7]);
  assign t[154] = (x[10]);
  assign t[155] = (x[10]);
  assign t[156] = (x[13]);
  assign t[157] = (x[13]);
  assign t[158] = (x[16]);
  assign t[159] = (x[16]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[19]);
  assign t[161] = (x[19]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[25]);
  assign t[165] = (x[25]);
  assign t[166] = (x[28]);
  assign t[167] = (x[28]);
  assign t[168] = (x[31]);
  assign t[169] = (x[31]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[34]);
  assign t[171] = (x[34]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[40]);
  assign t[175] = (x[40]);
  assign t[176] = (x[43]);
  assign t[177] = (x[43]);
  assign t[178] = (x[46]);
  assign t[179] = (x[46]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[49]);
  assign t[181] = (x[49]);
  assign t[182] = (x[52]);
  assign t[183] = (x[52]);
  assign t[184] = (x[55]);
  assign t[185] = (x[55]);
  assign t[186] = (x[58]);
  assign t[187] = (x[58]);
  assign t[188] = (x[61]);
  assign t[189] = (x[61]);
  assign t[18] = ~(t[25]);
  assign t[190] = (x[64]);
  assign t[191] = (x[64]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[43] | t[44]);
  assign t[23] = ~(t[45] | t[46]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[34] ^ t[35];
  assign t[27] = ~(t[47] ^ t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[53] & t[36]);
  assign t[32] = ~(t[54]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[55] ^ t[56];
  assign t[35] = t[41] ^ t[37];
  assign t[36] = ~(t[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[38] = (t[60]);
  assign t[39] = (t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[82] ^ x[2];
  assign t[61] = t[83] ^ x[5];
  assign t[62] = t[84] ^ x[9];
  assign t[63] = t[85] ^ x[12];
  assign t[64] = t[86] ^ x[15];
  assign t[65] = t[87] ^ x[18];
  assign t[66] = t[88] ^ x[21];
  assign t[67] = t[89] ^ x[24];
  assign t[68] = t[90] ^ x[27];
  assign t[69] = t[91] ^ x[30];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[33];
  assign t[71] = t[93] ^ x[36];
  assign t[72] = t[94] ^ x[39];
  assign t[73] = t[95] ^ x[42];
  assign t[74] = t[96] ^ x[45];
  assign t[75] = t[97] ^ x[48];
  assign t[76] = t[98] ^ x[51];
  assign t[77] = t[99] ^ x[54];
  assign t[78] = t[100] ^ x[57];
  assign t[79] = t[101] ^ x[60];
  assign t[7] = ~(t[40] & t[11]);
  assign t[80] = t[102] ^ x[63];
  assign t[81] = t[103] ^ x[66];
  assign t[82] = (t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[107]);
  assign t[84] = (t[108] & ~t[109]);
  assign t[85] = (t[110] & ~t[111]);
  assign t[86] = (t[112] & ~t[113]);
  assign t[87] = (t[114] & ~t[115]);
  assign t[88] = (t[116] & ~t[117]);
  assign t[89] = (t[118] & ~t[119]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[120] & ~t[121]);
  assign t[91] = (t[122] & ~t[123]);
  assign t[92] = (t[124] & ~t[125]);
  assign t[93] = (t[126] & ~t[127]);
  assign t[94] = (t[128] & ~t[129]);
  assign t[95] = (t[130] & ~t[131]);
  assign t[96] = (t[132] & ~t[133]);
  assign t[97] = (t[134] & ~t[135]);
  assign t[98] = (t[136] & ~t[137]);
  assign t[99] = (t[138] & ~t[139]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind411(x, y);
 input [66:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[140] & ~t[141]);
  assign t[101] = (t[142] & ~t[143]);
  assign t[102] = (t[144] & ~t[145]);
  assign t[103] = (t[146] & ~t[147]);
  assign t[104] = t[148] ^ x[2];
  assign t[105] = t[149] ^ x[1];
  assign t[106] = t[150] ^ x[5];
  assign t[107] = t[151] ^ x[4];
  assign t[108] = t[152] ^ x[9];
  assign t[109] = t[153] ^ x[8];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[154] ^ x[12];
  assign t[111] = t[155] ^ x[11];
  assign t[112] = t[156] ^ x[15];
  assign t[113] = t[157] ^ x[14];
  assign t[114] = t[158] ^ x[18];
  assign t[115] = t[159] ^ x[17];
  assign t[116] = t[160] ^ x[21];
  assign t[117] = t[161] ^ x[20];
  assign t[118] = t[162] ^ x[24];
  assign t[119] = t[163] ^ x[23];
  assign t[11] = ~(t[42] | t[16]);
  assign t[120] = t[164] ^ x[27];
  assign t[121] = t[165] ^ x[26];
  assign t[122] = t[166] ^ x[30];
  assign t[123] = t[167] ^ x[29];
  assign t[124] = t[168] ^ x[33];
  assign t[125] = t[169] ^ x[32];
  assign t[126] = t[170] ^ x[36];
  assign t[127] = t[171] ^ x[35];
  assign t[128] = t[172] ^ x[39];
  assign t[129] = t[173] ^ x[38];
  assign t[12] = ~(t[40]);
  assign t[130] = t[174] ^ x[42];
  assign t[131] = t[175] ^ x[41];
  assign t[132] = t[176] ^ x[45];
  assign t[133] = t[177] ^ x[44];
  assign t[134] = t[178] ^ x[48];
  assign t[135] = t[179] ^ x[47];
  assign t[136] = t[180] ^ x[51];
  assign t[137] = t[181] ^ x[50];
  assign t[138] = t[182] ^ x[54];
  assign t[139] = t[183] ^ x[53];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[57];
  assign t[141] = t[185] ^ x[56];
  assign t[142] = t[186] ^ x[60];
  assign t[143] = t[187] ^ x[59];
  assign t[144] = t[188] ^ x[63];
  assign t[145] = t[189] ^ x[62];
  assign t[146] = t[190] ^ x[66];
  assign t[147] = t[191] ^ x[65];
  assign t[148] = (x[0]);
  assign t[149] = (x[0]);
  assign t[14] = t[18] ? t[39] : t[19];
  assign t[150] = (x[3]);
  assign t[151] = (x[3]);
  assign t[152] = (x[7]);
  assign t[153] = (x[7]);
  assign t[154] = (x[10]);
  assign t[155] = (x[10]);
  assign t[156] = (x[13]);
  assign t[157] = (x[13]);
  assign t[158] = (x[16]);
  assign t[159] = (x[16]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[19]);
  assign t[161] = (x[19]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[25]);
  assign t[165] = (x[25]);
  assign t[166] = (x[28]);
  assign t[167] = (x[28]);
  assign t[168] = (x[31]);
  assign t[169] = (x[31]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[34]);
  assign t[171] = (x[34]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[40]);
  assign t[175] = (x[40]);
  assign t[176] = (x[43]);
  assign t[177] = (x[43]);
  assign t[178] = (x[46]);
  assign t[179] = (x[46]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[49]);
  assign t[181] = (x[49]);
  assign t[182] = (x[52]);
  assign t[183] = (x[52]);
  assign t[184] = (x[55]);
  assign t[185] = (x[55]);
  assign t[186] = (x[58]);
  assign t[187] = (x[58]);
  assign t[188] = (x[61]);
  assign t[189] = (x[61]);
  assign t[18] = ~(t[25]);
  assign t[190] = (x[64]);
  assign t[191] = (x[64]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[43] | t[44]);
  assign t[23] = ~(t[45] | t[46]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[34] ^ t[35];
  assign t[27] = ~(t[47] ^ t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[53] & t[36]);
  assign t[32] = ~(t[54]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[55] ^ t[56];
  assign t[35] = t[41] ^ t[37];
  assign t[36] = ~(t[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[38] = (t[60]);
  assign t[39] = (t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[82] ^ x[2];
  assign t[61] = t[83] ^ x[5];
  assign t[62] = t[84] ^ x[9];
  assign t[63] = t[85] ^ x[12];
  assign t[64] = t[86] ^ x[15];
  assign t[65] = t[87] ^ x[18];
  assign t[66] = t[88] ^ x[21];
  assign t[67] = t[89] ^ x[24];
  assign t[68] = t[90] ^ x[27];
  assign t[69] = t[91] ^ x[30];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[33];
  assign t[71] = t[93] ^ x[36];
  assign t[72] = t[94] ^ x[39];
  assign t[73] = t[95] ^ x[42];
  assign t[74] = t[96] ^ x[45];
  assign t[75] = t[97] ^ x[48];
  assign t[76] = t[98] ^ x[51];
  assign t[77] = t[99] ^ x[54];
  assign t[78] = t[100] ^ x[57];
  assign t[79] = t[101] ^ x[60];
  assign t[7] = ~(t[40] & t[11]);
  assign t[80] = t[102] ^ x[63];
  assign t[81] = t[103] ^ x[66];
  assign t[82] = (t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[107]);
  assign t[84] = (t[108] & ~t[109]);
  assign t[85] = (t[110] & ~t[111]);
  assign t[86] = (t[112] & ~t[113]);
  assign t[87] = (t[114] & ~t[115]);
  assign t[88] = (t[116] & ~t[117]);
  assign t[89] = (t[118] & ~t[119]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[120] & ~t[121]);
  assign t[91] = (t[122] & ~t[123]);
  assign t[92] = (t[124] & ~t[125]);
  assign t[93] = (t[126] & ~t[127]);
  assign t[94] = (t[128] & ~t[129]);
  assign t[95] = (t[130] & ~t[131]);
  assign t[96] = (t[132] & ~t[133]);
  assign t[97] = (t[134] & ~t[135]);
  assign t[98] = (t[136] & ~t[137]);
  assign t[99] = (t[138] & ~t[139]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind412(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind413(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind414(x, y);
 input [66:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[140] & ~t[141]);
  assign t[101] = (t[142] & ~t[143]);
  assign t[102] = (t[144] & ~t[145]);
  assign t[103] = (t[146] & ~t[147]);
  assign t[104] = t[148] ^ x[2];
  assign t[105] = t[149] ^ x[1];
  assign t[106] = t[150] ^ x[5];
  assign t[107] = t[151] ^ x[4];
  assign t[108] = t[152] ^ x[9];
  assign t[109] = t[153] ^ x[8];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[154] ^ x[12];
  assign t[111] = t[155] ^ x[11];
  assign t[112] = t[156] ^ x[15];
  assign t[113] = t[157] ^ x[14];
  assign t[114] = t[158] ^ x[18];
  assign t[115] = t[159] ^ x[17];
  assign t[116] = t[160] ^ x[21];
  assign t[117] = t[161] ^ x[20];
  assign t[118] = t[162] ^ x[24];
  assign t[119] = t[163] ^ x[23];
  assign t[11] = ~(t[42] | t[16]);
  assign t[120] = t[164] ^ x[27];
  assign t[121] = t[165] ^ x[26];
  assign t[122] = t[166] ^ x[30];
  assign t[123] = t[167] ^ x[29];
  assign t[124] = t[168] ^ x[33];
  assign t[125] = t[169] ^ x[32];
  assign t[126] = t[170] ^ x[36];
  assign t[127] = t[171] ^ x[35];
  assign t[128] = t[172] ^ x[39];
  assign t[129] = t[173] ^ x[38];
  assign t[12] = ~(t[40]);
  assign t[130] = t[174] ^ x[42];
  assign t[131] = t[175] ^ x[41];
  assign t[132] = t[176] ^ x[45];
  assign t[133] = t[177] ^ x[44];
  assign t[134] = t[178] ^ x[48];
  assign t[135] = t[179] ^ x[47];
  assign t[136] = t[180] ^ x[51];
  assign t[137] = t[181] ^ x[50];
  assign t[138] = t[182] ^ x[54];
  assign t[139] = t[183] ^ x[53];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[57];
  assign t[141] = t[185] ^ x[56];
  assign t[142] = t[186] ^ x[60];
  assign t[143] = t[187] ^ x[59];
  assign t[144] = t[188] ^ x[63];
  assign t[145] = t[189] ^ x[62];
  assign t[146] = t[190] ^ x[66];
  assign t[147] = t[191] ^ x[65];
  assign t[148] = (x[0]);
  assign t[149] = (x[0]);
  assign t[14] = t[18] ? t[39] : t[19];
  assign t[150] = (x[3]);
  assign t[151] = (x[3]);
  assign t[152] = (x[7]);
  assign t[153] = (x[7]);
  assign t[154] = (x[10]);
  assign t[155] = (x[10]);
  assign t[156] = (x[13]);
  assign t[157] = (x[13]);
  assign t[158] = (x[16]);
  assign t[159] = (x[16]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[19]);
  assign t[161] = (x[19]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[25]);
  assign t[165] = (x[25]);
  assign t[166] = (x[28]);
  assign t[167] = (x[28]);
  assign t[168] = (x[31]);
  assign t[169] = (x[31]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[34]);
  assign t[171] = (x[34]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[40]);
  assign t[175] = (x[40]);
  assign t[176] = (x[43]);
  assign t[177] = (x[43]);
  assign t[178] = (x[46]);
  assign t[179] = (x[46]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[49]);
  assign t[181] = (x[49]);
  assign t[182] = (x[52]);
  assign t[183] = (x[52]);
  assign t[184] = (x[55]);
  assign t[185] = (x[55]);
  assign t[186] = (x[58]);
  assign t[187] = (x[58]);
  assign t[188] = (x[61]);
  assign t[189] = (x[61]);
  assign t[18] = ~(t[25]);
  assign t[190] = (x[64]);
  assign t[191] = (x[64]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[43] | t[44]);
  assign t[23] = ~(t[45] | t[46]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[34] ^ t[35];
  assign t[27] = ~(t[47] ^ t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[53] & t[36]);
  assign t[32] = ~(t[54]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[55] ^ t[56];
  assign t[35] = t[41] ^ t[37];
  assign t[36] = ~(t[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[38] = (t[60]);
  assign t[39] = (t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[82] ^ x[2];
  assign t[61] = t[83] ^ x[5];
  assign t[62] = t[84] ^ x[9];
  assign t[63] = t[85] ^ x[12];
  assign t[64] = t[86] ^ x[15];
  assign t[65] = t[87] ^ x[18];
  assign t[66] = t[88] ^ x[21];
  assign t[67] = t[89] ^ x[24];
  assign t[68] = t[90] ^ x[27];
  assign t[69] = t[91] ^ x[30];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[33];
  assign t[71] = t[93] ^ x[36];
  assign t[72] = t[94] ^ x[39];
  assign t[73] = t[95] ^ x[42];
  assign t[74] = t[96] ^ x[45];
  assign t[75] = t[97] ^ x[48];
  assign t[76] = t[98] ^ x[51];
  assign t[77] = t[99] ^ x[54];
  assign t[78] = t[100] ^ x[57];
  assign t[79] = t[101] ^ x[60];
  assign t[7] = ~(t[40] & t[11]);
  assign t[80] = t[102] ^ x[63];
  assign t[81] = t[103] ^ x[66];
  assign t[82] = (t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[107]);
  assign t[84] = (t[108] & ~t[109]);
  assign t[85] = (t[110] & ~t[111]);
  assign t[86] = (t[112] & ~t[113]);
  assign t[87] = (t[114] & ~t[115]);
  assign t[88] = (t[116] & ~t[117]);
  assign t[89] = (t[118] & ~t[119]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[120] & ~t[121]);
  assign t[91] = (t[122] & ~t[123]);
  assign t[92] = (t[124] & ~t[125]);
  assign t[93] = (t[126] & ~t[127]);
  assign t[94] = (t[128] & ~t[129]);
  assign t[95] = (t[130] & ~t[131]);
  assign t[96] = (t[132] & ~t[133]);
  assign t[97] = (t[134] & ~t[135]);
  assign t[98] = (t[136] & ~t[137]);
  assign t[99] = (t[138] & ~t[139]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind415(x, y);
 input [66:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[140] & ~t[141]);
  assign t[101] = (t[142] & ~t[143]);
  assign t[102] = (t[144] & ~t[145]);
  assign t[103] = (t[146] & ~t[147]);
  assign t[104] = t[148] ^ x[2];
  assign t[105] = t[149] ^ x[1];
  assign t[106] = t[150] ^ x[5];
  assign t[107] = t[151] ^ x[4];
  assign t[108] = t[152] ^ x[9];
  assign t[109] = t[153] ^ x[8];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[154] ^ x[12];
  assign t[111] = t[155] ^ x[11];
  assign t[112] = t[156] ^ x[15];
  assign t[113] = t[157] ^ x[14];
  assign t[114] = t[158] ^ x[18];
  assign t[115] = t[159] ^ x[17];
  assign t[116] = t[160] ^ x[21];
  assign t[117] = t[161] ^ x[20];
  assign t[118] = t[162] ^ x[24];
  assign t[119] = t[163] ^ x[23];
  assign t[11] = ~(t[42] | t[16]);
  assign t[120] = t[164] ^ x[27];
  assign t[121] = t[165] ^ x[26];
  assign t[122] = t[166] ^ x[30];
  assign t[123] = t[167] ^ x[29];
  assign t[124] = t[168] ^ x[33];
  assign t[125] = t[169] ^ x[32];
  assign t[126] = t[170] ^ x[36];
  assign t[127] = t[171] ^ x[35];
  assign t[128] = t[172] ^ x[39];
  assign t[129] = t[173] ^ x[38];
  assign t[12] = ~(t[40]);
  assign t[130] = t[174] ^ x[42];
  assign t[131] = t[175] ^ x[41];
  assign t[132] = t[176] ^ x[45];
  assign t[133] = t[177] ^ x[44];
  assign t[134] = t[178] ^ x[48];
  assign t[135] = t[179] ^ x[47];
  assign t[136] = t[180] ^ x[51];
  assign t[137] = t[181] ^ x[50];
  assign t[138] = t[182] ^ x[54];
  assign t[139] = t[183] ^ x[53];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[57];
  assign t[141] = t[185] ^ x[56];
  assign t[142] = t[186] ^ x[60];
  assign t[143] = t[187] ^ x[59];
  assign t[144] = t[188] ^ x[63];
  assign t[145] = t[189] ^ x[62];
  assign t[146] = t[190] ^ x[66];
  assign t[147] = t[191] ^ x[65];
  assign t[148] = (x[0]);
  assign t[149] = (x[0]);
  assign t[14] = t[18] ? t[39] : t[19];
  assign t[150] = (x[3]);
  assign t[151] = (x[3]);
  assign t[152] = (x[7]);
  assign t[153] = (x[7]);
  assign t[154] = (x[10]);
  assign t[155] = (x[10]);
  assign t[156] = (x[13]);
  assign t[157] = (x[13]);
  assign t[158] = (x[16]);
  assign t[159] = (x[16]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[19]);
  assign t[161] = (x[19]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[25]);
  assign t[165] = (x[25]);
  assign t[166] = (x[28]);
  assign t[167] = (x[28]);
  assign t[168] = (x[31]);
  assign t[169] = (x[31]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[34]);
  assign t[171] = (x[34]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[40]);
  assign t[175] = (x[40]);
  assign t[176] = (x[43]);
  assign t[177] = (x[43]);
  assign t[178] = (x[46]);
  assign t[179] = (x[46]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[49]);
  assign t[181] = (x[49]);
  assign t[182] = (x[52]);
  assign t[183] = (x[52]);
  assign t[184] = (x[55]);
  assign t[185] = (x[55]);
  assign t[186] = (x[58]);
  assign t[187] = (x[58]);
  assign t[188] = (x[61]);
  assign t[189] = (x[61]);
  assign t[18] = ~(t[25]);
  assign t[190] = (x[64]);
  assign t[191] = (x[64]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[43] | t[44]);
  assign t[23] = ~(t[45] | t[46]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[34] ^ t[35];
  assign t[27] = ~(t[47] ^ t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[53] & t[36]);
  assign t[32] = ~(t[54]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[55] ^ t[56];
  assign t[35] = t[41] ^ t[37];
  assign t[36] = ~(t[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[38] = (t[60]);
  assign t[39] = (t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[82] ^ x[2];
  assign t[61] = t[83] ^ x[5];
  assign t[62] = t[84] ^ x[9];
  assign t[63] = t[85] ^ x[12];
  assign t[64] = t[86] ^ x[15];
  assign t[65] = t[87] ^ x[18];
  assign t[66] = t[88] ^ x[21];
  assign t[67] = t[89] ^ x[24];
  assign t[68] = t[90] ^ x[27];
  assign t[69] = t[91] ^ x[30];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[33];
  assign t[71] = t[93] ^ x[36];
  assign t[72] = t[94] ^ x[39];
  assign t[73] = t[95] ^ x[42];
  assign t[74] = t[96] ^ x[45];
  assign t[75] = t[97] ^ x[48];
  assign t[76] = t[98] ^ x[51];
  assign t[77] = t[99] ^ x[54];
  assign t[78] = t[100] ^ x[57];
  assign t[79] = t[101] ^ x[60];
  assign t[7] = ~(t[40] & t[11]);
  assign t[80] = t[102] ^ x[63];
  assign t[81] = t[103] ^ x[66];
  assign t[82] = (t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[107]);
  assign t[84] = (t[108] & ~t[109]);
  assign t[85] = (t[110] & ~t[111]);
  assign t[86] = (t[112] & ~t[113]);
  assign t[87] = (t[114] & ~t[115]);
  assign t[88] = (t[116] & ~t[117]);
  assign t[89] = (t[118] & ~t[119]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[120] & ~t[121]);
  assign t[91] = (t[122] & ~t[123]);
  assign t[92] = (t[124] & ~t[125]);
  assign t[93] = (t[126] & ~t[127]);
  assign t[94] = (t[128] & ~t[129]);
  assign t[95] = (t[130] & ~t[131]);
  assign t[96] = (t[132] & ~t[133]);
  assign t[97] = (t[134] & ~t[135]);
  assign t[98] = (t[136] & ~t[137]);
  assign t[99] = (t[138] & ~t[139]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind416(x, y);
 input [66:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[140] & ~t[141]);
  assign t[101] = (t[142] & ~t[143]);
  assign t[102] = (t[144] & ~t[145]);
  assign t[103] = (t[146] & ~t[147]);
  assign t[104] = t[148] ^ x[2];
  assign t[105] = t[149] ^ x[1];
  assign t[106] = t[150] ^ x[5];
  assign t[107] = t[151] ^ x[4];
  assign t[108] = t[152] ^ x[9];
  assign t[109] = t[153] ^ x[8];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[154] ^ x[12];
  assign t[111] = t[155] ^ x[11];
  assign t[112] = t[156] ^ x[15];
  assign t[113] = t[157] ^ x[14];
  assign t[114] = t[158] ^ x[18];
  assign t[115] = t[159] ^ x[17];
  assign t[116] = t[160] ^ x[21];
  assign t[117] = t[161] ^ x[20];
  assign t[118] = t[162] ^ x[24];
  assign t[119] = t[163] ^ x[23];
  assign t[11] = ~(t[42] | t[16]);
  assign t[120] = t[164] ^ x[27];
  assign t[121] = t[165] ^ x[26];
  assign t[122] = t[166] ^ x[30];
  assign t[123] = t[167] ^ x[29];
  assign t[124] = t[168] ^ x[33];
  assign t[125] = t[169] ^ x[32];
  assign t[126] = t[170] ^ x[36];
  assign t[127] = t[171] ^ x[35];
  assign t[128] = t[172] ^ x[39];
  assign t[129] = t[173] ^ x[38];
  assign t[12] = ~(t[40]);
  assign t[130] = t[174] ^ x[42];
  assign t[131] = t[175] ^ x[41];
  assign t[132] = t[176] ^ x[45];
  assign t[133] = t[177] ^ x[44];
  assign t[134] = t[178] ^ x[48];
  assign t[135] = t[179] ^ x[47];
  assign t[136] = t[180] ^ x[51];
  assign t[137] = t[181] ^ x[50];
  assign t[138] = t[182] ^ x[54];
  assign t[139] = t[183] ^ x[53];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[57];
  assign t[141] = t[185] ^ x[56];
  assign t[142] = t[186] ^ x[60];
  assign t[143] = t[187] ^ x[59];
  assign t[144] = t[188] ^ x[63];
  assign t[145] = t[189] ^ x[62];
  assign t[146] = t[190] ^ x[66];
  assign t[147] = t[191] ^ x[65];
  assign t[148] = (x[0]);
  assign t[149] = (x[0]);
  assign t[14] = t[18] ? t[39] : t[19];
  assign t[150] = (x[3]);
  assign t[151] = (x[3]);
  assign t[152] = (x[7]);
  assign t[153] = (x[7]);
  assign t[154] = (x[10]);
  assign t[155] = (x[10]);
  assign t[156] = (x[13]);
  assign t[157] = (x[13]);
  assign t[158] = (x[16]);
  assign t[159] = (x[16]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[19]);
  assign t[161] = (x[19]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[25]);
  assign t[165] = (x[25]);
  assign t[166] = (x[28]);
  assign t[167] = (x[28]);
  assign t[168] = (x[31]);
  assign t[169] = (x[31]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[34]);
  assign t[171] = (x[34]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[40]);
  assign t[175] = (x[40]);
  assign t[176] = (x[43]);
  assign t[177] = (x[43]);
  assign t[178] = (x[46]);
  assign t[179] = (x[46]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[49]);
  assign t[181] = (x[49]);
  assign t[182] = (x[52]);
  assign t[183] = (x[52]);
  assign t[184] = (x[55]);
  assign t[185] = (x[55]);
  assign t[186] = (x[58]);
  assign t[187] = (x[58]);
  assign t[188] = (x[61]);
  assign t[189] = (x[61]);
  assign t[18] = ~(t[25]);
  assign t[190] = (x[64]);
  assign t[191] = (x[64]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[43] | t[44]);
  assign t[23] = ~(t[45] | t[46]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[34] ^ t[35];
  assign t[27] = ~(t[47] ^ t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[53] & t[36]);
  assign t[32] = ~(t[54]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[55] ^ t[56];
  assign t[35] = t[41] ^ t[37];
  assign t[36] = ~(t[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[38] = (t[60]);
  assign t[39] = (t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[82] ^ x[2];
  assign t[61] = t[83] ^ x[5];
  assign t[62] = t[84] ^ x[9];
  assign t[63] = t[85] ^ x[12];
  assign t[64] = t[86] ^ x[15];
  assign t[65] = t[87] ^ x[18];
  assign t[66] = t[88] ^ x[21];
  assign t[67] = t[89] ^ x[24];
  assign t[68] = t[90] ^ x[27];
  assign t[69] = t[91] ^ x[30];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[33];
  assign t[71] = t[93] ^ x[36];
  assign t[72] = t[94] ^ x[39];
  assign t[73] = t[95] ^ x[42];
  assign t[74] = t[96] ^ x[45];
  assign t[75] = t[97] ^ x[48];
  assign t[76] = t[98] ^ x[51];
  assign t[77] = t[99] ^ x[54];
  assign t[78] = t[100] ^ x[57];
  assign t[79] = t[101] ^ x[60];
  assign t[7] = ~(t[40] & t[11]);
  assign t[80] = t[102] ^ x[63];
  assign t[81] = t[103] ^ x[66];
  assign t[82] = (t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[107]);
  assign t[84] = (t[108] & ~t[109]);
  assign t[85] = (t[110] & ~t[111]);
  assign t[86] = (t[112] & ~t[113]);
  assign t[87] = (t[114] & ~t[115]);
  assign t[88] = (t[116] & ~t[117]);
  assign t[89] = (t[118] & ~t[119]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[120] & ~t[121]);
  assign t[91] = (t[122] & ~t[123]);
  assign t[92] = (t[124] & ~t[125]);
  assign t[93] = (t[126] & ~t[127]);
  assign t[94] = (t[128] & ~t[129]);
  assign t[95] = (t[130] & ~t[131]);
  assign t[96] = (t[132] & ~t[133]);
  assign t[97] = (t[134] & ~t[135]);
  assign t[98] = (t[136] & ~t[137]);
  assign t[99] = (t[138] & ~t[139]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind417(x, y);
 input [66:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[140] & ~t[141]);
  assign t[101] = (t[142] & ~t[143]);
  assign t[102] = (t[144] & ~t[145]);
  assign t[103] = (t[146] & ~t[147]);
  assign t[104] = t[148] ^ x[2];
  assign t[105] = t[149] ^ x[1];
  assign t[106] = t[150] ^ x[5];
  assign t[107] = t[151] ^ x[4];
  assign t[108] = t[152] ^ x[9];
  assign t[109] = t[153] ^ x[8];
  assign t[10] = t[40] & t[15];
  assign t[110] = t[154] ^ x[12];
  assign t[111] = t[155] ^ x[11];
  assign t[112] = t[156] ^ x[15];
  assign t[113] = t[157] ^ x[14];
  assign t[114] = t[158] ^ x[18];
  assign t[115] = t[159] ^ x[17];
  assign t[116] = t[160] ^ x[21];
  assign t[117] = t[161] ^ x[20];
  assign t[118] = t[162] ^ x[24];
  assign t[119] = t[163] ^ x[23];
  assign t[11] = ~(t[42] | t[16]);
  assign t[120] = t[164] ^ x[27];
  assign t[121] = t[165] ^ x[26];
  assign t[122] = t[166] ^ x[30];
  assign t[123] = t[167] ^ x[29];
  assign t[124] = t[168] ^ x[33];
  assign t[125] = t[169] ^ x[32];
  assign t[126] = t[170] ^ x[36];
  assign t[127] = t[171] ^ x[35];
  assign t[128] = t[172] ^ x[39];
  assign t[129] = t[173] ^ x[38];
  assign t[12] = ~(t[40]);
  assign t[130] = t[174] ^ x[42];
  assign t[131] = t[175] ^ x[41];
  assign t[132] = t[176] ^ x[45];
  assign t[133] = t[177] ^ x[44];
  assign t[134] = t[178] ^ x[48];
  assign t[135] = t[179] ^ x[47];
  assign t[136] = t[180] ^ x[51];
  assign t[137] = t[181] ^ x[50];
  assign t[138] = t[182] ^ x[54];
  assign t[139] = t[183] ^ x[53];
  assign t[13] = ~(t[17]);
  assign t[140] = t[184] ^ x[57];
  assign t[141] = t[185] ^ x[56];
  assign t[142] = t[186] ^ x[60];
  assign t[143] = t[187] ^ x[59];
  assign t[144] = t[188] ^ x[63];
  assign t[145] = t[189] ^ x[62];
  assign t[146] = t[190] ^ x[66];
  assign t[147] = t[191] ^ x[65];
  assign t[148] = (x[0]);
  assign t[149] = (x[0]);
  assign t[14] = t[18] ? t[39] : t[19];
  assign t[150] = (x[3]);
  assign t[151] = (x[3]);
  assign t[152] = (x[7]);
  assign t[153] = (x[7]);
  assign t[154] = (x[10]);
  assign t[155] = (x[10]);
  assign t[156] = (x[13]);
  assign t[157] = (x[13]);
  assign t[158] = (x[16]);
  assign t[159] = (x[16]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[19]);
  assign t[161] = (x[19]);
  assign t[162] = (x[22]);
  assign t[163] = (x[22]);
  assign t[164] = (x[25]);
  assign t[165] = (x[25]);
  assign t[166] = (x[28]);
  assign t[167] = (x[28]);
  assign t[168] = (x[31]);
  assign t[169] = (x[31]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[34]);
  assign t[171] = (x[34]);
  assign t[172] = (x[37]);
  assign t[173] = (x[37]);
  assign t[174] = (x[40]);
  assign t[175] = (x[40]);
  assign t[176] = (x[43]);
  assign t[177] = (x[43]);
  assign t[178] = (x[46]);
  assign t[179] = (x[46]);
  assign t[17] = ~(t[24]);
  assign t[180] = (x[49]);
  assign t[181] = (x[49]);
  assign t[182] = (x[52]);
  assign t[183] = (x[52]);
  assign t[184] = (x[55]);
  assign t[185] = (x[55]);
  assign t[186] = (x[58]);
  assign t[187] = (x[58]);
  assign t[188] = (x[61]);
  assign t[189] = (x[61]);
  assign t[18] = ~(t[25]);
  assign t[190] = (x[64]);
  assign t[191] = (x[64]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[43] | t[44]);
  assign t[23] = ~(t[45] | t[46]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[34] ^ t[35];
  assign t[27] = ~(t[47] ^ t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[51] & t[52]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[53] & t[36]);
  assign t[32] = ~(t[54]);
  assign t[33] = ~(t[40]);
  assign t[34] = t[55] ^ t[56];
  assign t[35] = t[41] ^ t[37];
  assign t[36] = ~(t[57]);
  assign t[37] = t[58] ^ t[59];
  assign t[38] = (t[60]);
  assign t[39] = (t[61]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[62]);
  assign t[41] = (t[63]);
  assign t[42] = (t[64]);
  assign t[43] = (t[65]);
  assign t[44] = (t[66]);
  assign t[45] = (t[67]);
  assign t[46] = (t[68]);
  assign t[47] = (t[69]);
  assign t[48] = (t[70]);
  assign t[49] = (t[71]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[72]);
  assign t[51] = (t[73]);
  assign t[52] = (t[74]);
  assign t[53] = (t[75]);
  assign t[54] = (t[76]);
  assign t[55] = (t[77]);
  assign t[56] = (t[78]);
  assign t[57] = (t[79]);
  assign t[58] = (t[80]);
  assign t[59] = (t[81]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[82] ^ x[2];
  assign t[61] = t[83] ^ x[5];
  assign t[62] = t[84] ^ x[9];
  assign t[63] = t[85] ^ x[12];
  assign t[64] = t[86] ^ x[15];
  assign t[65] = t[87] ^ x[18];
  assign t[66] = t[88] ^ x[21];
  assign t[67] = t[89] ^ x[24];
  assign t[68] = t[90] ^ x[27];
  assign t[69] = t[91] ^ x[30];
  assign t[6] = ~(t[10]);
  assign t[70] = t[92] ^ x[33];
  assign t[71] = t[93] ^ x[36];
  assign t[72] = t[94] ^ x[39];
  assign t[73] = t[95] ^ x[42];
  assign t[74] = t[96] ^ x[45];
  assign t[75] = t[97] ^ x[48];
  assign t[76] = t[98] ^ x[51];
  assign t[77] = t[99] ^ x[54];
  assign t[78] = t[100] ^ x[57];
  assign t[79] = t[101] ^ x[60];
  assign t[7] = ~(t[40] & t[11]);
  assign t[80] = t[102] ^ x[63];
  assign t[81] = t[103] ^ x[66];
  assign t[82] = (t[104] & ~t[105]);
  assign t[83] = (t[106] & ~t[107]);
  assign t[84] = (t[108] & ~t[109]);
  assign t[85] = (t[110] & ~t[111]);
  assign t[86] = (t[112] & ~t[113]);
  assign t[87] = (t[114] & ~t[115]);
  assign t[88] = (t[116] & ~t[117]);
  assign t[89] = (t[118] & ~t[119]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[120] & ~t[121]);
  assign t[91] = (t[122] & ~t[123]);
  assign t[92] = (t[124] & ~t[125]);
  assign t[93] = (t[126] & ~t[127]);
  assign t[94] = (t[128] & ~t[129]);
  assign t[95] = (t[130] & ~t[131]);
  assign t[96] = (t[132] & ~t[133]);
  assign t[97] = (t[134] & ~t[135]);
  assign t[98] = (t[136] & ~t[137]);
  assign t[99] = (t[138] & ~t[139]);
  assign t[9] = t[13] ? t[14] : t[41];
  assign y = (t[0]);
endmodule

module R2ind418(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind419(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind420(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind421(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind422(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind423(x, y);
 input [60:0] x;
 output y;

 wire [175:0] t;
  assign t[0] = t[1] ? t[2] : t[36];
  assign t[100] = t[140] ^ x[9];
  assign t[101] = t[141] ^ x[8];
  assign t[102] = t[142] ^ x[12];
  assign t[103] = t[143] ^ x[11];
  assign t[104] = t[144] ^ x[15];
  assign t[105] = t[145] ^ x[14];
  assign t[106] = t[146] ^ x[18];
  assign t[107] = t[147] ^ x[17];
  assign t[108] = t[148] ^ x[21];
  assign t[109] = t[149] ^ x[20];
  assign t[10] = t[38] & t[15];
  assign t[110] = t[150] ^ x[24];
  assign t[111] = t[151] ^ x[23];
  assign t[112] = t[152] ^ x[27];
  assign t[113] = t[153] ^ x[26];
  assign t[114] = t[154] ^ x[30];
  assign t[115] = t[155] ^ x[29];
  assign t[116] = t[156] ^ x[33];
  assign t[117] = t[157] ^ x[32];
  assign t[118] = t[158] ^ x[36];
  assign t[119] = t[159] ^ x[35];
  assign t[11] = ~(t[40] | t[16]);
  assign t[120] = t[160] ^ x[39];
  assign t[121] = t[161] ^ x[38];
  assign t[122] = t[162] ^ x[42];
  assign t[123] = t[163] ^ x[41];
  assign t[124] = t[164] ^ x[45];
  assign t[125] = t[165] ^ x[44];
  assign t[126] = t[166] ^ x[48];
  assign t[127] = t[167] ^ x[47];
  assign t[128] = t[168] ^ x[51];
  assign t[129] = t[169] ^ x[50];
  assign t[12] = ~(t[38]);
  assign t[130] = t[170] ^ x[54];
  assign t[131] = t[171] ^ x[53];
  assign t[132] = t[172] ^ x[57];
  assign t[133] = t[173] ^ x[56];
  assign t[134] = t[174] ^ x[60];
  assign t[135] = t[175] ^ x[59];
  assign t[136] = (x[0]);
  assign t[137] = (x[0]);
  assign t[138] = (x[3]);
  assign t[139] = (x[3]);
  assign t[13] = ~(t[17]);
  assign t[140] = (x[7]);
  assign t[141] = (x[7]);
  assign t[142] = (x[10]);
  assign t[143] = (x[10]);
  assign t[144] = (x[13]);
  assign t[145] = (x[13]);
  assign t[146] = (x[16]);
  assign t[147] = (x[16]);
  assign t[148] = (x[19]);
  assign t[149] = (x[19]);
  assign t[14] = t[18] ? t[37] : t[19];
  assign t[150] = (x[22]);
  assign t[151] = (x[22]);
  assign t[152] = (x[25]);
  assign t[153] = (x[25]);
  assign t[154] = (x[28]);
  assign t[155] = (x[28]);
  assign t[156] = (x[31]);
  assign t[157] = (x[31]);
  assign t[158] = (x[34]);
  assign t[159] = (x[34]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[37]);
  assign t[161] = (x[37]);
  assign t[162] = (x[40]);
  assign t[163] = (x[40]);
  assign t[164] = (x[43]);
  assign t[165] = (x[43]);
  assign t[166] = (x[46]);
  assign t[167] = (x[46]);
  assign t[168] = (x[49]);
  assign t[169] = (x[49]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[170] = (x[52]);
  assign t[171] = (x[52]);
  assign t[172] = (x[55]);
  assign t[173] = (x[55]);
  assign t[174] = (x[58]);
  assign t[175] = (x[58]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[25]);
  assign t[19] = ~(t[26] ^ t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[28] | t[29]);
  assign t[21] = ~(t[30] | t[31]);
  assign t[22] = ~(t[41] | t[42]);
  assign t[23] = ~(t[43] | t[44]);
  assign t[24] = ~(t[32] | t[33]);
  assign t[25] = ~(t[20]);
  assign t[26] = t[45] ^ t[34];
  assign t[27] = ~(t[46] ^ t[47]);
  assign t[28] = ~(t[48] & t[49]);
  assign t[29] = ~(t[50] & t[51]);
  assign t[2] = t[4] ? t[37] : t[5];
  assign t[30] = ~(t[11]);
  assign t[31] = ~(t[52] & t[35]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ t[54];
  assign t[35] = ~(t[55]);
  assign t[36] = (t[56]);
  assign t[37] = (t[57]);
  assign t[38] = (t[58]);
  assign t[39] = (t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[60]);
  assign t[41] = (t[61]);
  assign t[42] = (t[62]);
  assign t[43] = (t[63]);
  assign t[44] = (t[64]);
  assign t[45] = (t[65]);
  assign t[46] = (t[66]);
  assign t[47] = (t[67]);
  assign t[48] = (t[68]);
  assign t[49] = (t[69]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[70]);
  assign t[51] = (t[71]);
  assign t[52] = (t[72]);
  assign t[53] = (t[73]);
  assign t[54] = (t[74]);
  assign t[55] = (t[75]);
  assign t[56] = t[76] ^ x[2];
  assign t[57] = t[77] ^ x[5];
  assign t[58] = t[78] ^ x[9];
  assign t[59] = t[79] ^ x[12];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[80] ^ x[15];
  assign t[61] = t[81] ^ x[18];
  assign t[62] = t[82] ^ x[21];
  assign t[63] = t[83] ^ x[24];
  assign t[64] = t[84] ^ x[27];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = t[86] ^ x[33];
  assign t[67] = t[87] ^ x[36];
  assign t[68] = t[88] ^ x[39];
  assign t[69] = t[89] ^ x[42];
  assign t[6] = ~(t[10]);
  assign t[70] = t[90] ^ x[45];
  assign t[71] = t[91] ^ x[48];
  assign t[72] = t[92] ^ x[51];
  assign t[73] = t[93] ^ x[54];
  assign t[74] = t[94] ^ x[57];
  assign t[75] = t[95] ^ x[60];
  assign t[76] = (t[96] & ~t[97]);
  assign t[77] = (t[98] & ~t[99]);
  assign t[78] = (t[100] & ~t[101]);
  assign t[79] = (t[102] & ~t[103]);
  assign t[7] = ~(t[38] & t[11]);
  assign t[80] = (t[104] & ~t[105]);
  assign t[81] = (t[106] & ~t[107]);
  assign t[82] = (t[108] & ~t[109]);
  assign t[83] = (t[110] & ~t[111]);
  assign t[84] = (t[112] & ~t[113]);
  assign t[85] = (t[114] & ~t[115]);
  assign t[86] = (t[116] & ~t[117]);
  assign t[87] = (t[118] & ~t[119]);
  assign t[88] = (t[120] & ~t[121]);
  assign t[89] = (t[122] & ~t[123]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[124] & ~t[125]);
  assign t[91] = (t[126] & ~t[127]);
  assign t[92] = (t[128] & ~t[129]);
  assign t[93] = (t[130] & ~t[131]);
  assign t[94] = (t[132] & ~t[133]);
  assign t[95] = (t[134] & ~t[135]);
  assign t[96] = t[136] ^ x[2];
  assign t[97] = t[137] ^ x[1];
  assign t[98] = t[138] ^ x[5];
  assign t[99] = t[139] ^ x[4];
  assign t[9] = t[13] ? t[14] : t[39];
  assign y = (t[0]);
endmodule

module R2ind424(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind425(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind426(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind427(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind428(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind429(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind430(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind431(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind432(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind433(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind434(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind435(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind436(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind437(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind438(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind439(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind440(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind441(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind442(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind443(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind444(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind445(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind446(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind447(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind448(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind449(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind450(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind451(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind452(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind453(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind454(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind455(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind456(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind457(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind458(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind459(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind460(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind461(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind462(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind463(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind464(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind465(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind466(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind467(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind468(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind469(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind470(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind471(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind472(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind473(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind474(x, y);
 input [69:0] x;
 output y;

 wire [200:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[137] & ~t[138]);
  assign t[101] = (t[139] & ~t[140]);
  assign t[102] = (t[141] & ~t[142]);
  assign t[103] = (t[143] & ~t[144]);
  assign t[104] = (t[145] & ~t[146]);
  assign t[105] = (t[147] & ~t[148]);
  assign t[106] = (t[149] & ~t[150]);
  assign t[107] = (t[151] & ~t[152]);
  assign t[108] = (t[153] & ~t[154]);
  assign t[109] = t[155] ^ x[2];
  assign t[10] = t[43] & t[15];
  assign t[110] = t[156] ^ x[1];
  assign t[111] = t[157] ^ x[5];
  assign t[112] = t[158] ^ x[4];
  assign t[113] = t[159] ^ x[9];
  assign t[114] = t[160] ^ x[8];
  assign t[115] = t[161] ^ x[12];
  assign t[116] = t[162] ^ x[11];
  assign t[117] = t[163] ^ x[15];
  assign t[118] = t[164] ^ x[14];
  assign t[119] = t[165] ^ x[18];
  assign t[11] = ~(t[16]);
  assign t[120] = t[166] ^ x[17];
  assign t[121] = t[167] ^ x[21];
  assign t[122] = t[168] ^ x[20];
  assign t[123] = t[169] ^ x[24];
  assign t[124] = t[170] ^ x[23];
  assign t[125] = t[171] ^ x[27];
  assign t[126] = t[172] ^ x[26];
  assign t[127] = t[173] ^ x[30];
  assign t[128] = t[174] ^ x[29];
  assign t[129] = t[175] ^ x[33];
  assign t[12] = ~(t[43]);
  assign t[130] = t[176] ^ x[32];
  assign t[131] = t[177] ^ x[36];
  assign t[132] = t[178] ^ x[35];
  assign t[133] = t[179] ^ x[39];
  assign t[134] = t[180] ^ x[38];
  assign t[135] = t[181] ^ x[42];
  assign t[136] = t[182] ^ x[41];
  assign t[137] = t[183] ^ x[45];
  assign t[138] = t[184] ^ x[44];
  assign t[139] = t[185] ^ x[48];
  assign t[13] = ~(t[17]);
  assign t[140] = t[186] ^ x[47];
  assign t[141] = t[187] ^ x[51];
  assign t[142] = t[188] ^ x[50];
  assign t[143] = t[189] ^ x[54];
  assign t[144] = t[190] ^ x[53];
  assign t[145] = t[191] ^ x[57];
  assign t[146] = t[192] ^ x[56];
  assign t[147] = t[193] ^ x[60];
  assign t[148] = t[194] ^ x[59];
  assign t[149] = t[195] ^ x[63];
  assign t[14] = t[18] ? t[44] : t[19];
  assign t[150] = t[196] ^ x[62];
  assign t[151] = t[197] ^ x[66];
  assign t[152] = t[198] ^ x[65];
  assign t[153] = t[199] ^ x[69];
  assign t[154] = t[200] ^ x[68];
  assign t[155] = (x[0]);
  assign t[156] = (x[0]);
  assign t[157] = (x[3]);
  assign t[158] = (x[3]);
  assign t[159] = (x[7]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[7]);
  assign t[161] = (x[10]);
  assign t[162] = (x[10]);
  assign t[163] = (x[13]);
  assign t[164] = (x[13]);
  assign t[165] = (x[16]);
  assign t[166] = (x[16]);
  assign t[167] = (x[19]);
  assign t[168] = (x[19]);
  assign t[169] = (x[22]);
  assign t[16] = ~(t[43] & t[22]);
  assign t[170] = (x[22]);
  assign t[171] = (x[25]);
  assign t[172] = (x[25]);
  assign t[173] = (x[28]);
  assign t[174] = (x[28]);
  assign t[175] = (x[31]);
  assign t[176] = (x[31]);
  assign t[177] = (x[34]);
  assign t[178] = (x[34]);
  assign t[179] = (x[37]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[37]);
  assign t[181] = (x[40]);
  assign t[182] = (x[40]);
  assign t[183] = (x[43]);
  assign t[184] = (x[43]);
  assign t[185] = (x[46]);
  assign t[186] = (x[46]);
  assign t[187] = (x[49]);
  assign t[188] = (x[49]);
  assign t[189] = (x[52]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[52]);
  assign t[191] = (x[55]);
  assign t[192] = (x[55]);
  assign t[193] = (x[58]);
  assign t[194] = (x[58]);
  assign t[195] = (x[61]);
  assign t[196] = (x[61]);
  assign t[197] = (x[64]);
  assign t[198] = (x[64]);
  assign t[199] = (x[67]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = (x[67]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[45] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[41] : t[5];
  assign t[30] = ~(t[52] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[43]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[42] ^ t[39];
  assign t[36] = ~(t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[63]);
  assign t[41] = (t[64]);
  assign t[42] = (t[65]);
  assign t[43] = (t[66]);
  assign t[44] = (t[67]);
  assign t[45] = (t[68]);
  assign t[46] = (t[69]);
  assign t[47] = (t[70]);
  assign t[48] = (t[71]);
  assign t[49] = (t[72]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[73]);
  assign t[51] = (t[74]);
  assign t[52] = (t[75]);
  assign t[53] = (t[76]);
  assign t[54] = (t[77]);
  assign t[55] = (t[78]);
  assign t[56] = (t[79]);
  assign t[57] = (t[80]);
  assign t[58] = (t[81]);
  assign t[59] = (t[82]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[83]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = t[86] ^ x[2];
  assign t[64] = t[87] ^ x[5];
  assign t[65] = t[88] ^ x[9];
  assign t[66] = t[89] ^ x[12];
  assign t[67] = t[90] ^ x[15];
  assign t[68] = t[91] ^ x[18];
  assign t[69] = t[92] ^ x[21];
  assign t[6] = ~(t[10]);
  assign t[70] = t[93] ^ x[24];
  assign t[71] = t[94] ^ x[27];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[33];
  assign t[74] = t[97] ^ x[36];
  assign t[75] = t[98] ^ x[39];
  assign t[76] = t[99] ^ x[42];
  assign t[77] = t[100] ^ x[45];
  assign t[78] = t[101] ^ x[48];
  assign t[79] = t[102] ^ x[51];
  assign t[7] = ~(t[11]);
  assign t[80] = t[103] ^ x[54];
  assign t[81] = t[104] ^ x[57];
  assign t[82] = t[105] ^ x[60];
  assign t[83] = t[106] ^ x[63];
  assign t[84] = t[107] ^ x[66];
  assign t[85] = t[108] ^ x[69];
  assign t[86] = (t[109] & ~t[110]);
  assign t[87] = (t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[114]);
  assign t[89] = (t[115] & ~t[116]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[117] & ~t[118]);
  assign t[91] = (t[119] & ~t[120]);
  assign t[92] = (t[121] & ~t[122]);
  assign t[93] = (t[123] & ~t[124]);
  assign t[94] = (t[125] & ~t[126]);
  assign t[95] = (t[127] & ~t[128]);
  assign t[96] = (t[129] & ~t[130]);
  assign t[97] = (t[131] & ~t[132]);
  assign t[98] = (t[133] & ~t[134]);
  assign t[99] = (t[135] & ~t[136]);
  assign t[9] = t[13] ? t[14] : t[42];
  assign y = (t[0]);
endmodule

module R2ind475(x, y);
 input [69:0] x;
 output y;

 wire [200:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[137] & ~t[138]);
  assign t[101] = (t[139] & ~t[140]);
  assign t[102] = (t[141] & ~t[142]);
  assign t[103] = (t[143] & ~t[144]);
  assign t[104] = (t[145] & ~t[146]);
  assign t[105] = (t[147] & ~t[148]);
  assign t[106] = (t[149] & ~t[150]);
  assign t[107] = (t[151] & ~t[152]);
  assign t[108] = (t[153] & ~t[154]);
  assign t[109] = t[155] ^ x[2];
  assign t[10] = t[43] & t[15];
  assign t[110] = t[156] ^ x[1];
  assign t[111] = t[157] ^ x[5];
  assign t[112] = t[158] ^ x[4];
  assign t[113] = t[159] ^ x[9];
  assign t[114] = t[160] ^ x[8];
  assign t[115] = t[161] ^ x[12];
  assign t[116] = t[162] ^ x[11];
  assign t[117] = t[163] ^ x[15];
  assign t[118] = t[164] ^ x[14];
  assign t[119] = t[165] ^ x[18];
  assign t[11] = ~(t[16]);
  assign t[120] = t[166] ^ x[17];
  assign t[121] = t[167] ^ x[21];
  assign t[122] = t[168] ^ x[20];
  assign t[123] = t[169] ^ x[24];
  assign t[124] = t[170] ^ x[23];
  assign t[125] = t[171] ^ x[27];
  assign t[126] = t[172] ^ x[26];
  assign t[127] = t[173] ^ x[30];
  assign t[128] = t[174] ^ x[29];
  assign t[129] = t[175] ^ x[33];
  assign t[12] = ~(t[43]);
  assign t[130] = t[176] ^ x[32];
  assign t[131] = t[177] ^ x[36];
  assign t[132] = t[178] ^ x[35];
  assign t[133] = t[179] ^ x[39];
  assign t[134] = t[180] ^ x[38];
  assign t[135] = t[181] ^ x[42];
  assign t[136] = t[182] ^ x[41];
  assign t[137] = t[183] ^ x[45];
  assign t[138] = t[184] ^ x[44];
  assign t[139] = t[185] ^ x[48];
  assign t[13] = ~(t[17]);
  assign t[140] = t[186] ^ x[47];
  assign t[141] = t[187] ^ x[51];
  assign t[142] = t[188] ^ x[50];
  assign t[143] = t[189] ^ x[54];
  assign t[144] = t[190] ^ x[53];
  assign t[145] = t[191] ^ x[57];
  assign t[146] = t[192] ^ x[56];
  assign t[147] = t[193] ^ x[60];
  assign t[148] = t[194] ^ x[59];
  assign t[149] = t[195] ^ x[63];
  assign t[14] = t[18] ? t[44] : t[19];
  assign t[150] = t[196] ^ x[62];
  assign t[151] = t[197] ^ x[66];
  assign t[152] = t[198] ^ x[65];
  assign t[153] = t[199] ^ x[69];
  assign t[154] = t[200] ^ x[68];
  assign t[155] = (x[0]);
  assign t[156] = (x[0]);
  assign t[157] = (x[3]);
  assign t[158] = (x[3]);
  assign t[159] = (x[7]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[7]);
  assign t[161] = (x[10]);
  assign t[162] = (x[10]);
  assign t[163] = (x[13]);
  assign t[164] = (x[13]);
  assign t[165] = (x[16]);
  assign t[166] = (x[16]);
  assign t[167] = (x[19]);
  assign t[168] = (x[19]);
  assign t[169] = (x[22]);
  assign t[16] = ~(t[43] & t[22]);
  assign t[170] = (x[22]);
  assign t[171] = (x[25]);
  assign t[172] = (x[25]);
  assign t[173] = (x[28]);
  assign t[174] = (x[28]);
  assign t[175] = (x[31]);
  assign t[176] = (x[31]);
  assign t[177] = (x[34]);
  assign t[178] = (x[34]);
  assign t[179] = (x[37]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[37]);
  assign t[181] = (x[40]);
  assign t[182] = (x[40]);
  assign t[183] = (x[43]);
  assign t[184] = (x[43]);
  assign t[185] = (x[46]);
  assign t[186] = (x[46]);
  assign t[187] = (x[49]);
  assign t[188] = (x[49]);
  assign t[189] = (x[52]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[52]);
  assign t[191] = (x[55]);
  assign t[192] = (x[55]);
  assign t[193] = (x[58]);
  assign t[194] = (x[58]);
  assign t[195] = (x[61]);
  assign t[196] = (x[61]);
  assign t[197] = (x[64]);
  assign t[198] = (x[64]);
  assign t[199] = (x[67]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = (x[67]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[45] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[41] : t[5];
  assign t[30] = ~(t[52] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[43]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[42] ^ t[39];
  assign t[36] = ~(t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[63]);
  assign t[41] = (t[64]);
  assign t[42] = (t[65]);
  assign t[43] = (t[66]);
  assign t[44] = (t[67]);
  assign t[45] = (t[68]);
  assign t[46] = (t[69]);
  assign t[47] = (t[70]);
  assign t[48] = (t[71]);
  assign t[49] = (t[72]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[73]);
  assign t[51] = (t[74]);
  assign t[52] = (t[75]);
  assign t[53] = (t[76]);
  assign t[54] = (t[77]);
  assign t[55] = (t[78]);
  assign t[56] = (t[79]);
  assign t[57] = (t[80]);
  assign t[58] = (t[81]);
  assign t[59] = (t[82]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[83]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = t[86] ^ x[2];
  assign t[64] = t[87] ^ x[5];
  assign t[65] = t[88] ^ x[9];
  assign t[66] = t[89] ^ x[12];
  assign t[67] = t[90] ^ x[15];
  assign t[68] = t[91] ^ x[18];
  assign t[69] = t[92] ^ x[21];
  assign t[6] = ~(t[10]);
  assign t[70] = t[93] ^ x[24];
  assign t[71] = t[94] ^ x[27];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[33];
  assign t[74] = t[97] ^ x[36];
  assign t[75] = t[98] ^ x[39];
  assign t[76] = t[99] ^ x[42];
  assign t[77] = t[100] ^ x[45];
  assign t[78] = t[101] ^ x[48];
  assign t[79] = t[102] ^ x[51];
  assign t[7] = ~(t[11]);
  assign t[80] = t[103] ^ x[54];
  assign t[81] = t[104] ^ x[57];
  assign t[82] = t[105] ^ x[60];
  assign t[83] = t[106] ^ x[63];
  assign t[84] = t[107] ^ x[66];
  assign t[85] = t[108] ^ x[69];
  assign t[86] = (t[109] & ~t[110]);
  assign t[87] = (t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[114]);
  assign t[89] = (t[115] & ~t[116]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[117] & ~t[118]);
  assign t[91] = (t[119] & ~t[120]);
  assign t[92] = (t[121] & ~t[122]);
  assign t[93] = (t[123] & ~t[124]);
  assign t[94] = (t[125] & ~t[126]);
  assign t[95] = (t[127] & ~t[128]);
  assign t[96] = (t[129] & ~t[130]);
  assign t[97] = (t[131] & ~t[132]);
  assign t[98] = (t[133] & ~t[134]);
  assign t[99] = (t[135] & ~t[136]);
  assign t[9] = t[13] ? t[14] : t[42];
  assign y = (t[0]);
endmodule

module R2ind476(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind477(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind478(x, y);
 input [69:0] x;
 output y;

 wire [200:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[137] & ~t[138]);
  assign t[101] = (t[139] & ~t[140]);
  assign t[102] = (t[141] & ~t[142]);
  assign t[103] = (t[143] & ~t[144]);
  assign t[104] = (t[145] & ~t[146]);
  assign t[105] = (t[147] & ~t[148]);
  assign t[106] = (t[149] & ~t[150]);
  assign t[107] = (t[151] & ~t[152]);
  assign t[108] = (t[153] & ~t[154]);
  assign t[109] = t[155] ^ x[2];
  assign t[10] = t[43] & t[15];
  assign t[110] = t[156] ^ x[1];
  assign t[111] = t[157] ^ x[5];
  assign t[112] = t[158] ^ x[4];
  assign t[113] = t[159] ^ x[9];
  assign t[114] = t[160] ^ x[8];
  assign t[115] = t[161] ^ x[12];
  assign t[116] = t[162] ^ x[11];
  assign t[117] = t[163] ^ x[15];
  assign t[118] = t[164] ^ x[14];
  assign t[119] = t[165] ^ x[18];
  assign t[11] = ~(t[16]);
  assign t[120] = t[166] ^ x[17];
  assign t[121] = t[167] ^ x[21];
  assign t[122] = t[168] ^ x[20];
  assign t[123] = t[169] ^ x[24];
  assign t[124] = t[170] ^ x[23];
  assign t[125] = t[171] ^ x[27];
  assign t[126] = t[172] ^ x[26];
  assign t[127] = t[173] ^ x[30];
  assign t[128] = t[174] ^ x[29];
  assign t[129] = t[175] ^ x[33];
  assign t[12] = ~(t[43]);
  assign t[130] = t[176] ^ x[32];
  assign t[131] = t[177] ^ x[36];
  assign t[132] = t[178] ^ x[35];
  assign t[133] = t[179] ^ x[39];
  assign t[134] = t[180] ^ x[38];
  assign t[135] = t[181] ^ x[42];
  assign t[136] = t[182] ^ x[41];
  assign t[137] = t[183] ^ x[45];
  assign t[138] = t[184] ^ x[44];
  assign t[139] = t[185] ^ x[48];
  assign t[13] = ~(t[17]);
  assign t[140] = t[186] ^ x[47];
  assign t[141] = t[187] ^ x[51];
  assign t[142] = t[188] ^ x[50];
  assign t[143] = t[189] ^ x[54];
  assign t[144] = t[190] ^ x[53];
  assign t[145] = t[191] ^ x[57];
  assign t[146] = t[192] ^ x[56];
  assign t[147] = t[193] ^ x[60];
  assign t[148] = t[194] ^ x[59];
  assign t[149] = t[195] ^ x[63];
  assign t[14] = t[18] ? t[44] : t[19];
  assign t[150] = t[196] ^ x[62];
  assign t[151] = t[197] ^ x[66];
  assign t[152] = t[198] ^ x[65];
  assign t[153] = t[199] ^ x[69];
  assign t[154] = t[200] ^ x[68];
  assign t[155] = (x[0]);
  assign t[156] = (x[0]);
  assign t[157] = (x[3]);
  assign t[158] = (x[3]);
  assign t[159] = (x[7]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[7]);
  assign t[161] = (x[10]);
  assign t[162] = (x[10]);
  assign t[163] = (x[13]);
  assign t[164] = (x[13]);
  assign t[165] = (x[16]);
  assign t[166] = (x[16]);
  assign t[167] = (x[19]);
  assign t[168] = (x[19]);
  assign t[169] = (x[22]);
  assign t[16] = ~(t[43] & t[22]);
  assign t[170] = (x[22]);
  assign t[171] = (x[25]);
  assign t[172] = (x[25]);
  assign t[173] = (x[28]);
  assign t[174] = (x[28]);
  assign t[175] = (x[31]);
  assign t[176] = (x[31]);
  assign t[177] = (x[34]);
  assign t[178] = (x[34]);
  assign t[179] = (x[37]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[37]);
  assign t[181] = (x[40]);
  assign t[182] = (x[40]);
  assign t[183] = (x[43]);
  assign t[184] = (x[43]);
  assign t[185] = (x[46]);
  assign t[186] = (x[46]);
  assign t[187] = (x[49]);
  assign t[188] = (x[49]);
  assign t[189] = (x[52]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[52]);
  assign t[191] = (x[55]);
  assign t[192] = (x[55]);
  assign t[193] = (x[58]);
  assign t[194] = (x[58]);
  assign t[195] = (x[61]);
  assign t[196] = (x[61]);
  assign t[197] = (x[64]);
  assign t[198] = (x[64]);
  assign t[199] = (x[67]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = (x[67]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[45] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[41] : t[5];
  assign t[30] = ~(t[52] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[43]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[42] ^ t[39];
  assign t[36] = ~(t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[63]);
  assign t[41] = (t[64]);
  assign t[42] = (t[65]);
  assign t[43] = (t[66]);
  assign t[44] = (t[67]);
  assign t[45] = (t[68]);
  assign t[46] = (t[69]);
  assign t[47] = (t[70]);
  assign t[48] = (t[71]);
  assign t[49] = (t[72]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[73]);
  assign t[51] = (t[74]);
  assign t[52] = (t[75]);
  assign t[53] = (t[76]);
  assign t[54] = (t[77]);
  assign t[55] = (t[78]);
  assign t[56] = (t[79]);
  assign t[57] = (t[80]);
  assign t[58] = (t[81]);
  assign t[59] = (t[82]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[83]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = t[86] ^ x[2];
  assign t[64] = t[87] ^ x[5];
  assign t[65] = t[88] ^ x[9];
  assign t[66] = t[89] ^ x[12];
  assign t[67] = t[90] ^ x[15];
  assign t[68] = t[91] ^ x[18];
  assign t[69] = t[92] ^ x[21];
  assign t[6] = ~(t[10]);
  assign t[70] = t[93] ^ x[24];
  assign t[71] = t[94] ^ x[27];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[33];
  assign t[74] = t[97] ^ x[36];
  assign t[75] = t[98] ^ x[39];
  assign t[76] = t[99] ^ x[42];
  assign t[77] = t[100] ^ x[45];
  assign t[78] = t[101] ^ x[48];
  assign t[79] = t[102] ^ x[51];
  assign t[7] = ~(t[11]);
  assign t[80] = t[103] ^ x[54];
  assign t[81] = t[104] ^ x[57];
  assign t[82] = t[105] ^ x[60];
  assign t[83] = t[106] ^ x[63];
  assign t[84] = t[107] ^ x[66];
  assign t[85] = t[108] ^ x[69];
  assign t[86] = (t[109] & ~t[110]);
  assign t[87] = (t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[114]);
  assign t[89] = (t[115] & ~t[116]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[117] & ~t[118]);
  assign t[91] = (t[119] & ~t[120]);
  assign t[92] = (t[121] & ~t[122]);
  assign t[93] = (t[123] & ~t[124]);
  assign t[94] = (t[125] & ~t[126]);
  assign t[95] = (t[127] & ~t[128]);
  assign t[96] = (t[129] & ~t[130]);
  assign t[97] = (t[131] & ~t[132]);
  assign t[98] = (t[133] & ~t[134]);
  assign t[99] = (t[135] & ~t[136]);
  assign t[9] = t[13] ? t[14] : t[42];
  assign y = (t[0]);
endmodule

module R2ind479(x, y);
 input [69:0] x;
 output y;

 wire [200:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[137] & ~t[138]);
  assign t[101] = (t[139] & ~t[140]);
  assign t[102] = (t[141] & ~t[142]);
  assign t[103] = (t[143] & ~t[144]);
  assign t[104] = (t[145] & ~t[146]);
  assign t[105] = (t[147] & ~t[148]);
  assign t[106] = (t[149] & ~t[150]);
  assign t[107] = (t[151] & ~t[152]);
  assign t[108] = (t[153] & ~t[154]);
  assign t[109] = t[155] ^ x[2];
  assign t[10] = t[43] & t[15];
  assign t[110] = t[156] ^ x[1];
  assign t[111] = t[157] ^ x[5];
  assign t[112] = t[158] ^ x[4];
  assign t[113] = t[159] ^ x[9];
  assign t[114] = t[160] ^ x[8];
  assign t[115] = t[161] ^ x[12];
  assign t[116] = t[162] ^ x[11];
  assign t[117] = t[163] ^ x[15];
  assign t[118] = t[164] ^ x[14];
  assign t[119] = t[165] ^ x[18];
  assign t[11] = ~(t[16]);
  assign t[120] = t[166] ^ x[17];
  assign t[121] = t[167] ^ x[21];
  assign t[122] = t[168] ^ x[20];
  assign t[123] = t[169] ^ x[24];
  assign t[124] = t[170] ^ x[23];
  assign t[125] = t[171] ^ x[27];
  assign t[126] = t[172] ^ x[26];
  assign t[127] = t[173] ^ x[30];
  assign t[128] = t[174] ^ x[29];
  assign t[129] = t[175] ^ x[33];
  assign t[12] = ~(t[43]);
  assign t[130] = t[176] ^ x[32];
  assign t[131] = t[177] ^ x[36];
  assign t[132] = t[178] ^ x[35];
  assign t[133] = t[179] ^ x[39];
  assign t[134] = t[180] ^ x[38];
  assign t[135] = t[181] ^ x[42];
  assign t[136] = t[182] ^ x[41];
  assign t[137] = t[183] ^ x[45];
  assign t[138] = t[184] ^ x[44];
  assign t[139] = t[185] ^ x[48];
  assign t[13] = ~(t[17]);
  assign t[140] = t[186] ^ x[47];
  assign t[141] = t[187] ^ x[51];
  assign t[142] = t[188] ^ x[50];
  assign t[143] = t[189] ^ x[54];
  assign t[144] = t[190] ^ x[53];
  assign t[145] = t[191] ^ x[57];
  assign t[146] = t[192] ^ x[56];
  assign t[147] = t[193] ^ x[60];
  assign t[148] = t[194] ^ x[59];
  assign t[149] = t[195] ^ x[63];
  assign t[14] = t[18] ? t[44] : t[19];
  assign t[150] = t[196] ^ x[62];
  assign t[151] = t[197] ^ x[66];
  assign t[152] = t[198] ^ x[65];
  assign t[153] = t[199] ^ x[69];
  assign t[154] = t[200] ^ x[68];
  assign t[155] = (x[0]);
  assign t[156] = (x[0]);
  assign t[157] = (x[3]);
  assign t[158] = (x[3]);
  assign t[159] = (x[7]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[7]);
  assign t[161] = (x[10]);
  assign t[162] = (x[10]);
  assign t[163] = (x[13]);
  assign t[164] = (x[13]);
  assign t[165] = (x[16]);
  assign t[166] = (x[16]);
  assign t[167] = (x[19]);
  assign t[168] = (x[19]);
  assign t[169] = (x[22]);
  assign t[16] = ~(t[43] & t[22]);
  assign t[170] = (x[22]);
  assign t[171] = (x[25]);
  assign t[172] = (x[25]);
  assign t[173] = (x[28]);
  assign t[174] = (x[28]);
  assign t[175] = (x[31]);
  assign t[176] = (x[31]);
  assign t[177] = (x[34]);
  assign t[178] = (x[34]);
  assign t[179] = (x[37]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[37]);
  assign t[181] = (x[40]);
  assign t[182] = (x[40]);
  assign t[183] = (x[43]);
  assign t[184] = (x[43]);
  assign t[185] = (x[46]);
  assign t[186] = (x[46]);
  assign t[187] = (x[49]);
  assign t[188] = (x[49]);
  assign t[189] = (x[52]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[52]);
  assign t[191] = (x[55]);
  assign t[192] = (x[55]);
  assign t[193] = (x[58]);
  assign t[194] = (x[58]);
  assign t[195] = (x[61]);
  assign t[196] = (x[61]);
  assign t[197] = (x[64]);
  assign t[198] = (x[64]);
  assign t[199] = (x[67]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = (x[67]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[45] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[41] : t[5];
  assign t[30] = ~(t[52] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[43]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[42] ^ t[39];
  assign t[36] = ~(t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[63]);
  assign t[41] = (t[64]);
  assign t[42] = (t[65]);
  assign t[43] = (t[66]);
  assign t[44] = (t[67]);
  assign t[45] = (t[68]);
  assign t[46] = (t[69]);
  assign t[47] = (t[70]);
  assign t[48] = (t[71]);
  assign t[49] = (t[72]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[73]);
  assign t[51] = (t[74]);
  assign t[52] = (t[75]);
  assign t[53] = (t[76]);
  assign t[54] = (t[77]);
  assign t[55] = (t[78]);
  assign t[56] = (t[79]);
  assign t[57] = (t[80]);
  assign t[58] = (t[81]);
  assign t[59] = (t[82]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[83]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = t[86] ^ x[2];
  assign t[64] = t[87] ^ x[5];
  assign t[65] = t[88] ^ x[9];
  assign t[66] = t[89] ^ x[12];
  assign t[67] = t[90] ^ x[15];
  assign t[68] = t[91] ^ x[18];
  assign t[69] = t[92] ^ x[21];
  assign t[6] = ~(t[10]);
  assign t[70] = t[93] ^ x[24];
  assign t[71] = t[94] ^ x[27];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[33];
  assign t[74] = t[97] ^ x[36];
  assign t[75] = t[98] ^ x[39];
  assign t[76] = t[99] ^ x[42];
  assign t[77] = t[100] ^ x[45];
  assign t[78] = t[101] ^ x[48];
  assign t[79] = t[102] ^ x[51];
  assign t[7] = ~(t[11]);
  assign t[80] = t[103] ^ x[54];
  assign t[81] = t[104] ^ x[57];
  assign t[82] = t[105] ^ x[60];
  assign t[83] = t[106] ^ x[63];
  assign t[84] = t[107] ^ x[66];
  assign t[85] = t[108] ^ x[69];
  assign t[86] = (t[109] & ~t[110]);
  assign t[87] = (t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[114]);
  assign t[89] = (t[115] & ~t[116]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[117] & ~t[118]);
  assign t[91] = (t[119] & ~t[120]);
  assign t[92] = (t[121] & ~t[122]);
  assign t[93] = (t[123] & ~t[124]);
  assign t[94] = (t[125] & ~t[126]);
  assign t[95] = (t[127] & ~t[128]);
  assign t[96] = (t[129] & ~t[130]);
  assign t[97] = (t[131] & ~t[132]);
  assign t[98] = (t[133] & ~t[134]);
  assign t[99] = (t[135] & ~t[136]);
  assign t[9] = t[13] ? t[14] : t[42];
  assign y = (t[0]);
endmodule

module R2ind480(x, y);
 input [69:0] x;
 output y;

 wire [200:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[137] & ~t[138]);
  assign t[101] = (t[139] & ~t[140]);
  assign t[102] = (t[141] & ~t[142]);
  assign t[103] = (t[143] & ~t[144]);
  assign t[104] = (t[145] & ~t[146]);
  assign t[105] = (t[147] & ~t[148]);
  assign t[106] = (t[149] & ~t[150]);
  assign t[107] = (t[151] & ~t[152]);
  assign t[108] = (t[153] & ~t[154]);
  assign t[109] = t[155] ^ x[2];
  assign t[10] = t[43] & t[15];
  assign t[110] = t[156] ^ x[1];
  assign t[111] = t[157] ^ x[5];
  assign t[112] = t[158] ^ x[4];
  assign t[113] = t[159] ^ x[9];
  assign t[114] = t[160] ^ x[8];
  assign t[115] = t[161] ^ x[12];
  assign t[116] = t[162] ^ x[11];
  assign t[117] = t[163] ^ x[15];
  assign t[118] = t[164] ^ x[14];
  assign t[119] = t[165] ^ x[18];
  assign t[11] = ~(t[16]);
  assign t[120] = t[166] ^ x[17];
  assign t[121] = t[167] ^ x[21];
  assign t[122] = t[168] ^ x[20];
  assign t[123] = t[169] ^ x[24];
  assign t[124] = t[170] ^ x[23];
  assign t[125] = t[171] ^ x[27];
  assign t[126] = t[172] ^ x[26];
  assign t[127] = t[173] ^ x[30];
  assign t[128] = t[174] ^ x[29];
  assign t[129] = t[175] ^ x[33];
  assign t[12] = ~(t[43]);
  assign t[130] = t[176] ^ x[32];
  assign t[131] = t[177] ^ x[36];
  assign t[132] = t[178] ^ x[35];
  assign t[133] = t[179] ^ x[39];
  assign t[134] = t[180] ^ x[38];
  assign t[135] = t[181] ^ x[42];
  assign t[136] = t[182] ^ x[41];
  assign t[137] = t[183] ^ x[45];
  assign t[138] = t[184] ^ x[44];
  assign t[139] = t[185] ^ x[48];
  assign t[13] = ~(t[17]);
  assign t[140] = t[186] ^ x[47];
  assign t[141] = t[187] ^ x[51];
  assign t[142] = t[188] ^ x[50];
  assign t[143] = t[189] ^ x[54];
  assign t[144] = t[190] ^ x[53];
  assign t[145] = t[191] ^ x[57];
  assign t[146] = t[192] ^ x[56];
  assign t[147] = t[193] ^ x[60];
  assign t[148] = t[194] ^ x[59];
  assign t[149] = t[195] ^ x[63];
  assign t[14] = t[18] ? t[44] : t[19];
  assign t[150] = t[196] ^ x[62];
  assign t[151] = t[197] ^ x[66];
  assign t[152] = t[198] ^ x[65];
  assign t[153] = t[199] ^ x[69];
  assign t[154] = t[200] ^ x[68];
  assign t[155] = (x[0]);
  assign t[156] = (x[0]);
  assign t[157] = (x[3]);
  assign t[158] = (x[3]);
  assign t[159] = (x[7]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[7]);
  assign t[161] = (x[10]);
  assign t[162] = (x[10]);
  assign t[163] = (x[13]);
  assign t[164] = (x[13]);
  assign t[165] = (x[16]);
  assign t[166] = (x[16]);
  assign t[167] = (x[19]);
  assign t[168] = (x[19]);
  assign t[169] = (x[22]);
  assign t[16] = ~(t[43] & t[22]);
  assign t[170] = (x[22]);
  assign t[171] = (x[25]);
  assign t[172] = (x[25]);
  assign t[173] = (x[28]);
  assign t[174] = (x[28]);
  assign t[175] = (x[31]);
  assign t[176] = (x[31]);
  assign t[177] = (x[34]);
  assign t[178] = (x[34]);
  assign t[179] = (x[37]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[37]);
  assign t[181] = (x[40]);
  assign t[182] = (x[40]);
  assign t[183] = (x[43]);
  assign t[184] = (x[43]);
  assign t[185] = (x[46]);
  assign t[186] = (x[46]);
  assign t[187] = (x[49]);
  assign t[188] = (x[49]);
  assign t[189] = (x[52]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[52]);
  assign t[191] = (x[55]);
  assign t[192] = (x[55]);
  assign t[193] = (x[58]);
  assign t[194] = (x[58]);
  assign t[195] = (x[61]);
  assign t[196] = (x[61]);
  assign t[197] = (x[64]);
  assign t[198] = (x[64]);
  assign t[199] = (x[67]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = (x[67]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[45] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[41] : t[5];
  assign t[30] = ~(t[52] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[43]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[42] ^ t[39];
  assign t[36] = ~(t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[63]);
  assign t[41] = (t[64]);
  assign t[42] = (t[65]);
  assign t[43] = (t[66]);
  assign t[44] = (t[67]);
  assign t[45] = (t[68]);
  assign t[46] = (t[69]);
  assign t[47] = (t[70]);
  assign t[48] = (t[71]);
  assign t[49] = (t[72]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[73]);
  assign t[51] = (t[74]);
  assign t[52] = (t[75]);
  assign t[53] = (t[76]);
  assign t[54] = (t[77]);
  assign t[55] = (t[78]);
  assign t[56] = (t[79]);
  assign t[57] = (t[80]);
  assign t[58] = (t[81]);
  assign t[59] = (t[82]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[83]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = t[86] ^ x[2];
  assign t[64] = t[87] ^ x[5];
  assign t[65] = t[88] ^ x[9];
  assign t[66] = t[89] ^ x[12];
  assign t[67] = t[90] ^ x[15];
  assign t[68] = t[91] ^ x[18];
  assign t[69] = t[92] ^ x[21];
  assign t[6] = ~(t[10]);
  assign t[70] = t[93] ^ x[24];
  assign t[71] = t[94] ^ x[27];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[33];
  assign t[74] = t[97] ^ x[36];
  assign t[75] = t[98] ^ x[39];
  assign t[76] = t[99] ^ x[42];
  assign t[77] = t[100] ^ x[45];
  assign t[78] = t[101] ^ x[48];
  assign t[79] = t[102] ^ x[51];
  assign t[7] = ~(t[11]);
  assign t[80] = t[103] ^ x[54];
  assign t[81] = t[104] ^ x[57];
  assign t[82] = t[105] ^ x[60];
  assign t[83] = t[106] ^ x[63];
  assign t[84] = t[107] ^ x[66];
  assign t[85] = t[108] ^ x[69];
  assign t[86] = (t[109] & ~t[110]);
  assign t[87] = (t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[114]);
  assign t[89] = (t[115] & ~t[116]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[117] & ~t[118]);
  assign t[91] = (t[119] & ~t[120]);
  assign t[92] = (t[121] & ~t[122]);
  assign t[93] = (t[123] & ~t[124]);
  assign t[94] = (t[125] & ~t[126]);
  assign t[95] = (t[127] & ~t[128]);
  assign t[96] = (t[129] & ~t[130]);
  assign t[97] = (t[131] & ~t[132]);
  assign t[98] = (t[133] & ~t[134]);
  assign t[99] = (t[135] & ~t[136]);
  assign t[9] = t[13] ? t[14] : t[42];
  assign y = (t[0]);
endmodule

module R2ind481(x, y);
 input [69:0] x;
 output y;

 wire [200:0] t;
  assign t[0] = t[1] ? t[2] : t[40];
  assign t[100] = (t[137] & ~t[138]);
  assign t[101] = (t[139] & ~t[140]);
  assign t[102] = (t[141] & ~t[142]);
  assign t[103] = (t[143] & ~t[144]);
  assign t[104] = (t[145] & ~t[146]);
  assign t[105] = (t[147] & ~t[148]);
  assign t[106] = (t[149] & ~t[150]);
  assign t[107] = (t[151] & ~t[152]);
  assign t[108] = (t[153] & ~t[154]);
  assign t[109] = t[155] ^ x[2];
  assign t[10] = t[43] & t[15];
  assign t[110] = t[156] ^ x[1];
  assign t[111] = t[157] ^ x[5];
  assign t[112] = t[158] ^ x[4];
  assign t[113] = t[159] ^ x[9];
  assign t[114] = t[160] ^ x[8];
  assign t[115] = t[161] ^ x[12];
  assign t[116] = t[162] ^ x[11];
  assign t[117] = t[163] ^ x[15];
  assign t[118] = t[164] ^ x[14];
  assign t[119] = t[165] ^ x[18];
  assign t[11] = ~(t[16]);
  assign t[120] = t[166] ^ x[17];
  assign t[121] = t[167] ^ x[21];
  assign t[122] = t[168] ^ x[20];
  assign t[123] = t[169] ^ x[24];
  assign t[124] = t[170] ^ x[23];
  assign t[125] = t[171] ^ x[27];
  assign t[126] = t[172] ^ x[26];
  assign t[127] = t[173] ^ x[30];
  assign t[128] = t[174] ^ x[29];
  assign t[129] = t[175] ^ x[33];
  assign t[12] = ~(t[43]);
  assign t[130] = t[176] ^ x[32];
  assign t[131] = t[177] ^ x[36];
  assign t[132] = t[178] ^ x[35];
  assign t[133] = t[179] ^ x[39];
  assign t[134] = t[180] ^ x[38];
  assign t[135] = t[181] ^ x[42];
  assign t[136] = t[182] ^ x[41];
  assign t[137] = t[183] ^ x[45];
  assign t[138] = t[184] ^ x[44];
  assign t[139] = t[185] ^ x[48];
  assign t[13] = ~(t[17]);
  assign t[140] = t[186] ^ x[47];
  assign t[141] = t[187] ^ x[51];
  assign t[142] = t[188] ^ x[50];
  assign t[143] = t[189] ^ x[54];
  assign t[144] = t[190] ^ x[53];
  assign t[145] = t[191] ^ x[57];
  assign t[146] = t[192] ^ x[56];
  assign t[147] = t[193] ^ x[60];
  assign t[148] = t[194] ^ x[59];
  assign t[149] = t[195] ^ x[63];
  assign t[14] = t[18] ? t[44] : t[19];
  assign t[150] = t[196] ^ x[62];
  assign t[151] = t[197] ^ x[66];
  assign t[152] = t[198] ^ x[65];
  assign t[153] = t[199] ^ x[69];
  assign t[154] = t[200] ^ x[68];
  assign t[155] = (x[0]);
  assign t[156] = (x[0]);
  assign t[157] = (x[3]);
  assign t[158] = (x[3]);
  assign t[159] = (x[7]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[7]);
  assign t[161] = (x[10]);
  assign t[162] = (x[10]);
  assign t[163] = (x[13]);
  assign t[164] = (x[13]);
  assign t[165] = (x[16]);
  assign t[166] = (x[16]);
  assign t[167] = (x[19]);
  assign t[168] = (x[19]);
  assign t[169] = (x[22]);
  assign t[16] = ~(t[43] & t[22]);
  assign t[170] = (x[22]);
  assign t[171] = (x[25]);
  assign t[172] = (x[25]);
  assign t[173] = (x[28]);
  assign t[174] = (x[28]);
  assign t[175] = (x[31]);
  assign t[176] = (x[31]);
  assign t[177] = (x[34]);
  assign t[178] = (x[34]);
  assign t[179] = (x[37]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[37]);
  assign t[181] = (x[40]);
  assign t[182] = (x[40]);
  assign t[183] = (x[43]);
  assign t[184] = (x[43]);
  assign t[185] = (x[46]);
  assign t[186] = (x[46]);
  assign t[187] = (x[49]);
  assign t[188] = (x[49]);
  assign t[189] = (x[52]);
  assign t[18] = ~(t[24]);
  assign t[190] = (x[52]);
  assign t[191] = (x[55]);
  assign t[192] = (x[55]);
  assign t[193] = (x[58]);
  assign t[194] = (x[58]);
  assign t[195] = (x[61]);
  assign t[196] = (x[61]);
  assign t[197] = (x[64]);
  assign t[198] = (x[64]);
  assign t[199] = (x[67]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[200] = (x[67]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[45] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[34] ^ t[35];
  assign t[26] = ~(t[46] ^ t[47]);
  assign t[27] = ~(t[48] & t[49]);
  assign t[28] = ~(t[50] & t[51]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[41] : t[5];
  assign t[30] = ~(t[52] & t[36]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[53]);
  assign t[33] = ~(t[43]);
  assign t[34] = t[54] ^ t[55];
  assign t[35] = t[42] ^ t[39];
  assign t[36] = ~(t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = ~(t[59] | t[60]);
  assign t[39] = t[61] ^ t[62];
  assign t[3] = ~(t[6]);
  assign t[40] = (t[63]);
  assign t[41] = (t[64]);
  assign t[42] = (t[65]);
  assign t[43] = (t[66]);
  assign t[44] = (t[67]);
  assign t[45] = (t[68]);
  assign t[46] = (t[69]);
  assign t[47] = (t[70]);
  assign t[48] = (t[71]);
  assign t[49] = (t[72]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[73]);
  assign t[51] = (t[74]);
  assign t[52] = (t[75]);
  assign t[53] = (t[76]);
  assign t[54] = (t[77]);
  assign t[55] = (t[78]);
  assign t[56] = (t[79]);
  assign t[57] = (t[80]);
  assign t[58] = (t[81]);
  assign t[59] = (t[82]);
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = (t[83]);
  assign t[61] = (t[84]);
  assign t[62] = (t[85]);
  assign t[63] = t[86] ^ x[2];
  assign t[64] = t[87] ^ x[5];
  assign t[65] = t[88] ^ x[9];
  assign t[66] = t[89] ^ x[12];
  assign t[67] = t[90] ^ x[15];
  assign t[68] = t[91] ^ x[18];
  assign t[69] = t[92] ^ x[21];
  assign t[6] = ~(t[10]);
  assign t[70] = t[93] ^ x[24];
  assign t[71] = t[94] ^ x[27];
  assign t[72] = t[95] ^ x[30];
  assign t[73] = t[96] ^ x[33];
  assign t[74] = t[97] ^ x[36];
  assign t[75] = t[98] ^ x[39];
  assign t[76] = t[99] ^ x[42];
  assign t[77] = t[100] ^ x[45];
  assign t[78] = t[101] ^ x[48];
  assign t[79] = t[102] ^ x[51];
  assign t[7] = ~(t[11]);
  assign t[80] = t[103] ^ x[54];
  assign t[81] = t[104] ^ x[57];
  assign t[82] = t[105] ^ x[60];
  assign t[83] = t[106] ^ x[63];
  assign t[84] = t[107] ^ x[66];
  assign t[85] = t[108] ^ x[69];
  assign t[86] = (t[109] & ~t[110]);
  assign t[87] = (t[111] & ~t[112]);
  assign t[88] = (t[113] & ~t[114]);
  assign t[89] = (t[115] & ~t[116]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[117] & ~t[118]);
  assign t[91] = (t[119] & ~t[120]);
  assign t[92] = (t[121] & ~t[122]);
  assign t[93] = (t[123] & ~t[124]);
  assign t[94] = (t[125] & ~t[126]);
  assign t[95] = (t[127] & ~t[128]);
  assign t[96] = (t[129] & ~t[130]);
  assign t[97] = (t[131] & ~t[132]);
  assign t[98] = (t[133] & ~t[134]);
  assign t[99] = (t[135] & ~t[136]);
  assign t[9] = t[13] ? t[14] : t[42];
  assign y = (t[0]);
endmodule

module R2ind482(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind483(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind484(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind485(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind486(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind487(x, y);
 input [63:0] x;
 output y;

 wire [184:0] t;
  assign t[0] = t[1] ? t[2] : t[38];
  assign t[100] = (t[141] & ~t[142]);
  assign t[101] = t[143] ^ x[2];
  assign t[102] = t[144] ^ x[1];
  assign t[103] = t[145] ^ x[5];
  assign t[104] = t[146] ^ x[4];
  assign t[105] = t[147] ^ x[9];
  assign t[106] = t[148] ^ x[8];
  assign t[107] = t[149] ^ x[12];
  assign t[108] = t[150] ^ x[11];
  assign t[109] = t[151] ^ x[15];
  assign t[10] = t[41] & t[15];
  assign t[110] = t[152] ^ x[14];
  assign t[111] = t[153] ^ x[18];
  assign t[112] = t[154] ^ x[17];
  assign t[113] = t[155] ^ x[21];
  assign t[114] = t[156] ^ x[20];
  assign t[115] = t[157] ^ x[24];
  assign t[116] = t[158] ^ x[23];
  assign t[117] = t[159] ^ x[27];
  assign t[118] = t[160] ^ x[26];
  assign t[119] = t[161] ^ x[30];
  assign t[11] = ~(t[16]);
  assign t[120] = t[162] ^ x[29];
  assign t[121] = t[163] ^ x[33];
  assign t[122] = t[164] ^ x[32];
  assign t[123] = t[165] ^ x[36];
  assign t[124] = t[166] ^ x[35];
  assign t[125] = t[167] ^ x[39];
  assign t[126] = t[168] ^ x[38];
  assign t[127] = t[169] ^ x[42];
  assign t[128] = t[170] ^ x[41];
  assign t[129] = t[171] ^ x[45];
  assign t[12] = ~(t[41]);
  assign t[130] = t[172] ^ x[44];
  assign t[131] = t[173] ^ x[48];
  assign t[132] = t[174] ^ x[47];
  assign t[133] = t[175] ^ x[51];
  assign t[134] = t[176] ^ x[50];
  assign t[135] = t[177] ^ x[54];
  assign t[136] = t[178] ^ x[53];
  assign t[137] = t[179] ^ x[57];
  assign t[138] = t[180] ^ x[56];
  assign t[139] = t[181] ^ x[60];
  assign t[13] = ~(t[17]);
  assign t[140] = t[182] ^ x[59];
  assign t[141] = t[183] ^ x[63];
  assign t[142] = t[184] ^ x[62];
  assign t[143] = (x[0]);
  assign t[144] = (x[0]);
  assign t[145] = (x[3]);
  assign t[146] = (x[3]);
  assign t[147] = (x[7]);
  assign t[148] = (x[7]);
  assign t[149] = (x[10]);
  assign t[14] = t[18] ? t[42] : t[19];
  assign t[150] = (x[10]);
  assign t[151] = (x[13]);
  assign t[152] = (x[13]);
  assign t[153] = (x[16]);
  assign t[154] = (x[16]);
  assign t[155] = (x[19]);
  assign t[156] = (x[19]);
  assign t[157] = (x[22]);
  assign t[158] = (x[22]);
  assign t[159] = (x[25]);
  assign t[15] = t[20] & t[21];
  assign t[160] = (x[25]);
  assign t[161] = (x[28]);
  assign t[162] = (x[28]);
  assign t[163] = (x[31]);
  assign t[164] = (x[31]);
  assign t[165] = (x[34]);
  assign t[166] = (x[34]);
  assign t[167] = (x[37]);
  assign t[168] = (x[37]);
  assign t[169] = (x[40]);
  assign t[16] = ~(t[41] & t[22]);
  assign t[170] = (x[40]);
  assign t[171] = (x[43]);
  assign t[172] = (x[43]);
  assign t[173] = (x[46]);
  assign t[174] = (x[46]);
  assign t[175] = (x[49]);
  assign t[176] = (x[49]);
  assign t[177] = (x[52]);
  assign t[178] = (x[52]);
  assign t[179] = (x[55]);
  assign t[17] = ~(t[23]);
  assign t[180] = (x[55]);
  assign t[181] = (x[58]);
  assign t[182] = (x[58]);
  assign t[183] = (x[61]);
  assign t[184] = (x[61]);
  assign t[18] = ~(t[24]);
  assign t[19] = ~(t[25] ^ t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[30]);
  assign t[22] = ~(t[43] | t[31]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[24] = ~(t[20]);
  assign t[25] = t[44] ^ t[34];
  assign t[26] = ~(t[45] ^ t[46]);
  assign t[27] = ~(t[47] & t[48]);
  assign t[28] = ~(t[49] & t[50]);
  assign t[29] = ~(t[22]);
  assign t[2] = t[4] ? t[39] : t[5];
  assign t[30] = ~(t[51] & t[35]);
  assign t[31] = ~(t[36] & t[37]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[41]);
  assign t[34] = t[40] ^ t[53];
  assign t[35] = ~(t[54]);
  assign t[36] = ~(t[55] | t[56]);
  assign t[37] = ~(t[57] | t[58]);
  assign t[38] = (t[59]);
  assign t[39] = (t[60]);
  assign t[3] = ~(t[6]);
  assign t[40] = (t[61]);
  assign t[41] = (t[62]);
  assign t[42] = (t[63]);
  assign t[43] = (t[64]);
  assign t[44] = (t[65]);
  assign t[45] = (t[66]);
  assign t[46] = (t[67]);
  assign t[47] = (t[68]);
  assign t[48] = (t[69]);
  assign t[49] = (t[70]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[71]);
  assign t[51] = (t[72]);
  assign t[52] = (t[73]);
  assign t[53] = (t[74]);
  assign t[54] = (t[75]);
  assign t[55] = (t[76]);
  assign t[56] = (t[77]);
  assign t[57] = (t[78]);
  assign t[58] = (t[79]);
  assign t[59] = t[80] ^ x[2];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[81] ^ x[5];
  assign t[61] = t[82] ^ x[9];
  assign t[62] = t[83] ^ x[12];
  assign t[63] = t[84] ^ x[15];
  assign t[64] = t[85] ^ x[18];
  assign t[65] = t[86] ^ x[21];
  assign t[66] = t[87] ^ x[24];
  assign t[67] = t[88] ^ x[27];
  assign t[68] = t[89] ^ x[30];
  assign t[69] = t[90] ^ x[33];
  assign t[6] = ~(t[10]);
  assign t[70] = t[91] ^ x[36];
  assign t[71] = t[92] ^ x[39];
  assign t[72] = t[93] ^ x[42];
  assign t[73] = t[94] ^ x[45];
  assign t[74] = t[95] ^ x[48];
  assign t[75] = t[96] ^ x[51];
  assign t[76] = t[97] ^ x[54];
  assign t[77] = t[98] ^ x[57];
  assign t[78] = t[99] ^ x[60];
  assign t[79] = t[100] ^ x[63];
  assign t[7] = ~(t[11]);
  assign t[80] = (t[101] & ~t[102]);
  assign t[81] = (t[103] & ~t[104]);
  assign t[82] = (t[105] & ~t[106]);
  assign t[83] = (t[107] & ~t[108]);
  assign t[84] = (t[109] & ~t[110]);
  assign t[85] = (t[111] & ~t[112]);
  assign t[86] = (t[113] & ~t[114]);
  assign t[87] = (t[115] & ~t[116]);
  assign t[88] = (t[117] & ~t[118]);
  assign t[89] = (t[119] & ~t[120]);
  assign t[8] = ~(t[12]);
  assign t[90] = (t[121] & ~t[122]);
  assign t[91] = (t[123] & ~t[124]);
  assign t[92] = (t[125] & ~t[126]);
  assign t[93] = (t[127] & ~t[128]);
  assign t[94] = (t[129] & ~t[130]);
  assign t[95] = (t[131] & ~t[132]);
  assign t[96] = (t[133] & ~t[134]);
  assign t[97] = (t[135] & ~t[136]);
  assign t[98] = (t[137] & ~t[138]);
  assign t[99] = (t[139] & ~t[140]);
  assign t[9] = t[13] ? t[14] : t[40];
  assign y = (t[0]);
endmodule

module R2ind488(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind489(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind490(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind491(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind492(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind493(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind494(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind495(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind496(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind497(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind498(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind499(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind500(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind501(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind502(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind503(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind504(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind505(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind506(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind507(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind508(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind509(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind510(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind511(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind512(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind513(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind514(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind515(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind516(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind517(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind518(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind519(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind520(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind521(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind522(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind523(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind524(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind525(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind526(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind527(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind528(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind529(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind530(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind531(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind532(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind533(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind534(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind535(x, y);
 input [45:0] x;
 output y;

 wire [129:0] t;
  assign t[0] = t[1] ? t[2] : t[25];
  assign t[100] = (x[0]);
  assign t[101] = (x[0]);
  assign t[102] = (x[3]);
  assign t[103] = (x[3]);
  assign t[104] = (x[7]);
  assign t[105] = (x[7]);
  assign t[106] = (x[10]);
  assign t[107] = (x[10]);
  assign t[108] = (x[13]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[13]);
  assign t[110] = (x[16]);
  assign t[111] = (x[16]);
  assign t[112] = (x[19]);
  assign t[113] = (x[19]);
  assign t[114] = (x[22]);
  assign t[115] = (x[22]);
  assign t[116] = (x[25]);
  assign t[117] = (x[25]);
  assign t[118] = (x[28]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[28]);
  assign t[120] = (x[31]);
  assign t[121] = (x[31]);
  assign t[122] = (x[34]);
  assign t[123] = (x[34]);
  assign t[124] = (x[37]);
  assign t[125] = (x[37]);
  assign t[126] = (x[40]);
  assign t[127] = (x[40]);
  assign t[128] = (x[43]);
  assign t[129] = (x[43]);
  assign t[12] = t[14] & t[15];
  assign t[13] = ~(t[28] & t[16]);
  assign t[14] = ~(t[17] | t[18]);
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[29] | t[21]);
  assign t[17] = ~(t[30] & t[31]);
  assign t[18] = ~(t[32] & t[33]);
  assign t[19] = ~(t[16]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[34] & t[22]);
  assign t[21] = ~(t[23] & t[24]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[36] | t[37]);
  assign t[24] = ~(t[38] | t[39]);
  assign t[25] = (t[40]);
  assign t[26] = (t[41]);
  assign t[27] = (t[42]);
  assign t[28] = (t[43]);
  assign t[29] = (t[44]);
  assign t[2] = t[4] ? t[26] : t[5];
  assign t[30] = (t[45]);
  assign t[31] = (t[46]);
  assign t[32] = (t[47]);
  assign t[33] = (t[48]);
  assign t[34] = (t[49]);
  assign t[35] = (t[50]);
  assign t[36] = (t[51]);
  assign t[37] = (t[52]);
  assign t[38] = (t[53]);
  assign t[39] = (t[54]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[55] ^ x[2];
  assign t[41] = t[56] ^ x[5];
  assign t[42] = t[57] ^ x[9];
  assign t[43] = t[58] ^ x[12];
  assign t[44] = t[59] ^ x[15];
  assign t[45] = t[60] ^ x[18];
  assign t[46] = t[61] ^ x[21];
  assign t[47] = t[62] ^ x[24];
  assign t[48] = t[63] ^ x[27];
  assign t[49] = t[64] ^ x[30];
  assign t[4] = ~(t[7]);
  assign t[50] = t[65] ^ x[33];
  assign t[51] = t[66] ^ x[36];
  assign t[52] = t[67] ^ x[39];
  assign t[53] = t[68] ^ x[42];
  assign t[54] = t[69] ^ x[45];
  assign t[55] = (t[70] & ~t[71]);
  assign t[56] = (t[72] & ~t[73]);
  assign t[57] = (t[74] & ~t[75]);
  assign t[58] = (t[76] & ~t[77]);
  assign t[59] = (t[78] & ~t[79]);
  assign t[5] = t[8] ? t[27] : x[6];
  assign t[60] = (t[80] & ~t[81]);
  assign t[61] = (t[82] & ~t[83]);
  assign t[62] = (t[84] & ~t[85]);
  assign t[63] = (t[86] & ~t[87]);
  assign t[64] = (t[88] & ~t[89]);
  assign t[65] = (t[90] & ~t[91]);
  assign t[66] = (t[92] & ~t[93]);
  assign t[67] = (t[94] & ~t[95]);
  assign t[68] = (t[96] & ~t[97]);
  assign t[69] = (t[98] & ~t[99]);
  assign t[6] = ~(t[9]);
  assign t[70] = t[100] ^ x[2];
  assign t[71] = t[101] ^ x[1];
  assign t[72] = t[102] ^ x[5];
  assign t[73] = t[103] ^ x[4];
  assign t[74] = t[104] ^ x[9];
  assign t[75] = t[105] ^ x[8];
  assign t[76] = t[106] ^ x[12];
  assign t[77] = t[107] ^ x[11];
  assign t[78] = t[108] ^ x[15];
  assign t[79] = t[109] ^ x[14];
  assign t[7] = ~(t[10]);
  assign t[80] = t[110] ^ x[18];
  assign t[81] = t[111] ^ x[17];
  assign t[82] = t[112] ^ x[21];
  assign t[83] = t[113] ^ x[20];
  assign t[84] = t[114] ^ x[24];
  assign t[85] = t[115] ^ x[23];
  assign t[86] = t[116] ^ x[27];
  assign t[87] = t[117] ^ x[26];
  assign t[88] = t[118] ^ x[30];
  assign t[89] = t[119] ^ x[29];
  assign t[8] = ~(t[11]);
  assign t[90] = t[120] ^ x[33];
  assign t[91] = t[121] ^ x[32];
  assign t[92] = t[122] ^ x[36];
  assign t[93] = t[123] ^ x[35];
  assign t[94] = t[124] ^ x[39];
  assign t[95] = t[125] ^ x[38];
  assign t[96] = t[126] ^ x[42];
  assign t[97] = t[127] ^ x[41];
  assign t[98] = t[128] ^ x[45];
  assign t[99] = t[129] ^ x[44];
  assign t[9] = t[28] & t[12];
  assign y = (t[0]);
endmodule

module R2ind536(x, y);
 input [129:0] x;
 output y;

 wire [442:0] t;
  assign t[0] = t[1] ? t[2] : t[142];
  assign t[100] = t[114] ^ t[115];
  assign t[101] = t[80] ^ t[104];
  assign t[102] = t[116] ^ t[82];
  assign t[103] = t[116] & t[80];
  assign t[104] = t[111] & t[116];
  assign t[105] = t[82] & t[111];
  assign t[106] = t[178] ^ t[179];
  assign t[107] = t[180] ^ t[181];
  assign t[108] = t[26] ? t[182] : t[117];
  assign t[109] = t[118] ^ t[119];
  assign t[10] = t[144] & t[16];
  assign t[110] = t[61] ^ t[120];
  assign t[111] = t[121] ^ t[122];
  assign t[112] = t[123] ^ t[124];
  assign t[113] = t[125] ^ t[126];
  assign t[114] = t[125] & t[126];
  assign t[115] = t[61] & t[127];
  assign t[116] = t[128] ^ t[122];
  assign t[117] = t[183] ^ t[184];
  assign t[118] = t[110] & t[78];
  assign t[119] = t[62] & t[60];
  assign t[11] = ~(t[17]);
  assign t[120] = t[93] ^ t[129];
  assign t[121] = t[130] ^ t[131];
  assign t[122] = t[132] ^ t[115];
  assign t[123] = t[120] & t[68];
  assign t[124] = t[133] & t[66];
  assign t[125] = t[76] ^ t[58];
  assign t[126] = t[66] ^ t[93];
  assign t[127] = t[74] ^ t[134];
  assign t[128] = t[135] ^ t[136];
  assign t[129] = t[57] ^ t[68];
  assign t[12] = ~(t[144]);
  assign t[130] = t[137] ^ t[119];
  assign t[131] = t[79] & t[92];
  assign t[132] = t[48] & t[138];
  assign t[133] = t[62] ^ t[48];
  assign t[134] = t[108] ^ t[58];
  assign t[135] = t[139] ^ t[124];
  assign t[136] = t[140] & t[141];
  assign t[137] = t[62] ^ t[60];
  assign t[138] = t[61] ^ t[75];
  assign t[139] = t[66] ^ t[134];
  assign t[13] = ~(t[18]);
  assign t[140] = t[125] ^ t[79];
  assign t[141] = t[68] ^ t[66];
  assign t[142] = (t[185]);
  assign t[143] = (t[186]);
  assign t[144] = (t[187]);
  assign t[145] = (t[188]);
  assign t[146] = (t[189]);
  assign t[147] = (t[190]);
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[22] ? t[145] : t[23];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[24];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[144] & t[25]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = (t[225]);
  assign t[183] = (t[226]);
  assign t[184] = (t[227]);
  assign t[185] = t[228] ^ x[2];
  assign t[186] = t[229] ^ x[5];
  assign t[187] = t[230] ^ x[9];
  assign t[188] = t[231] ^ x[12];
  assign t[189] = t[232] ^ x[15];
  assign t[18] = ~(t[26]);
  assign t[190] = t[233] ^ x[18];
  assign t[191] = t[234] ^ x[21];
  assign t[192] = t[235] ^ x[24];
  assign t[193] = t[236] ^ x[27];
  assign t[194] = t[237] ^ x[30];
  assign t[195] = t[238] ^ x[33];
  assign t[196] = t[239] ^ x[36];
  assign t[197] = t[240] ^ x[39];
  assign t[198] = t[241] ^ x[42];
  assign t[199] = t[242] ^ x[45];
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[48];
  assign t[201] = t[244] ^ x[51];
  assign t[202] = t[245] ^ x[54];
  assign t[203] = t[246] ^ x[57];
  assign t[204] = t[247] ^ x[60];
  assign t[205] = t[248] ^ x[63];
  assign t[206] = t[249] ^ x[66];
  assign t[207] = t[250] ^ x[69];
  assign t[208] = t[251] ^ x[72];
  assign t[209] = t[252] ^ x[75];
  assign t[20] = ~(t[29] ^ t[30]);
  assign t[210] = t[253] ^ x[78];
  assign t[211] = t[254] ^ x[81];
  assign t[212] = t[255] ^ x[84];
  assign t[213] = t[256] ^ x[87];
  assign t[214] = t[257] ^ x[90];
  assign t[215] = t[258] ^ x[93];
  assign t[216] = t[259] ^ x[96];
  assign t[217] = t[260] ^ x[99];
  assign t[218] = t[261] ^ x[102];
  assign t[219] = t[262] ^ x[105];
  assign t[21] = t[146] ^ t[147];
  assign t[220] = t[263] ^ x[108];
  assign t[221] = t[264] ^ x[111];
  assign t[222] = t[265] ^ x[114];
  assign t[223] = t[266] ^ x[117];
  assign t[224] = t[267] ^ x[120];
  assign t[225] = t[268] ^ x[123];
  assign t[226] = t[269] ^ x[126];
  assign t[227] = t[270] ^ x[129];
  assign t[228] = (t[271] & ~t[272]);
  assign t[229] = (t[273] & ~t[274]);
  assign t[22] = ~(t[31]);
  assign t[230] = (t[275] & ~t[276]);
  assign t[231] = (t[277] & ~t[278]);
  assign t[232] = (t[279] & ~t[280]);
  assign t[233] = (t[281] & ~t[282]);
  assign t[234] = (t[283] & ~t[284]);
  assign t[235] = (t[285] & ~t[286]);
  assign t[236] = (t[287] & ~t[288]);
  assign t[237] = (t[289] & ~t[290]);
  assign t[238] = (t[291] & ~t[292]);
  assign t[239] = (t[293] & ~t[294]);
  assign t[23] = ~(t[32] ^ t[33]);
  assign t[240] = (t[295] & ~t[296]);
  assign t[241] = (t[297] & ~t[298]);
  assign t[242] = (t[299] & ~t[300]);
  assign t[243] = (t[301] & ~t[302]);
  assign t[244] = (t[303] & ~t[304]);
  assign t[245] = (t[305] & ~t[306]);
  assign t[246] = (t[307] & ~t[308]);
  assign t[247] = (t[309] & ~t[310]);
  assign t[248] = (t[311] & ~t[312]);
  assign t[249] = (t[313] & ~t[314]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[250] = (t[315] & ~t[316]);
  assign t[251] = (t[317] & ~t[318]);
  assign t[252] = (t[319] & ~t[320]);
  assign t[253] = (t[321] & ~t[322]);
  assign t[254] = (t[323] & ~t[324]);
  assign t[255] = (t[325] & ~t[326]);
  assign t[256] = (t[327] & ~t[328]);
  assign t[257] = (t[329] & ~t[330]);
  assign t[258] = (t[331] & ~t[332]);
  assign t[259] = (t[333] & ~t[334]);
  assign t[25] = ~(t[148] | t[36]);
  assign t[260] = (t[335] & ~t[336]);
  assign t[261] = (t[337] & ~t[338]);
  assign t[262] = (t[339] & ~t[340]);
  assign t[263] = (t[341] & ~t[342]);
  assign t[264] = (t[343] & ~t[344]);
  assign t[265] = (t[345] & ~t[346]);
  assign t[266] = (t[347] & ~t[348]);
  assign t[267] = (t[349] & ~t[350]);
  assign t[268] = (t[351] & ~t[352]);
  assign t[269] = (t[353] & ~t[354]);
  assign t[26] = ~(t[37] | t[38]);
  assign t[270] = (t[355] & ~t[356]);
  assign t[271] = t[357] ^ x[2];
  assign t[272] = t[358] ^ x[1];
  assign t[273] = t[359] ^ x[5];
  assign t[274] = t[360] ^ x[4];
  assign t[275] = t[361] ^ x[9];
  assign t[276] = t[362] ^ x[8];
  assign t[277] = t[363] ^ x[12];
  assign t[278] = t[364] ^ x[11];
  assign t[279] = t[365] ^ x[15];
  assign t[27] = ~(t[149] & t[150]);
  assign t[280] = t[366] ^ x[14];
  assign t[281] = t[367] ^ x[18];
  assign t[282] = t[368] ^ x[17];
  assign t[283] = t[369] ^ x[21];
  assign t[284] = t[370] ^ x[20];
  assign t[285] = t[371] ^ x[24];
  assign t[286] = t[372] ^ x[23];
  assign t[287] = t[373] ^ x[27];
  assign t[288] = t[374] ^ x[26];
  assign t[289] = t[375] ^ x[30];
  assign t[28] = ~(t[151] & t[152]);
  assign t[290] = t[376] ^ x[29];
  assign t[291] = t[377] ^ x[33];
  assign t[292] = t[378] ^ x[32];
  assign t[293] = t[379] ^ x[36];
  assign t[294] = t[380] ^ x[35];
  assign t[295] = t[381] ^ x[39];
  assign t[296] = t[382] ^ x[38];
  assign t[297] = t[383] ^ x[42];
  assign t[298] = t[384] ^ x[41];
  assign t[299] = t[385] ^ x[45];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[143] : t[5];
  assign t[300] = t[386] ^ x[44];
  assign t[301] = t[387] ^ x[48];
  assign t[302] = t[388] ^ x[47];
  assign t[303] = t[389] ^ x[51];
  assign t[304] = t[390] ^ x[50];
  assign t[305] = t[391] ^ x[54];
  assign t[306] = t[392] ^ x[53];
  assign t[307] = t[393] ^ x[57];
  assign t[308] = t[394] ^ x[56];
  assign t[309] = t[395] ^ x[60];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[396] ^ x[59];
  assign t[311] = t[397] ^ x[63];
  assign t[312] = t[398] ^ x[62];
  assign t[313] = t[399] ^ x[66];
  assign t[314] = t[400] ^ x[65];
  assign t[315] = t[401] ^ x[69];
  assign t[316] = t[402] ^ x[68];
  assign t[317] = t[403] ^ x[72];
  assign t[318] = t[404] ^ x[71];
  assign t[319] = t[405] ^ x[75];
  assign t[31] = ~(t[19]);
  assign t[320] = t[406] ^ x[74];
  assign t[321] = t[407] ^ x[78];
  assign t[322] = t[408] ^ x[77];
  assign t[323] = t[409] ^ x[81];
  assign t[324] = t[410] ^ x[80];
  assign t[325] = t[411] ^ x[84];
  assign t[326] = t[412] ^ x[83];
  assign t[327] = t[413] ^ x[87];
  assign t[328] = t[414] ^ x[86];
  assign t[329] = t[415] ^ x[90];
  assign t[32] = t[153] ^ t[43];
  assign t[330] = t[416] ^ x[89];
  assign t[331] = t[417] ^ x[93];
  assign t[332] = t[418] ^ x[92];
  assign t[333] = t[419] ^ x[96];
  assign t[334] = t[420] ^ x[95];
  assign t[335] = t[421] ^ x[99];
  assign t[336] = t[422] ^ x[98];
  assign t[337] = t[423] ^ x[102];
  assign t[338] = t[424] ^ x[101];
  assign t[339] = t[425] ^ x[105];
  assign t[33] = ~(t[154] ^ t[155]);
  assign t[340] = t[426] ^ x[104];
  assign t[341] = t[427] ^ x[108];
  assign t[342] = t[428] ^ x[107];
  assign t[343] = t[429] ^ x[111];
  assign t[344] = t[430] ^ x[110];
  assign t[345] = t[431] ^ x[114];
  assign t[346] = t[432] ^ x[113];
  assign t[347] = t[433] ^ x[117];
  assign t[348] = t[434] ^ x[116];
  assign t[349] = t[435] ^ x[120];
  assign t[34] = ~(t[25]);
  assign t[350] = t[436] ^ x[119];
  assign t[351] = t[437] ^ x[123];
  assign t[352] = t[438] ^ x[122];
  assign t[353] = t[439] ^ x[126];
  assign t[354] = t[440] ^ x[125];
  assign t[355] = t[441] ^ x[129];
  assign t[356] = t[442] ^ x[128];
  assign t[357] = (x[0]);
  assign t[358] = (x[0]);
  assign t[359] = (x[3]);
  assign t[35] = ~(t[156] & t[44]);
  assign t[360] = (x[3]);
  assign t[361] = (x[7]);
  assign t[362] = (x[7]);
  assign t[363] = (x[10]);
  assign t[364] = (x[10]);
  assign t[365] = (x[13]);
  assign t[366] = (x[13]);
  assign t[367] = (x[16]);
  assign t[368] = (x[16]);
  assign t[369] = (x[19]);
  assign t[36] = ~(t[45] & t[46]);
  assign t[370] = (x[19]);
  assign t[371] = (x[22]);
  assign t[372] = (x[22]);
  assign t[373] = (x[25]);
  assign t[374] = (x[25]);
  assign t[375] = (x[28]);
  assign t[376] = (x[28]);
  assign t[377] = (x[31]);
  assign t[378] = (x[31]);
  assign t[379] = (x[34]);
  assign t[37] = ~(t[157]);
  assign t[380] = (x[34]);
  assign t[381] = (x[37]);
  assign t[382] = (x[37]);
  assign t[383] = (x[40]);
  assign t[384] = (x[40]);
  assign t[385] = (x[43]);
  assign t[386] = (x[43]);
  assign t[387] = (x[46]);
  assign t[388] = (x[46]);
  assign t[389] = (x[49]);
  assign t[38] = ~(t[144]);
  assign t[390] = (x[49]);
  assign t[391] = (x[52]);
  assign t[392] = (x[52]);
  assign t[393] = (x[55]);
  assign t[394] = (x[55]);
  assign t[395] = (x[58]);
  assign t[396] = (x[58]);
  assign t[397] = (x[61]);
  assign t[398] = (x[61]);
  assign t[399] = (x[64]);
  assign t[39] = t[47] & t[48];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[64]);
  assign t[401] = (x[67]);
  assign t[402] = (x[67]);
  assign t[403] = (x[70]);
  assign t[404] = (x[70]);
  assign t[405] = (x[73]);
  assign t[406] = (x[73]);
  assign t[407] = (x[76]);
  assign t[408] = (x[76]);
  assign t[409] = (x[79]);
  assign t[40] = t[49] ^ t[50];
  assign t[410] = (x[79]);
  assign t[411] = (x[82]);
  assign t[412] = (x[82]);
  assign t[413] = (x[85]);
  assign t[414] = (x[85]);
  assign t[415] = (x[88]);
  assign t[416] = (x[88]);
  assign t[417] = (x[91]);
  assign t[418] = (x[91]);
  assign t[419] = (x[94]);
  assign t[41] = t[51] ^ t[52];
  assign t[420] = (x[94]);
  assign t[421] = (x[97]);
  assign t[422] = (x[97]);
  assign t[423] = (x[100]);
  assign t[424] = (x[100]);
  assign t[425] = (x[103]);
  assign t[426] = (x[103]);
  assign t[427] = (x[106]);
  assign t[428] = (x[106]);
  assign t[429] = (x[109]);
  assign t[42] = t[53] ^ t[54];
  assign t[430] = (x[109]);
  assign t[431] = (x[112]);
  assign t[432] = (x[112]);
  assign t[433] = (x[115]);
  assign t[434] = (x[115]);
  assign t[435] = (x[118]);
  assign t[436] = (x[118]);
  assign t[437] = (x[121]);
  assign t[438] = (x[121]);
  assign t[439] = (x[124]);
  assign t[43] = t[146] ^ t[158];
  assign t[440] = (x[124]);
  assign t[441] = (x[127]);
  assign t[442] = (x[127]);
  assign t[44] = ~(t[159]);
  assign t[45] = ~(t[160] | t[161]);
  assign t[46] = ~(t[162] | t[163]);
  assign t[47] = t[55] ^ t[56];
  assign t[48] = t[57] ^ t[58];
  assign t[49] = t[59] & t[60];
  assign t[4] = ~(t[7]);
  assign t[50] = t[55] & t[61];
  assign t[51] = t[59] & t[62];
  assign t[52] = t[63] ^ t[64];
  assign t[53] = t[65] & t[66];
  assign t[54] = t[67] & t[68];
  assign t[55] = t[69] ^ t[67];
  assign t[56] = t[70] ^ t[71];
  assign t[57] = t[26] ? t[164] : t[72];
  assign t[58] = t[26] ? t[165] : t[73];
  assign t[59] = t[69] ^ t[70];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[74] ^ t[75];
  assign t[61] = t[76] ^ t[57];
  assign t[62] = t[76] ^ t[77];
  assign t[63] = t[69] & t[78];
  assign t[64] = t[70] & t[79];
  assign t[65] = t[67] ^ t[71];
  assign t[66] = t[61] ^ t[74];
  assign t[67] = t[80] ^ t[81];
  assign t[68] = t[26] ? t[166] : t[21];
  assign t[69] = t[82] ^ t[83];
  assign t[6] = ~(t[10]);
  assign t[70] = t[84] ^ t[85];
  assign t[71] = t[86] ^ t[87];
  assign t[72] = t[167] ^ t[168];
  assign t[73] = t[169] ^ t[170];
  assign t[74] = t[88] ^ t[77];
  assign t[75] = t[89] ^ t[58];
  assign t[76] = t[26] ? t[171] : t[90];
  assign t[77] = t[26] ? t[172] : t[91];
  assign t[78] = t[92] ^ t[60];
  assign t[79] = t[93] ^ t[94];
  assign t[7] = ~(t[11]);
  assign t[80] = t[95] ^ t[96];
  assign t[81] = t[97] & t[98];
  assign t[82] = t[99] ^ t[100];
  assign t[83] = t[101] & t[102];
  assign t[84] = t[102] & t[103];
  assign t[85] = t[102] ^ t[104];
  assign t[86] = t[98] & t[105];
  assign t[87] = t[98] ^ t[104];
  assign t[88] = t[26] ? t[173] : t[106];
  assign t[89] = t[26] ? t[174] : t[107];
  assign t[8] = ~(t[12]);
  assign t[90] = t[158] ^ t[175];
  assign t[91] = t[176] ^ t[177];
  assign t[92] = t[68] ^ t[93];
  assign t[93] = t[108] ^ t[89];
  assign t[94] = t[77] ^ t[68];
  assign t[95] = t[109] ^ t[100];
  assign t[96] = t[110] ^ t[78];
  assign t[97] = t[82] ^ t[104];
  assign t[98] = t[111] ^ t[80];
  assign t[99] = t[112] ^ t[113];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind537(x, y);
 input [129:0] x;
 output y;

 wire [442:0] t;
  assign t[0] = t[1] ? t[2] : t[142];
  assign t[100] = t[114] ^ t[115];
  assign t[101] = t[80] ^ t[104];
  assign t[102] = t[116] ^ t[82];
  assign t[103] = t[116] & t[80];
  assign t[104] = t[111] & t[116];
  assign t[105] = t[82] & t[111];
  assign t[106] = t[178] ^ t[179];
  assign t[107] = t[180] ^ t[181];
  assign t[108] = t[26] ? t[182] : t[117];
  assign t[109] = t[118] ^ t[119];
  assign t[10] = t[144] & t[16];
  assign t[110] = t[61] ^ t[120];
  assign t[111] = t[121] ^ t[122];
  assign t[112] = t[123] ^ t[124];
  assign t[113] = t[125] ^ t[126];
  assign t[114] = t[125] & t[126];
  assign t[115] = t[61] & t[127];
  assign t[116] = t[128] ^ t[122];
  assign t[117] = t[183] ^ t[184];
  assign t[118] = t[110] & t[78];
  assign t[119] = t[62] & t[60];
  assign t[11] = ~(t[17]);
  assign t[120] = t[93] ^ t[129];
  assign t[121] = t[130] ^ t[131];
  assign t[122] = t[132] ^ t[115];
  assign t[123] = t[120] & t[68];
  assign t[124] = t[133] & t[66];
  assign t[125] = t[76] ^ t[58];
  assign t[126] = t[66] ^ t[93];
  assign t[127] = t[74] ^ t[134];
  assign t[128] = t[135] ^ t[136];
  assign t[129] = t[57] ^ t[68];
  assign t[12] = ~(t[144]);
  assign t[130] = t[137] ^ t[119];
  assign t[131] = t[79] & t[92];
  assign t[132] = t[48] & t[138];
  assign t[133] = t[62] ^ t[48];
  assign t[134] = t[108] ^ t[58];
  assign t[135] = t[139] ^ t[124];
  assign t[136] = t[140] & t[141];
  assign t[137] = t[62] ^ t[60];
  assign t[138] = t[61] ^ t[75];
  assign t[139] = t[66] ^ t[134];
  assign t[13] = ~(t[18]);
  assign t[140] = t[125] ^ t[79];
  assign t[141] = t[68] ^ t[66];
  assign t[142] = (t[185]);
  assign t[143] = (t[186]);
  assign t[144] = (t[187]);
  assign t[145] = (t[188]);
  assign t[146] = (t[189]);
  assign t[147] = (t[190]);
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[22] ? t[145] : t[23];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[24];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[144] & t[25]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = (t[225]);
  assign t[183] = (t[226]);
  assign t[184] = (t[227]);
  assign t[185] = t[228] ^ x[2];
  assign t[186] = t[229] ^ x[5];
  assign t[187] = t[230] ^ x[9];
  assign t[188] = t[231] ^ x[12];
  assign t[189] = t[232] ^ x[15];
  assign t[18] = ~(t[26]);
  assign t[190] = t[233] ^ x[18];
  assign t[191] = t[234] ^ x[21];
  assign t[192] = t[235] ^ x[24];
  assign t[193] = t[236] ^ x[27];
  assign t[194] = t[237] ^ x[30];
  assign t[195] = t[238] ^ x[33];
  assign t[196] = t[239] ^ x[36];
  assign t[197] = t[240] ^ x[39];
  assign t[198] = t[241] ^ x[42];
  assign t[199] = t[242] ^ x[45];
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[48];
  assign t[201] = t[244] ^ x[51];
  assign t[202] = t[245] ^ x[54];
  assign t[203] = t[246] ^ x[57];
  assign t[204] = t[247] ^ x[60];
  assign t[205] = t[248] ^ x[63];
  assign t[206] = t[249] ^ x[66];
  assign t[207] = t[250] ^ x[69];
  assign t[208] = t[251] ^ x[72];
  assign t[209] = t[252] ^ x[75];
  assign t[20] = ~(t[29] ^ t[30]);
  assign t[210] = t[253] ^ x[78];
  assign t[211] = t[254] ^ x[81];
  assign t[212] = t[255] ^ x[84];
  assign t[213] = t[256] ^ x[87];
  assign t[214] = t[257] ^ x[90];
  assign t[215] = t[258] ^ x[93];
  assign t[216] = t[259] ^ x[96];
  assign t[217] = t[260] ^ x[99];
  assign t[218] = t[261] ^ x[102];
  assign t[219] = t[262] ^ x[105];
  assign t[21] = t[146] ^ t[147];
  assign t[220] = t[263] ^ x[108];
  assign t[221] = t[264] ^ x[111];
  assign t[222] = t[265] ^ x[114];
  assign t[223] = t[266] ^ x[117];
  assign t[224] = t[267] ^ x[120];
  assign t[225] = t[268] ^ x[123];
  assign t[226] = t[269] ^ x[126];
  assign t[227] = t[270] ^ x[129];
  assign t[228] = (t[271] & ~t[272]);
  assign t[229] = (t[273] & ~t[274]);
  assign t[22] = ~(t[31]);
  assign t[230] = (t[275] & ~t[276]);
  assign t[231] = (t[277] & ~t[278]);
  assign t[232] = (t[279] & ~t[280]);
  assign t[233] = (t[281] & ~t[282]);
  assign t[234] = (t[283] & ~t[284]);
  assign t[235] = (t[285] & ~t[286]);
  assign t[236] = (t[287] & ~t[288]);
  assign t[237] = (t[289] & ~t[290]);
  assign t[238] = (t[291] & ~t[292]);
  assign t[239] = (t[293] & ~t[294]);
  assign t[23] = ~(t[32] ^ t[33]);
  assign t[240] = (t[295] & ~t[296]);
  assign t[241] = (t[297] & ~t[298]);
  assign t[242] = (t[299] & ~t[300]);
  assign t[243] = (t[301] & ~t[302]);
  assign t[244] = (t[303] & ~t[304]);
  assign t[245] = (t[305] & ~t[306]);
  assign t[246] = (t[307] & ~t[308]);
  assign t[247] = (t[309] & ~t[310]);
  assign t[248] = (t[311] & ~t[312]);
  assign t[249] = (t[313] & ~t[314]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[250] = (t[315] & ~t[316]);
  assign t[251] = (t[317] & ~t[318]);
  assign t[252] = (t[319] & ~t[320]);
  assign t[253] = (t[321] & ~t[322]);
  assign t[254] = (t[323] & ~t[324]);
  assign t[255] = (t[325] & ~t[326]);
  assign t[256] = (t[327] & ~t[328]);
  assign t[257] = (t[329] & ~t[330]);
  assign t[258] = (t[331] & ~t[332]);
  assign t[259] = (t[333] & ~t[334]);
  assign t[25] = ~(t[148] | t[36]);
  assign t[260] = (t[335] & ~t[336]);
  assign t[261] = (t[337] & ~t[338]);
  assign t[262] = (t[339] & ~t[340]);
  assign t[263] = (t[341] & ~t[342]);
  assign t[264] = (t[343] & ~t[344]);
  assign t[265] = (t[345] & ~t[346]);
  assign t[266] = (t[347] & ~t[348]);
  assign t[267] = (t[349] & ~t[350]);
  assign t[268] = (t[351] & ~t[352]);
  assign t[269] = (t[353] & ~t[354]);
  assign t[26] = ~(t[37] | t[38]);
  assign t[270] = (t[355] & ~t[356]);
  assign t[271] = t[357] ^ x[2];
  assign t[272] = t[358] ^ x[1];
  assign t[273] = t[359] ^ x[5];
  assign t[274] = t[360] ^ x[4];
  assign t[275] = t[361] ^ x[9];
  assign t[276] = t[362] ^ x[8];
  assign t[277] = t[363] ^ x[12];
  assign t[278] = t[364] ^ x[11];
  assign t[279] = t[365] ^ x[15];
  assign t[27] = ~(t[149] & t[150]);
  assign t[280] = t[366] ^ x[14];
  assign t[281] = t[367] ^ x[18];
  assign t[282] = t[368] ^ x[17];
  assign t[283] = t[369] ^ x[21];
  assign t[284] = t[370] ^ x[20];
  assign t[285] = t[371] ^ x[24];
  assign t[286] = t[372] ^ x[23];
  assign t[287] = t[373] ^ x[27];
  assign t[288] = t[374] ^ x[26];
  assign t[289] = t[375] ^ x[30];
  assign t[28] = ~(t[151] & t[152]);
  assign t[290] = t[376] ^ x[29];
  assign t[291] = t[377] ^ x[33];
  assign t[292] = t[378] ^ x[32];
  assign t[293] = t[379] ^ x[36];
  assign t[294] = t[380] ^ x[35];
  assign t[295] = t[381] ^ x[39];
  assign t[296] = t[382] ^ x[38];
  assign t[297] = t[383] ^ x[42];
  assign t[298] = t[384] ^ x[41];
  assign t[299] = t[385] ^ x[45];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[143] : t[5];
  assign t[300] = t[386] ^ x[44];
  assign t[301] = t[387] ^ x[48];
  assign t[302] = t[388] ^ x[47];
  assign t[303] = t[389] ^ x[51];
  assign t[304] = t[390] ^ x[50];
  assign t[305] = t[391] ^ x[54];
  assign t[306] = t[392] ^ x[53];
  assign t[307] = t[393] ^ x[57];
  assign t[308] = t[394] ^ x[56];
  assign t[309] = t[395] ^ x[60];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[396] ^ x[59];
  assign t[311] = t[397] ^ x[63];
  assign t[312] = t[398] ^ x[62];
  assign t[313] = t[399] ^ x[66];
  assign t[314] = t[400] ^ x[65];
  assign t[315] = t[401] ^ x[69];
  assign t[316] = t[402] ^ x[68];
  assign t[317] = t[403] ^ x[72];
  assign t[318] = t[404] ^ x[71];
  assign t[319] = t[405] ^ x[75];
  assign t[31] = ~(t[19]);
  assign t[320] = t[406] ^ x[74];
  assign t[321] = t[407] ^ x[78];
  assign t[322] = t[408] ^ x[77];
  assign t[323] = t[409] ^ x[81];
  assign t[324] = t[410] ^ x[80];
  assign t[325] = t[411] ^ x[84];
  assign t[326] = t[412] ^ x[83];
  assign t[327] = t[413] ^ x[87];
  assign t[328] = t[414] ^ x[86];
  assign t[329] = t[415] ^ x[90];
  assign t[32] = t[153] ^ t[43];
  assign t[330] = t[416] ^ x[89];
  assign t[331] = t[417] ^ x[93];
  assign t[332] = t[418] ^ x[92];
  assign t[333] = t[419] ^ x[96];
  assign t[334] = t[420] ^ x[95];
  assign t[335] = t[421] ^ x[99];
  assign t[336] = t[422] ^ x[98];
  assign t[337] = t[423] ^ x[102];
  assign t[338] = t[424] ^ x[101];
  assign t[339] = t[425] ^ x[105];
  assign t[33] = ~(t[154] ^ t[155]);
  assign t[340] = t[426] ^ x[104];
  assign t[341] = t[427] ^ x[108];
  assign t[342] = t[428] ^ x[107];
  assign t[343] = t[429] ^ x[111];
  assign t[344] = t[430] ^ x[110];
  assign t[345] = t[431] ^ x[114];
  assign t[346] = t[432] ^ x[113];
  assign t[347] = t[433] ^ x[117];
  assign t[348] = t[434] ^ x[116];
  assign t[349] = t[435] ^ x[120];
  assign t[34] = ~(t[25]);
  assign t[350] = t[436] ^ x[119];
  assign t[351] = t[437] ^ x[123];
  assign t[352] = t[438] ^ x[122];
  assign t[353] = t[439] ^ x[126];
  assign t[354] = t[440] ^ x[125];
  assign t[355] = t[441] ^ x[129];
  assign t[356] = t[442] ^ x[128];
  assign t[357] = (x[0]);
  assign t[358] = (x[0]);
  assign t[359] = (x[3]);
  assign t[35] = ~(t[156] & t[44]);
  assign t[360] = (x[3]);
  assign t[361] = (x[7]);
  assign t[362] = (x[7]);
  assign t[363] = (x[10]);
  assign t[364] = (x[10]);
  assign t[365] = (x[13]);
  assign t[366] = (x[13]);
  assign t[367] = (x[16]);
  assign t[368] = (x[16]);
  assign t[369] = (x[19]);
  assign t[36] = ~(t[45] & t[46]);
  assign t[370] = (x[19]);
  assign t[371] = (x[22]);
  assign t[372] = (x[22]);
  assign t[373] = (x[25]);
  assign t[374] = (x[25]);
  assign t[375] = (x[28]);
  assign t[376] = (x[28]);
  assign t[377] = (x[31]);
  assign t[378] = (x[31]);
  assign t[379] = (x[34]);
  assign t[37] = ~(t[157]);
  assign t[380] = (x[34]);
  assign t[381] = (x[37]);
  assign t[382] = (x[37]);
  assign t[383] = (x[40]);
  assign t[384] = (x[40]);
  assign t[385] = (x[43]);
  assign t[386] = (x[43]);
  assign t[387] = (x[46]);
  assign t[388] = (x[46]);
  assign t[389] = (x[49]);
  assign t[38] = ~(t[144]);
  assign t[390] = (x[49]);
  assign t[391] = (x[52]);
  assign t[392] = (x[52]);
  assign t[393] = (x[55]);
  assign t[394] = (x[55]);
  assign t[395] = (x[58]);
  assign t[396] = (x[58]);
  assign t[397] = (x[61]);
  assign t[398] = (x[61]);
  assign t[399] = (x[64]);
  assign t[39] = t[47] & t[48];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[64]);
  assign t[401] = (x[67]);
  assign t[402] = (x[67]);
  assign t[403] = (x[70]);
  assign t[404] = (x[70]);
  assign t[405] = (x[73]);
  assign t[406] = (x[73]);
  assign t[407] = (x[76]);
  assign t[408] = (x[76]);
  assign t[409] = (x[79]);
  assign t[40] = t[49] ^ t[50];
  assign t[410] = (x[79]);
  assign t[411] = (x[82]);
  assign t[412] = (x[82]);
  assign t[413] = (x[85]);
  assign t[414] = (x[85]);
  assign t[415] = (x[88]);
  assign t[416] = (x[88]);
  assign t[417] = (x[91]);
  assign t[418] = (x[91]);
  assign t[419] = (x[94]);
  assign t[41] = t[51] ^ t[52];
  assign t[420] = (x[94]);
  assign t[421] = (x[97]);
  assign t[422] = (x[97]);
  assign t[423] = (x[100]);
  assign t[424] = (x[100]);
  assign t[425] = (x[103]);
  assign t[426] = (x[103]);
  assign t[427] = (x[106]);
  assign t[428] = (x[106]);
  assign t[429] = (x[109]);
  assign t[42] = t[53] ^ t[54];
  assign t[430] = (x[109]);
  assign t[431] = (x[112]);
  assign t[432] = (x[112]);
  assign t[433] = (x[115]);
  assign t[434] = (x[115]);
  assign t[435] = (x[118]);
  assign t[436] = (x[118]);
  assign t[437] = (x[121]);
  assign t[438] = (x[121]);
  assign t[439] = (x[124]);
  assign t[43] = t[146] ^ t[158];
  assign t[440] = (x[124]);
  assign t[441] = (x[127]);
  assign t[442] = (x[127]);
  assign t[44] = ~(t[159]);
  assign t[45] = ~(t[160] | t[161]);
  assign t[46] = ~(t[162] | t[163]);
  assign t[47] = t[55] ^ t[56];
  assign t[48] = t[57] ^ t[58];
  assign t[49] = t[59] & t[60];
  assign t[4] = ~(t[7]);
  assign t[50] = t[55] & t[61];
  assign t[51] = t[59] & t[62];
  assign t[52] = t[63] ^ t[64];
  assign t[53] = t[65] & t[66];
  assign t[54] = t[67] & t[68];
  assign t[55] = t[69] ^ t[67];
  assign t[56] = t[70] ^ t[71];
  assign t[57] = t[26] ? t[164] : t[72];
  assign t[58] = t[26] ? t[165] : t[73];
  assign t[59] = t[69] ^ t[70];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[74] ^ t[75];
  assign t[61] = t[76] ^ t[57];
  assign t[62] = t[76] ^ t[77];
  assign t[63] = t[69] & t[78];
  assign t[64] = t[70] & t[79];
  assign t[65] = t[67] ^ t[71];
  assign t[66] = t[61] ^ t[74];
  assign t[67] = t[80] ^ t[81];
  assign t[68] = t[26] ? t[166] : t[21];
  assign t[69] = t[82] ^ t[83];
  assign t[6] = ~(t[10]);
  assign t[70] = t[84] ^ t[85];
  assign t[71] = t[86] ^ t[87];
  assign t[72] = t[167] ^ t[168];
  assign t[73] = t[169] ^ t[170];
  assign t[74] = t[88] ^ t[77];
  assign t[75] = t[89] ^ t[58];
  assign t[76] = t[26] ? t[171] : t[90];
  assign t[77] = t[26] ? t[172] : t[91];
  assign t[78] = t[92] ^ t[60];
  assign t[79] = t[93] ^ t[94];
  assign t[7] = ~(t[11]);
  assign t[80] = t[95] ^ t[96];
  assign t[81] = t[97] & t[98];
  assign t[82] = t[99] ^ t[100];
  assign t[83] = t[101] & t[102];
  assign t[84] = t[102] & t[103];
  assign t[85] = t[102] ^ t[104];
  assign t[86] = t[98] & t[105];
  assign t[87] = t[98] ^ t[104];
  assign t[88] = t[26] ? t[173] : t[106];
  assign t[89] = t[26] ? t[174] : t[107];
  assign t[8] = ~(t[12]);
  assign t[90] = t[158] ^ t[175];
  assign t[91] = t[176] ^ t[177];
  assign t[92] = t[68] ^ t[93];
  assign t[93] = t[108] ^ t[89];
  assign t[94] = t[77] ^ t[68];
  assign t[95] = t[109] ^ t[100];
  assign t[96] = t[110] ^ t[78];
  assign t[97] = t[82] ^ t[104];
  assign t[98] = t[111] ^ t[80];
  assign t[99] = t[112] ^ t[113];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind538(x, y);
 input [132:0] x;
 output y;

 wire [450:0] t;
  assign t[0] = t[1] ? t[2] : t[143];
  assign t[100] = t[115] ^ t[116];
  assign t[101] = t[117] ^ t[118];
  assign t[102] = t[91] ^ t[73];
  assign t[103] = t[119] ^ t[104];
  assign t[104] = t[26] ? t[183] : t[21];
  assign t[105] = t[62] ^ t[103];
  assign t[106] = t[120] ^ t[121];
  assign t[107] = t[122] ^ t[118];
  assign t[108] = t[123] ^ t[101];
  assign t[109] = t[124] ^ t[66];
  assign t[10] = t[145] & t[16];
  assign t[110] = t[125] ^ t[126];
  assign t[111] = t[82] ^ t[73];
  assign t[112] = t[92] ^ t[91];
  assign t[113] = t[112] & t[127];
  assign t[114] = t[112] ^ t[73];
  assign t[115] = t[128] ^ t[129];
  assign t[116] = t[130] ^ t[87];
  assign t[117] = t[130] & t[87];
  assign t[118] = t[62] & t[131];
  assign t[119] = t[26] ? t[184] : t[132];
  assign t[11] = ~(t[17]);
  assign t[120] = t[133] ^ t[129];
  assign t[121] = t[134] & t[135];
  assign t[122] = t[64] & t[68];
  assign t[123] = t[136] ^ t[137];
  assign t[124] = t[62] ^ t[138];
  assign t[125] = t[139] ^ t[137];
  assign t[126] = t[67] & t[49];
  assign t[127] = t[82] & t[92];
  assign t[128] = t[138] & t[59];
  assign t[129] = t[140] & t[105];
  assign t[12] = ~(t[145]);
  assign t[130] = t[78] ^ t[81];
  assign t[131] = t[103] ^ t[141];
  assign t[132] = t[185] ^ t[186];
  assign t[133] = t[105] ^ t[141];
  assign t[134] = t[130] ^ t[67];
  assign t[135] = t[59] ^ t[105];
  assign t[136] = t[124] & t[66];
  assign t[137] = t[89] & t[84];
  assign t[138] = t[60] ^ t[142];
  assign t[139] = t[89] ^ t[84];
  assign t[13] = ~(t[18]);
  assign t[140] = t[89] ^ t[64];
  assign t[141] = t[75] ^ t[81];
  assign t[142] = t[79] ^ t[59];
  assign t[143] = (t[187]);
  assign t[144] = (t[188]);
  assign t[145] = (t[189]);
  assign t[146] = (t[190]);
  assign t[147] = (t[191]);
  assign t[148] = (t[192]);
  assign t[149] = (t[193]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[194]);
  assign t[151] = (t[195]);
  assign t[152] = (t[196]);
  assign t[153] = (t[197]);
  assign t[154] = (t[198]);
  assign t[155] = (t[199]);
  assign t[156] = (t[200]);
  assign t[157] = (t[201]);
  assign t[158] = (t[202]);
  assign t[159] = (t[203]);
  assign t[15] = t[22] ? t[146] : t[23];
  assign t[160] = (t[204]);
  assign t[161] = (t[205]);
  assign t[162] = (t[206]);
  assign t[163] = (t[207]);
  assign t[164] = (t[208]);
  assign t[165] = (t[209]);
  assign t[166] = (t[210]);
  assign t[167] = (t[211]);
  assign t[168] = (t[212]);
  assign t[169] = (t[213]);
  assign t[16] = t[19] & t[24];
  assign t[170] = (t[214]);
  assign t[171] = (t[215]);
  assign t[172] = (t[216]);
  assign t[173] = (t[217]);
  assign t[174] = (t[218]);
  assign t[175] = (t[219]);
  assign t[176] = (t[220]);
  assign t[177] = (t[221]);
  assign t[178] = (t[222]);
  assign t[179] = (t[223]);
  assign t[17] = ~(t[145] & t[25]);
  assign t[180] = (t[224]);
  assign t[181] = (t[225]);
  assign t[182] = (t[226]);
  assign t[183] = (t[227]);
  assign t[184] = (t[228]);
  assign t[185] = (t[229]);
  assign t[186] = (t[230]);
  assign t[187] = t[231] ^ x[2];
  assign t[188] = t[232] ^ x[5];
  assign t[189] = t[233] ^ x[9];
  assign t[18] = ~(t[26]);
  assign t[190] = t[234] ^ x[12];
  assign t[191] = t[235] ^ x[15];
  assign t[192] = t[236] ^ x[18];
  assign t[193] = t[237] ^ x[21];
  assign t[194] = t[238] ^ x[24];
  assign t[195] = t[239] ^ x[27];
  assign t[196] = t[240] ^ x[30];
  assign t[197] = t[241] ^ x[33];
  assign t[198] = t[242] ^ x[36];
  assign t[199] = t[243] ^ x[39];
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[244] ^ x[42];
  assign t[201] = t[245] ^ x[45];
  assign t[202] = t[246] ^ x[48];
  assign t[203] = t[247] ^ x[51];
  assign t[204] = t[248] ^ x[54];
  assign t[205] = t[249] ^ x[57];
  assign t[206] = t[250] ^ x[60];
  assign t[207] = t[251] ^ x[63];
  assign t[208] = t[252] ^ x[66];
  assign t[209] = t[253] ^ x[69];
  assign t[20] = ~(t[29] ^ t[30]);
  assign t[210] = t[254] ^ x[72];
  assign t[211] = t[255] ^ x[75];
  assign t[212] = t[256] ^ x[78];
  assign t[213] = t[257] ^ x[81];
  assign t[214] = t[258] ^ x[84];
  assign t[215] = t[259] ^ x[87];
  assign t[216] = t[260] ^ x[90];
  assign t[217] = t[261] ^ x[93];
  assign t[218] = t[262] ^ x[96];
  assign t[219] = t[263] ^ x[99];
  assign t[21] = t[147] ^ t[148];
  assign t[220] = t[264] ^ x[102];
  assign t[221] = t[265] ^ x[105];
  assign t[222] = t[266] ^ x[108];
  assign t[223] = t[267] ^ x[111];
  assign t[224] = t[268] ^ x[114];
  assign t[225] = t[269] ^ x[117];
  assign t[226] = t[270] ^ x[120];
  assign t[227] = t[271] ^ x[123];
  assign t[228] = t[272] ^ x[126];
  assign t[229] = t[273] ^ x[129];
  assign t[22] = ~(t[31]);
  assign t[230] = t[274] ^ x[132];
  assign t[231] = (t[275] & ~t[276]);
  assign t[232] = (t[277] & ~t[278]);
  assign t[233] = (t[279] & ~t[280]);
  assign t[234] = (t[281] & ~t[282]);
  assign t[235] = (t[283] & ~t[284]);
  assign t[236] = (t[285] & ~t[286]);
  assign t[237] = (t[287] & ~t[288]);
  assign t[238] = (t[289] & ~t[290]);
  assign t[239] = (t[291] & ~t[292]);
  assign t[23] = ~(t[32] ^ t[33]);
  assign t[240] = (t[293] & ~t[294]);
  assign t[241] = (t[295] & ~t[296]);
  assign t[242] = (t[297] & ~t[298]);
  assign t[243] = (t[299] & ~t[300]);
  assign t[244] = (t[301] & ~t[302]);
  assign t[245] = (t[303] & ~t[304]);
  assign t[246] = (t[305] & ~t[306]);
  assign t[247] = (t[307] & ~t[308]);
  assign t[248] = (t[309] & ~t[310]);
  assign t[249] = (t[311] & ~t[312]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[250] = (t[313] & ~t[314]);
  assign t[251] = (t[315] & ~t[316]);
  assign t[252] = (t[317] & ~t[318]);
  assign t[253] = (t[319] & ~t[320]);
  assign t[254] = (t[321] & ~t[322]);
  assign t[255] = (t[323] & ~t[324]);
  assign t[256] = (t[325] & ~t[326]);
  assign t[257] = (t[327] & ~t[328]);
  assign t[258] = (t[329] & ~t[330]);
  assign t[259] = (t[331] & ~t[332]);
  assign t[25] = ~(t[149] | t[36]);
  assign t[260] = (t[333] & ~t[334]);
  assign t[261] = (t[335] & ~t[336]);
  assign t[262] = (t[337] & ~t[338]);
  assign t[263] = (t[339] & ~t[340]);
  assign t[264] = (t[341] & ~t[342]);
  assign t[265] = (t[343] & ~t[344]);
  assign t[266] = (t[345] & ~t[346]);
  assign t[267] = (t[347] & ~t[348]);
  assign t[268] = (t[349] & ~t[350]);
  assign t[269] = (t[351] & ~t[352]);
  assign t[26] = ~(t[37] | t[38]);
  assign t[270] = (t[353] & ~t[354]);
  assign t[271] = (t[355] & ~t[356]);
  assign t[272] = (t[357] & ~t[358]);
  assign t[273] = (t[359] & ~t[360]);
  assign t[274] = (t[361] & ~t[362]);
  assign t[275] = t[363] ^ x[2];
  assign t[276] = t[364] ^ x[1];
  assign t[277] = t[365] ^ x[5];
  assign t[278] = t[366] ^ x[4];
  assign t[279] = t[367] ^ x[9];
  assign t[27] = ~(t[150] & t[151]);
  assign t[280] = t[368] ^ x[8];
  assign t[281] = t[369] ^ x[12];
  assign t[282] = t[370] ^ x[11];
  assign t[283] = t[371] ^ x[15];
  assign t[284] = t[372] ^ x[14];
  assign t[285] = t[373] ^ x[18];
  assign t[286] = t[374] ^ x[17];
  assign t[287] = t[375] ^ x[21];
  assign t[288] = t[376] ^ x[20];
  assign t[289] = t[377] ^ x[24];
  assign t[28] = ~(t[152] & t[153]);
  assign t[290] = t[378] ^ x[23];
  assign t[291] = t[379] ^ x[27];
  assign t[292] = t[380] ^ x[26];
  assign t[293] = t[381] ^ x[30];
  assign t[294] = t[382] ^ x[29];
  assign t[295] = t[383] ^ x[33];
  assign t[296] = t[384] ^ x[32];
  assign t[297] = t[385] ^ x[36];
  assign t[298] = t[386] ^ x[35];
  assign t[299] = t[387] ^ x[39];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[144] : t[5];
  assign t[300] = t[388] ^ x[38];
  assign t[301] = t[389] ^ x[42];
  assign t[302] = t[390] ^ x[41];
  assign t[303] = t[391] ^ x[45];
  assign t[304] = t[392] ^ x[44];
  assign t[305] = t[393] ^ x[48];
  assign t[306] = t[394] ^ x[47];
  assign t[307] = t[395] ^ x[51];
  assign t[308] = t[396] ^ x[50];
  assign t[309] = t[397] ^ x[54];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[398] ^ x[53];
  assign t[311] = t[399] ^ x[57];
  assign t[312] = t[400] ^ x[56];
  assign t[313] = t[401] ^ x[60];
  assign t[314] = t[402] ^ x[59];
  assign t[315] = t[403] ^ x[63];
  assign t[316] = t[404] ^ x[62];
  assign t[317] = t[405] ^ x[66];
  assign t[318] = t[406] ^ x[65];
  assign t[319] = t[407] ^ x[69];
  assign t[31] = ~(t[19]);
  assign t[320] = t[408] ^ x[68];
  assign t[321] = t[409] ^ x[72];
  assign t[322] = t[410] ^ x[71];
  assign t[323] = t[411] ^ x[75];
  assign t[324] = t[412] ^ x[74];
  assign t[325] = t[413] ^ x[78];
  assign t[326] = t[414] ^ x[77];
  assign t[327] = t[415] ^ x[81];
  assign t[328] = t[416] ^ x[80];
  assign t[329] = t[417] ^ x[84];
  assign t[32] = t[43] ^ t[44];
  assign t[330] = t[418] ^ x[83];
  assign t[331] = t[419] ^ x[87];
  assign t[332] = t[420] ^ x[86];
  assign t[333] = t[421] ^ x[90];
  assign t[334] = t[422] ^ x[89];
  assign t[335] = t[423] ^ x[93];
  assign t[336] = t[424] ^ x[92];
  assign t[337] = t[425] ^ x[96];
  assign t[338] = t[426] ^ x[95];
  assign t[339] = t[427] ^ x[99];
  assign t[33] = ~(t[154] ^ t[155]);
  assign t[340] = t[428] ^ x[98];
  assign t[341] = t[429] ^ x[102];
  assign t[342] = t[430] ^ x[101];
  assign t[343] = t[431] ^ x[105];
  assign t[344] = t[432] ^ x[104];
  assign t[345] = t[433] ^ x[108];
  assign t[346] = t[434] ^ x[107];
  assign t[347] = t[435] ^ x[111];
  assign t[348] = t[436] ^ x[110];
  assign t[349] = t[437] ^ x[114];
  assign t[34] = ~(t[25]);
  assign t[350] = t[438] ^ x[113];
  assign t[351] = t[439] ^ x[117];
  assign t[352] = t[440] ^ x[116];
  assign t[353] = t[441] ^ x[120];
  assign t[354] = t[442] ^ x[119];
  assign t[355] = t[443] ^ x[123];
  assign t[356] = t[444] ^ x[122];
  assign t[357] = t[445] ^ x[126];
  assign t[358] = t[446] ^ x[125];
  assign t[359] = t[447] ^ x[129];
  assign t[35] = ~(t[156] & t[45]);
  assign t[360] = t[448] ^ x[128];
  assign t[361] = t[449] ^ x[132];
  assign t[362] = t[450] ^ x[131];
  assign t[363] = (x[0]);
  assign t[364] = (x[0]);
  assign t[365] = (x[3]);
  assign t[366] = (x[3]);
  assign t[367] = (x[7]);
  assign t[368] = (x[7]);
  assign t[369] = (x[10]);
  assign t[36] = ~(t[46] & t[47]);
  assign t[370] = (x[10]);
  assign t[371] = (x[13]);
  assign t[372] = (x[13]);
  assign t[373] = (x[16]);
  assign t[374] = (x[16]);
  assign t[375] = (x[19]);
  assign t[376] = (x[19]);
  assign t[377] = (x[22]);
  assign t[378] = (x[22]);
  assign t[379] = (x[25]);
  assign t[37] = ~(t[157]);
  assign t[380] = (x[25]);
  assign t[381] = (x[28]);
  assign t[382] = (x[28]);
  assign t[383] = (x[31]);
  assign t[384] = (x[31]);
  assign t[385] = (x[34]);
  assign t[386] = (x[34]);
  assign t[387] = (x[37]);
  assign t[388] = (x[37]);
  assign t[389] = (x[40]);
  assign t[38] = ~(t[145]);
  assign t[390] = (x[40]);
  assign t[391] = (x[43]);
  assign t[392] = (x[43]);
  assign t[393] = (x[46]);
  assign t[394] = (x[46]);
  assign t[395] = (x[49]);
  assign t[396] = (x[49]);
  assign t[397] = (x[52]);
  assign t[398] = (x[52]);
  assign t[399] = (x[55]);
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[55]);
  assign t[401] = (x[58]);
  assign t[402] = (x[58]);
  assign t[403] = (x[61]);
  assign t[404] = (x[61]);
  assign t[405] = (x[64]);
  assign t[406] = (x[64]);
  assign t[407] = (x[67]);
  assign t[408] = (x[67]);
  assign t[409] = (x[70]);
  assign t[40] = t[50] ^ t[51];
  assign t[410] = (x[70]);
  assign t[411] = (x[73]);
  assign t[412] = (x[73]);
  assign t[413] = (x[76]);
  assign t[414] = (x[76]);
  assign t[415] = (x[79]);
  assign t[416] = (x[79]);
  assign t[417] = (x[82]);
  assign t[418] = (x[82]);
  assign t[419] = (x[85]);
  assign t[41] = t[52] ^ t[53];
  assign t[420] = (x[85]);
  assign t[421] = (x[88]);
  assign t[422] = (x[88]);
  assign t[423] = (x[91]);
  assign t[424] = (x[91]);
  assign t[425] = (x[94]);
  assign t[426] = (x[94]);
  assign t[427] = (x[97]);
  assign t[428] = (x[97]);
  assign t[429] = (x[100]);
  assign t[42] = t[54] ^ t[55];
  assign t[430] = (x[100]);
  assign t[431] = (x[103]);
  assign t[432] = (x[103]);
  assign t[433] = (x[106]);
  assign t[434] = (x[106]);
  assign t[435] = (x[109]);
  assign t[436] = (x[109]);
  assign t[437] = (x[112]);
  assign t[438] = (x[112]);
  assign t[439] = (x[115]);
  assign t[43] = t[158] ^ t[159];
  assign t[440] = (x[115]);
  assign t[441] = (x[118]);
  assign t[442] = (x[118]);
  assign t[443] = (x[121]);
  assign t[444] = (x[121]);
  assign t[445] = (x[124]);
  assign t[446] = (x[124]);
  assign t[447] = (x[127]);
  assign t[448] = (x[127]);
  assign t[449] = (x[130]);
  assign t[44] = t[147] ^ t[56];
  assign t[450] = (x[130]);
  assign t[45] = ~(t[160]);
  assign t[46] = ~(t[161] | t[162]);
  assign t[47] = ~(t[163] | t[164]);
  assign t[48] = t[57] ^ t[58];
  assign t[49] = t[59] ^ t[60];
  assign t[4] = ~(t[7]);
  assign t[50] = t[61] & t[62];
  assign t[51] = t[63] & t[64];
  assign t[52] = t[65] & t[66];
  assign t[53] = t[48] & t[67];
  assign t[54] = t[63] & t[68];
  assign t[55] = t[69] ^ t[70];
  assign t[56] = t[165] ^ t[166];
  assign t[57] = t[71] & t[72];
  assign t[58] = t[71] ^ t[73];
  assign t[59] = t[26] ? t[167] : t[74];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[75] ^ t[76];
  assign t[61] = t[65] ^ t[77];
  assign t[62] = t[78] ^ t[79];
  assign t[63] = t[61] ^ t[80];
  assign t[64] = t[79] ^ t[81];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[49] ^ t[84];
  assign t[67] = t[60] ^ t[85];
  assign t[68] = t[62] ^ t[86];
  assign t[69] = t[80] & t[87];
  assign t[6] = ~(t[10]);
  assign t[70] = t[88] & t[89];
  assign t[71] = t[90] ^ t[82];
  assign t[72] = t[90] & t[91];
  assign t[73] = t[92] & t[90];
  assign t[74] = t[166] ^ t[168];
  assign t[75] = t[26] ? t[169] : t[93];
  assign t[76] = t[26] ? t[170] : t[94];
  assign t[77] = t[91] ^ t[95];
  assign t[78] = t[26] ? t[171] : t[96];
  assign t[79] = t[26] ? t[172] : t[97];
  assign t[7] = ~(t[11]);
  assign t[80] = t[48] ^ t[98];
  assign t[81] = t[26] ? t[173] : t[99];
  assign t[82] = t[100] ^ t[101];
  assign t[83] = t[102] & t[71];
  assign t[84] = t[103] ^ t[86];
  assign t[85] = t[104] ^ t[59];
  assign t[86] = t[76] ^ t[81];
  assign t[87] = t[105] ^ t[60];
  assign t[88] = t[65] ^ t[48];
  assign t[89] = t[78] ^ t[104];
  assign t[8] = ~(t[12]);
  assign t[90] = t[106] ^ t[107];
  assign t[91] = t[108] ^ t[109];
  assign t[92] = t[110] ^ t[107];
  assign t[93] = t[174] ^ t[175];
  assign t[94] = t[176] ^ t[177];
  assign t[95] = t[111] & t[112];
  assign t[96] = t[165] ^ t[178];
  assign t[97] = t[179] ^ t[180];
  assign t[98] = t[113] ^ t[114];
  assign t[99] = t[181] ^ t[182];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind539(x, y);
 input [132:0] x;
 output y;

 wire [450:0] t;
  assign t[0] = t[1] ? t[2] : t[143];
  assign t[100] = t[115] ^ t[116];
  assign t[101] = t[117] ^ t[118];
  assign t[102] = t[91] ^ t[73];
  assign t[103] = t[119] ^ t[104];
  assign t[104] = t[26] ? t[183] : t[21];
  assign t[105] = t[62] ^ t[103];
  assign t[106] = t[120] ^ t[121];
  assign t[107] = t[122] ^ t[118];
  assign t[108] = t[123] ^ t[101];
  assign t[109] = t[124] ^ t[66];
  assign t[10] = t[145] & t[16];
  assign t[110] = t[125] ^ t[126];
  assign t[111] = t[82] ^ t[73];
  assign t[112] = t[92] ^ t[91];
  assign t[113] = t[112] & t[127];
  assign t[114] = t[112] ^ t[73];
  assign t[115] = t[128] ^ t[129];
  assign t[116] = t[130] ^ t[87];
  assign t[117] = t[130] & t[87];
  assign t[118] = t[62] & t[131];
  assign t[119] = t[26] ? t[184] : t[132];
  assign t[11] = ~(t[17]);
  assign t[120] = t[133] ^ t[129];
  assign t[121] = t[134] & t[135];
  assign t[122] = t[64] & t[68];
  assign t[123] = t[136] ^ t[137];
  assign t[124] = t[62] ^ t[138];
  assign t[125] = t[139] ^ t[137];
  assign t[126] = t[67] & t[49];
  assign t[127] = t[82] & t[92];
  assign t[128] = t[138] & t[59];
  assign t[129] = t[140] & t[105];
  assign t[12] = ~(t[145]);
  assign t[130] = t[78] ^ t[81];
  assign t[131] = t[103] ^ t[141];
  assign t[132] = t[185] ^ t[186];
  assign t[133] = t[105] ^ t[141];
  assign t[134] = t[130] ^ t[67];
  assign t[135] = t[59] ^ t[105];
  assign t[136] = t[124] & t[66];
  assign t[137] = t[89] & t[84];
  assign t[138] = t[60] ^ t[142];
  assign t[139] = t[89] ^ t[84];
  assign t[13] = ~(t[18]);
  assign t[140] = t[89] ^ t[64];
  assign t[141] = t[75] ^ t[81];
  assign t[142] = t[79] ^ t[59];
  assign t[143] = (t[187]);
  assign t[144] = (t[188]);
  assign t[145] = (t[189]);
  assign t[146] = (t[190]);
  assign t[147] = (t[191]);
  assign t[148] = (t[192]);
  assign t[149] = (t[193]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[194]);
  assign t[151] = (t[195]);
  assign t[152] = (t[196]);
  assign t[153] = (t[197]);
  assign t[154] = (t[198]);
  assign t[155] = (t[199]);
  assign t[156] = (t[200]);
  assign t[157] = (t[201]);
  assign t[158] = (t[202]);
  assign t[159] = (t[203]);
  assign t[15] = t[22] ? t[146] : t[23];
  assign t[160] = (t[204]);
  assign t[161] = (t[205]);
  assign t[162] = (t[206]);
  assign t[163] = (t[207]);
  assign t[164] = (t[208]);
  assign t[165] = (t[209]);
  assign t[166] = (t[210]);
  assign t[167] = (t[211]);
  assign t[168] = (t[212]);
  assign t[169] = (t[213]);
  assign t[16] = t[19] & t[24];
  assign t[170] = (t[214]);
  assign t[171] = (t[215]);
  assign t[172] = (t[216]);
  assign t[173] = (t[217]);
  assign t[174] = (t[218]);
  assign t[175] = (t[219]);
  assign t[176] = (t[220]);
  assign t[177] = (t[221]);
  assign t[178] = (t[222]);
  assign t[179] = (t[223]);
  assign t[17] = ~(t[145] & t[25]);
  assign t[180] = (t[224]);
  assign t[181] = (t[225]);
  assign t[182] = (t[226]);
  assign t[183] = (t[227]);
  assign t[184] = (t[228]);
  assign t[185] = (t[229]);
  assign t[186] = (t[230]);
  assign t[187] = t[231] ^ x[2];
  assign t[188] = t[232] ^ x[5];
  assign t[189] = t[233] ^ x[9];
  assign t[18] = ~(t[26]);
  assign t[190] = t[234] ^ x[12];
  assign t[191] = t[235] ^ x[15];
  assign t[192] = t[236] ^ x[18];
  assign t[193] = t[237] ^ x[21];
  assign t[194] = t[238] ^ x[24];
  assign t[195] = t[239] ^ x[27];
  assign t[196] = t[240] ^ x[30];
  assign t[197] = t[241] ^ x[33];
  assign t[198] = t[242] ^ x[36];
  assign t[199] = t[243] ^ x[39];
  assign t[19] = ~(t[27] | t[28]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[244] ^ x[42];
  assign t[201] = t[245] ^ x[45];
  assign t[202] = t[246] ^ x[48];
  assign t[203] = t[247] ^ x[51];
  assign t[204] = t[248] ^ x[54];
  assign t[205] = t[249] ^ x[57];
  assign t[206] = t[250] ^ x[60];
  assign t[207] = t[251] ^ x[63];
  assign t[208] = t[252] ^ x[66];
  assign t[209] = t[253] ^ x[69];
  assign t[20] = ~(t[29] ^ t[30]);
  assign t[210] = t[254] ^ x[72];
  assign t[211] = t[255] ^ x[75];
  assign t[212] = t[256] ^ x[78];
  assign t[213] = t[257] ^ x[81];
  assign t[214] = t[258] ^ x[84];
  assign t[215] = t[259] ^ x[87];
  assign t[216] = t[260] ^ x[90];
  assign t[217] = t[261] ^ x[93];
  assign t[218] = t[262] ^ x[96];
  assign t[219] = t[263] ^ x[99];
  assign t[21] = t[147] ^ t[148];
  assign t[220] = t[264] ^ x[102];
  assign t[221] = t[265] ^ x[105];
  assign t[222] = t[266] ^ x[108];
  assign t[223] = t[267] ^ x[111];
  assign t[224] = t[268] ^ x[114];
  assign t[225] = t[269] ^ x[117];
  assign t[226] = t[270] ^ x[120];
  assign t[227] = t[271] ^ x[123];
  assign t[228] = t[272] ^ x[126];
  assign t[229] = t[273] ^ x[129];
  assign t[22] = ~(t[31]);
  assign t[230] = t[274] ^ x[132];
  assign t[231] = (t[275] & ~t[276]);
  assign t[232] = (t[277] & ~t[278]);
  assign t[233] = (t[279] & ~t[280]);
  assign t[234] = (t[281] & ~t[282]);
  assign t[235] = (t[283] & ~t[284]);
  assign t[236] = (t[285] & ~t[286]);
  assign t[237] = (t[287] & ~t[288]);
  assign t[238] = (t[289] & ~t[290]);
  assign t[239] = (t[291] & ~t[292]);
  assign t[23] = ~(t[32] ^ t[33]);
  assign t[240] = (t[293] & ~t[294]);
  assign t[241] = (t[295] & ~t[296]);
  assign t[242] = (t[297] & ~t[298]);
  assign t[243] = (t[299] & ~t[300]);
  assign t[244] = (t[301] & ~t[302]);
  assign t[245] = (t[303] & ~t[304]);
  assign t[246] = (t[305] & ~t[306]);
  assign t[247] = (t[307] & ~t[308]);
  assign t[248] = (t[309] & ~t[310]);
  assign t[249] = (t[311] & ~t[312]);
  assign t[24] = ~(t[34] | t[35]);
  assign t[250] = (t[313] & ~t[314]);
  assign t[251] = (t[315] & ~t[316]);
  assign t[252] = (t[317] & ~t[318]);
  assign t[253] = (t[319] & ~t[320]);
  assign t[254] = (t[321] & ~t[322]);
  assign t[255] = (t[323] & ~t[324]);
  assign t[256] = (t[325] & ~t[326]);
  assign t[257] = (t[327] & ~t[328]);
  assign t[258] = (t[329] & ~t[330]);
  assign t[259] = (t[331] & ~t[332]);
  assign t[25] = ~(t[149] | t[36]);
  assign t[260] = (t[333] & ~t[334]);
  assign t[261] = (t[335] & ~t[336]);
  assign t[262] = (t[337] & ~t[338]);
  assign t[263] = (t[339] & ~t[340]);
  assign t[264] = (t[341] & ~t[342]);
  assign t[265] = (t[343] & ~t[344]);
  assign t[266] = (t[345] & ~t[346]);
  assign t[267] = (t[347] & ~t[348]);
  assign t[268] = (t[349] & ~t[350]);
  assign t[269] = (t[351] & ~t[352]);
  assign t[26] = ~(t[37] | t[38]);
  assign t[270] = (t[353] & ~t[354]);
  assign t[271] = (t[355] & ~t[356]);
  assign t[272] = (t[357] & ~t[358]);
  assign t[273] = (t[359] & ~t[360]);
  assign t[274] = (t[361] & ~t[362]);
  assign t[275] = t[363] ^ x[2];
  assign t[276] = t[364] ^ x[1];
  assign t[277] = t[365] ^ x[5];
  assign t[278] = t[366] ^ x[4];
  assign t[279] = t[367] ^ x[9];
  assign t[27] = ~(t[150] & t[151]);
  assign t[280] = t[368] ^ x[8];
  assign t[281] = t[369] ^ x[12];
  assign t[282] = t[370] ^ x[11];
  assign t[283] = t[371] ^ x[15];
  assign t[284] = t[372] ^ x[14];
  assign t[285] = t[373] ^ x[18];
  assign t[286] = t[374] ^ x[17];
  assign t[287] = t[375] ^ x[21];
  assign t[288] = t[376] ^ x[20];
  assign t[289] = t[377] ^ x[24];
  assign t[28] = ~(t[152] & t[153]);
  assign t[290] = t[378] ^ x[23];
  assign t[291] = t[379] ^ x[27];
  assign t[292] = t[380] ^ x[26];
  assign t[293] = t[381] ^ x[30];
  assign t[294] = t[382] ^ x[29];
  assign t[295] = t[383] ^ x[33];
  assign t[296] = t[384] ^ x[32];
  assign t[297] = t[385] ^ x[36];
  assign t[298] = t[386] ^ x[35];
  assign t[299] = t[387] ^ x[39];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[144] : t[5];
  assign t[300] = t[388] ^ x[38];
  assign t[301] = t[389] ^ x[42];
  assign t[302] = t[390] ^ x[41];
  assign t[303] = t[391] ^ x[45];
  assign t[304] = t[392] ^ x[44];
  assign t[305] = t[393] ^ x[48];
  assign t[306] = t[394] ^ x[47];
  assign t[307] = t[395] ^ x[51];
  assign t[308] = t[396] ^ x[50];
  assign t[309] = t[397] ^ x[54];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[398] ^ x[53];
  assign t[311] = t[399] ^ x[57];
  assign t[312] = t[400] ^ x[56];
  assign t[313] = t[401] ^ x[60];
  assign t[314] = t[402] ^ x[59];
  assign t[315] = t[403] ^ x[63];
  assign t[316] = t[404] ^ x[62];
  assign t[317] = t[405] ^ x[66];
  assign t[318] = t[406] ^ x[65];
  assign t[319] = t[407] ^ x[69];
  assign t[31] = ~(t[19]);
  assign t[320] = t[408] ^ x[68];
  assign t[321] = t[409] ^ x[72];
  assign t[322] = t[410] ^ x[71];
  assign t[323] = t[411] ^ x[75];
  assign t[324] = t[412] ^ x[74];
  assign t[325] = t[413] ^ x[78];
  assign t[326] = t[414] ^ x[77];
  assign t[327] = t[415] ^ x[81];
  assign t[328] = t[416] ^ x[80];
  assign t[329] = t[417] ^ x[84];
  assign t[32] = t[43] ^ t[44];
  assign t[330] = t[418] ^ x[83];
  assign t[331] = t[419] ^ x[87];
  assign t[332] = t[420] ^ x[86];
  assign t[333] = t[421] ^ x[90];
  assign t[334] = t[422] ^ x[89];
  assign t[335] = t[423] ^ x[93];
  assign t[336] = t[424] ^ x[92];
  assign t[337] = t[425] ^ x[96];
  assign t[338] = t[426] ^ x[95];
  assign t[339] = t[427] ^ x[99];
  assign t[33] = ~(t[154] ^ t[155]);
  assign t[340] = t[428] ^ x[98];
  assign t[341] = t[429] ^ x[102];
  assign t[342] = t[430] ^ x[101];
  assign t[343] = t[431] ^ x[105];
  assign t[344] = t[432] ^ x[104];
  assign t[345] = t[433] ^ x[108];
  assign t[346] = t[434] ^ x[107];
  assign t[347] = t[435] ^ x[111];
  assign t[348] = t[436] ^ x[110];
  assign t[349] = t[437] ^ x[114];
  assign t[34] = ~(t[25]);
  assign t[350] = t[438] ^ x[113];
  assign t[351] = t[439] ^ x[117];
  assign t[352] = t[440] ^ x[116];
  assign t[353] = t[441] ^ x[120];
  assign t[354] = t[442] ^ x[119];
  assign t[355] = t[443] ^ x[123];
  assign t[356] = t[444] ^ x[122];
  assign t[357] = t[445] ^ x[126];
  assign t[358] = t[446] ^ x[125];
  assign t[359] = t[447] ^ x[129];
  assign t[35] = ~(t[156] & t[45]);
  assign t[360] = t[448] ^ x[128];
  assign t[361] = t[449] ^ x[132];
  assign t[362] = t[450] ^ x[131];
  assign t[363] = (x[0]);
  assign t[364] = (x[0]);
  assign t[365] = (x[3]);
  assign t[366] = (x[3]);
  assign t[367] = (x[7]);
  assign t[368] = (x[7]);
  assign t[369] = (x[10]);
  assign t[36] = ~(t[46] & t[47]);
  assign t[370] = (x[10]);
  assign t[371] = (x[13]);
  assign t[372] = (x[13]);
  assign t[373] = (x[16]);
  assign t[374] = (x[16]);
  assign t[375] = (x[19]);
  assign t[376] = (x[19]);
  assign t[377] = (x[22]);
  assign t[378] = (x[22]);
  assign t[379] = (x[25]);
  assign t[37] = ~(t[157]);
  assign t[380] = (x[25]);
  assign t[381] = (x[28]);
  assign t[382] = (x[28]);
  assign t[383] = (x[31]);
  assign t[384] = (x[31]);
  assign t[385] = (x[34]);
  assign t[386] = (x[34]);
  assign t[387] = (x[37]);
  assign t[388] = (x[37]);
  assign t[389] = (x[40]);
  assign t[38] = ~(t[145]);
  assign t[390] = (x[40]);
  assign t[391] = (x[43]);
  assign t[392] = (x[43]);
  assign t[393] = (x[46]);
  assign t[394] = (x[46]);
  assign t[395] = (x[49]);
  assign t[396] = (x[49]);
  assign t[397] = (x[52]);
  assign t[398] = (x[52]);
  assign t[399] = (x[55]);
  assign t[39] = t[48] & t[49];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[55]);
  assign t[401] = (x[58]);
  assign t[402] = (x[58]);
  assign t[403] = (x[61]);
  assign t[404] = (x[61]);
  assign t[405] = (x[64]);
  assign t[406] = (x[64]);
  assign t[407] = (x[67]);
  assign t[408] = (x[67]);
  assign t[409] = (x[70]);
  assign t[40] = t[50] ^ t[51];
  assign t[410] = (x[70]);
  assign t[411] = (x[73]);
  assign t[412] = (x[73]);
  assign t[413] = (x[76]);
  assign t[414] = (x[76]);
  assign t[415] = (x[79]);
  assign t[416] = (x[79]);
  assign t[417] = (x[82]);
  assign t[418] = (x[82]);
  assign t[419] = (x[85]);
  assign t[41] = t[52] ^ t[53];
  assign t[420] = (x[85]);
  assign t[421] = (x[88]);
  assign t[422] = (x[88]);
  assign t[423] = (x[91]);
  assign t[424] = (x[91]);
  assign t[425] = (x[94]);
  assign t[426] = (x[94]);
  assign t[427] = (x[97]);
  assign t[428] = (x[97]);
  assign t[429] = (x[100]);
  assign t[42] = t[54] ^ t[55];
  assign t[430] = (x[100]);
  assign t[431] = (x[103]);
  assign t[432] = (x[103]);
  assign t[433] = (x[106]);
  assign t[434] = (x[106]);
  assign t[435] = (x[109]);
  assign t[436] = (x[109]);
  assign t[437] = (x[112]);
  assign t[438] = (x[112]);
  assign t[439] = (x[115]);
  assign t[43] = t[158] ^ t[159];
  assign t[440] = (x[115]);
  assign t[441] = (x[118]);
  assign t[442] = (x[118]);
  assign t[443] = (x[121]);
  assign t[444] = (x[121]);
  assign t[445] = (x[124]);
  assign t[446] = (x[124]);
  assign t[447] = (x[127]);
  assign t[448] = (x[127]);
  assign t[449] = (x[130]);
  assign t[44] = t[147] ^ t[56];
  assign t[450] = (x[130]);
  assign t[45] = ~(t[160]);
  assign t[46] = ~(t[161] | t[162]);
  assign t[47] = ~(t[163] | t[164]);
  assign t[48] = t[57] ^ t[58];
  assign t[49] = t[59] ^ t[60];
  assign t[4] = ~(t[7]);
  assign t[50] = t[61] & t[62];
  assign t[51] = t[63] & t[64];
  assign t[52] = t[65] & t[66];
  assign t[53] = t[48] & t[67];
  assign t[54] = t[63] & t[68];
  assign t[55] = t[69] ^ t[70];
  assign t[56] = t[165] ^ t[166];
  assign t[57] = t[71] & t[72];
  assign t[58] = t[71] ^ t[73];
  assign t[59] = t[26] ? t[167] : t[74];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[75] ^ t[76];
  assign t[61] = t[65] ^ t[77];
  assign t[62] = t[78] ^ t[79];
  assign t[63] = t[61] ^ t[80];
  assign t[64] = t[79] ^ t[81];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[49] ^ t[84];
  assign t[67] = t[60] ^ t[85];
  assign t[68] = t[62] ^ t[86];
  assign t[69] = t[80] & t[87];
  assign t[6] = ~(t[10]);
  assign t[70] = t[88] & t[89];
  assign t[71] = t[90] ^ t[82];
  assign t[72] = t[90] & t[91];
  assign t[73] = t[92] & t[90];
  assign t[74] = t[166] ^ t[168];
  assign t[75] = t[26] ? t[169] : t[93];
  assign t[76] = t[26] ? t[170] : t[94];
  assign t[77] = t[91] ^ t[95];
  assign t[78] = t[26] ? t[171] : t[96];
  assign t[79] = t[26] ? t[172] : t[97];
  assign t[7] = ~(t[11]);
  assign t[80] = t[48] ^ t[98];
  assign t[81] = t[26] ? t[173] : t[99];
  assign t[82] = t[100] ^ t[101];
  assign t[83] = t[102] & t[71];
  assign t[84] = t[103] ^ t[86];
  assign t[85] = t[104] ^ t[59];
  assign t[86] = t[76] ^ t[81];
  assign t[87] = t[105] ^ t[60];
  assign t[88] = t[65] ^ t[48];
  assign t[89] = t[78] ^ t[104];
  assign t[8] = ~(t[12]);
  assign t[90] = t[106] ^ t[107];
  assign t[91] = t[108] ^ t[109];
  assign t[92] = t[110] ^ t[107];
  assign t[93] = t[174] ^ t[175];
  assign t[94] = t[176] ^ t[177];
  assign t[95] = t[111] & t[112];
  assign t[96] = t[165] ^ t[178];
  assign t[97] = t[179] ^ t[180];
  assign t[98] = t[113] ^ t[114];
  assign t[99] = t[181] ^ t[182];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind540(x, y);
 input [129:0] x;
 output y;

 wire [448:0] t;
  assign t[0] = t[1] ? t[2] : t[148];
  assign t[100] = t[178] ^ t[179];
  assign t[101] = t[122] ^ t[97];
  assign t[102] = t[61] ^ t[123];
  assign t[103] = t[78] ^ t[120];
  assign t[104] = t[124] ^ t[83];
  assign t[105] = t[25] ? t[180] : t[125];
  assign t[106] = t[99] & t[126];
  assign t[107] = t[99] ^ t[120];
  assign t[108] = t[104] & t[127];
  assign t[109] = t[104] ^ t[120];
  assign t[10] = t[150] & t[16];
  assign t[110] = t[93] ^ t[71];
  assign t[111] = t[85] ^ t[128];
  assign t[112] = t[25] ? t[181] : t[129];
  assign t[113] = t[182] ^ t[183];
  assign t[114] = t[184] ^ t[185];
  assign t[115] = t[164] ^ t[186];
  assign t[116] = t[130] ^ t[131];
  assign t[117] = t[110] ^ t[76];
  assign t[118] = t[110] & t[76];
  assign t[119] = t[74] & t[132];
  assign t[11] = ~(t[17]);
  assign t[120] = t[124] & t[121];
  assign t[121] = t[133] ^ t[134];
  assign t[122] = t[135] ^ t[136];
  assign t[123] = t[88] ^ t[73];
  assign t[124] = t[137] ^ t[134];
  assign t[125] = t[187] ^ t[188];
  assign t[126] = t[121] & t[83];
  assign t[127] = t[78] & t[124];
  assign t[128] = t[95] ^ t[82];
  assign t[129] = t[189] ^ t[190];
  assign t[12] = ~(t[150]);
  assign t[130] = t[65] & t[82];
  assign t[131] = t[138] & t[81];
  assign t[132] = t[92] ^ t[139];
  assign t[133] = t[140] ^ t[141];
  assign t[134] = t[142] ^ t[119];
  assign t[135] = t[61] & t[123];
  assign t[136] = t[77] & t[73];
  assign t[137] = t[143] ^ t[144];
  assign t[138] = t[77] ^ t[54];
  assign t[139] = t[105] ^ t[71];
  assign t[13] = ~(t[18]);
  assign t[140] = t[145] ^ t[131];
  assign t[141] = t[90] & t[146];
  assign t[142] = t[54] & t[57];
  assign t[143] = t[147] ^ t[136];
  assign t[144] = t[111] & t[88];
  assign t[145] = t[81] ^ t[139];
  assign t[146] = t[82] ^ t[81];
  assign t[147] = t[77] ^ t[73];
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[19] ? t[151] : t[22];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[150] & t[24]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = (t[225]);
  assign t[183] = (t[226]);
  assign t[184] = (t[227]);
  assign t[185] = (t[228]);
  assign t[186] = (t[229]);
  assign t[187] = (t[230]);
  assign t[188] = (t[231]);
  assign t[189] = (t[232]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[233]);
  assign t[191] = t[234] ^ x[2];
  assign t[192] = t[235] ^ x[5];
  assign t[193] = t[236] ^ x[9];
  assign t[194] = t[237] ^ x[12];
  assign t[195] = t[238] ^ x[15];
  assign t[196] = t[239] ^ x[18];
  assign t[197] = t[240] ^ x[21];
  assign t[198] = t[241] ^ x[24];
  assign t[199] = t[242] ^ x[27];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[30];
  assign t[201] = t[244] ^ x[33];
  assign t[202] = t[245] ^ x[36];
  assign t[203] = t[246] ^ x[39];
  assign t[204] = t[247] ^ x[42];
  assign t[205] = t[248] ^ x[45];
  assign t[206] = t[249] ^ x[48];
  assign t[207] = t[250] ^ x[51];
  assign t[208] = t[251] ^ x[54];
  assign t[209] = t[252] ^ x[57];
  assign t[20] = t[28] ^ t[29];
  assign t[210] = t[253] ^ x[60];
  assign t[211] = t[254] ^ x[63];
  assign t[212] = t[255] ^ x[66];
  assign t[213] = t[256] ^ x[69];
  assign t[214] = t[257] ^ x[72];
  assign t[215] = t[258] ^ x[75];
  assign t[216] = t[259] ^ x[78];
  assign t[217] = t[260] ^ x[81];
  assign t[218] = t[261] ^ x[84];
  assign t[219] = t[262] ^ x[87];
  assign t[21] = t[152] ^ t[153];
  assign t[220] = t[263] ^ x[90];
  assign t[221] = t[264] ^ x[93];
  assign t[222] = t[265] ^ x[96];
  assign t[223] = t[266] ^ x[99];
  assign t[224] = t[267] ^ x[102];
  assign t[225] = t[268] ^ x[105];
  assign t[226] = t[269] ^ x[108];
  assign t[227] = t[270] ^ x[111];
  assign t[228] = t[271] ^ x[114];
  assign t[229] = t[272] ^ x[117];
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = t[273] ^ x[120];
  assign t[231] = t[274] ^ x[123];
  assign t[232] = t[275] ^ x[126];
  assign t[233] = t[276] ^ x[129];
  assign t[234] = (t[277] & ~t[278]);
  assign t[235] = (t[279] & ~t[280]);
  assign t[236] = (t[281] & ~t[282]);
  assign t[237] = (t[283] & ~t[284]);
  assign t[238] = (t[285] & ~t[286]);
  assign t[239] = (t[287] & ~t[288]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[289] & ~t[290]);
  assign t[241] = (t[291] & ~t[292]);
  assign t[242] = (t[293] & ~t[294]);
  assign t[243] = (t[295] & ~t[296]);
  assign t[244] = (t[297] & ~t[298]);
  assign t[245] = (t[299] & ~t[300]);
  assign t[246] = (t[301] & ~t[302]);
  assign t[247] = (t[303] & ~t[304]);
  assign t[248] = (t[305] & ~t[306]);
  assign t[249] = (t[307] & ~t[308]);
  assign t[24] = ~(t[154] | t[34]);
  assign t[250] = (t[309] & ~t[310]);
  assign t[251] = (t[311] & ~t[312]);
  assign t[252] = (t[313] & ~t[314]);
  assign t[253] = (t[315] & ~t[316]);
  assign t[254] = (t[317] & ~t[318]);
  assign t[255] = (t[319] & ~t[320]);
  assign t[256] = (t[321] & ~t[322]);
  assign t[257] = (t[323] & ~t[324]);
  assign t[258] = (t[325] & ~t[326]);
  assign t[259] = (t[327] & ~t[328]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[329] & ~t[330]);
  assign t[261] = (t[331] & ~t[332]);
  assign t[262] = (t[333] & ~t[334]);
  assign t[263] = (t[335] & ~t[336]);
  assign t[264] = (t[337] & ~t[338]);
  assign t[265] = (t[339] & ~t[340]);
  assign t[266] = (t[341] & ~t[342]);
  assign t[267] = (t[343] & ~t[344]);
  assign t[268] = (t[345] & ~t[346]);
  assign t[269] = (t[347] & ~t[348]);
  assign t[26] = ~(t[155] & t[156]);
  assign t[270] = (t[349] & ~t[350]);
  assign t[271] = (t[351] & ~t[352]);
  assign t[272] = (t[353] & ~t[354]);
  assign t[273] = (t[355] & ~t[356]);
  assign t[274] = (t[357] & ~t[358]);
  assign t[275] = (t[359] & ~t[360]);
  assign t[276] = (t[361] & ~t[362]);
  assign t[277] = t[363] ^ x[2];
  assign t[278] = t[364] ^ x[1];
  assign t[279] = t[365] ^ x[5];
  assign t[27] = ~(t[157] & t[158]);
  assign t[280] = t[366] ^ x[4];
  assign t[281] = t[367] ^ x[9];
  assign t[282] = t[368] ^ x[8];
  assign t[283] = t[369] ^ x[12];
  assign t[284] = t[370] ^ x[11];
  assign t[285] = t[371] ^ x[15];
  assign t[286] = t[372] ^ x[14];
  assign t[287] = t[373] ^ x[18];
  assign t[288] = t[374] ^ x[17];
  assign t[289] = t[375] ^ x[21];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[376] ^ x[20];
  assign t[291] = t[377] ^ x[24];
  assign t[292] = t[378] ^ x[23];
  assign t[293] = t[379] ^ x[27];
  assign t[294] = t[380] ^ x[26];
  assign t[295] = t[381] ^ x[30];
  assign t[296] = t[382] ^ x[29];
  assign t[297] = t[383] ^ x[33];
  assign t[298] = t[384] ^ x[32];
  assign t[299] = t[385] ^ x[36];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[149] : t[5];
  assign t[300] = t[386] ^ x[35];
  assign t[301] = t[387] ^ x[39];
  assign t[302] = t[388] ^ x[38];
  assign t[303] = t[389] ^ x[42];
  assign t[304] = t[390] ^ x[41];
  assign t[305] = t[391] ^ x[45];
  assign t[306] = t[392] ^ x[44];
  assign t[307] = t[393] ^ x[48];
  assign t[308] = t[394] ^ x[47];
  assign t[309] = t[395] ^ x[51];
  assign t[30] = t[159] ^ t[41];
  assign t[310] = t[396] ^ x[50];
  assign t[311] = t[397] ^ x[54];
  assign t[312] = t[398] ^ x[53];
  assign t[313] = t[399] ^ x[57];
  assign t[314] = t[400] ^ x[56];
  assign t[315] = t[401] ^ x[60];
  assign t[316] = t[402] ^ x[59];
  assign t[317] = t[403] ^ x[63];
  assign t[318] = t[404] ^ x[62];
  assign t[319] = t[405] ^ x[66];
  assign t[31] = ~(t[160] ^ t[161]);
  assign t[320] = t[406] ^ x[65];
  assign t[321] = t[407] ^ x[69];
  assign t[322] = t[408] ^ x[68];
  assign t[323] = t[409] ^ x[72];
  assign t[324] = t[410] ^ x[71];
  assign t[325] = t[411] ^ x[75];
  assign t[326] = t[412] ^ x[74];
  assign t[327] = t[413] ^ x[78];
  assign t[328] = t[414] ^ x[77];
  assign t[329] = t[415] ^ x[81];
  assign t[32] = ~(t[24]);
  assign t[330] = t[416] ^ x[80];
  assign t[331] = t[417] ^ x[84];
  assign t[332] = t[418] ^ x[83];
  assign t[333] = t[419] ^ x[87];
  assign t[334] = t[420] ^ x[86];
  assign t[335] = t[421] ^ x[90];
  assign t[336] = t[422] ^ x[89];
  assign t[337] = t[423] ^ x[93];
  assign t[338] = t[424] ^ x[92];
  assign t[339] = t[425] ^ x[96];
  assign t[33] = ~(t[162] & t[42]);
  assign t[340] = t[426] ^ x[95];
  assign t[341] = t[427] ^ x[99];
  assign t[342] = t[428] ^ x[98];
  assign t[343] = t[429] ^ x[102];
  assign t[344] = t[430] ^ x[101];
  assign t[345] = t[431] ^ x[105];
  assign t[346] = t[432] ^ x[104];
  assign t[347] = t[433] ^ x[108];
  assign t[348] = t[434] ^ x[107];
  assign t[349] = t[435] ^ x[111];
  assign t[34] = ~(t[43] & t[44]);
  assign t[350] = t[436] ^ x[110];
  assign t[351] = t[437] ^ x[114];
  assign t[352] = t[438] ^ x[113];
  assign t[353] = t[439] ^ x[117];
  assign t[354] = t[440] ^ x[116];
  assign t[355] = t[441] ^ x[120];
  assign t[356] = t[442] ^ x[119];
  assign t[357] = t[443] ^ x[123];
  assign t[358] = t[444] ^ x[122];
  assign t[359] = t[445] ^ x[126];
  assign t[35] = ~(t[163]);
  assign t[360] = t[446] ^ x[125];
  assign t[361] = t[447] ^ x[129];
  assign t[362] = t[448] ^ x[128];
  assign t[363] = (x[0]);
  assign t[364] = (x[0]);
  assign t[365] = (x[3]);
  assign t[366] = (x[3]);
  assign t[367] = (x[7]);
  assign t[368] = (x[7]);
  assign t[369] = (x[10]);
  assign t[36] = ~(t[150]);
  assign t[370] = (x[10]);
  assign t[371] = (x[13]);
  assign t[372] = (x[13]);
  assign t[373] = (x[16]);
  assign t[374] = (x[16]);
  assign t[375] = (x[19]);
  assign t[376] = (x[19]);
  assign t[377] = (x[22]);
  assign t[378] = (x[22]);
  assign t[379] = (x[25]);
  assign t[37] = t[45] ^ t[46];
  assign t[380] = (x[25]);
  assign t[381] = (x[28]);
  assign t[382] = (x[28]);
  assign t[383] = (x[31]);
  assign t[384] = (x[31]);
  assign t[385] = (x[34]);
  assign t[386] = (x[34]);
  assign t[387] = (x[37]);
  assign t[388] = (x[37]);
  assign t[389] = (x[40]);
  assign t[38] = t[47] ^ t[48];
  assign t[390] = (x[40]);
  assign t[391] = (x[43]);
  assign t[392] = (x[43]);
  assign t[393] = (x[46]);
  assign t[394] = (x[46]);
  assign t[395] = (x[49]);
  assign t[396] = (x[49]);
  assign t[397] = (x[52]);
  assign t[398] = (x[52]);
  assign t[399] = (x[55]);
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[55]);
  assign t[401] = (x[58]);
  assign t[402] = (x[58]);
  assign t[403] = (x[61]);
  assign t[404] = (x[61]);
  assign t[405] = (x[64]);
  assign t[406] = (x[64]);
  assign t[407] = (x[67]);
  assign t[408] = (x[67]);
  assign t[409] = (x[70]);
  assign t[40] = t[51] ^ t[52];
  assign t[410] = (x[70]);
  assign t[411] = (x[73]);
  assign t[412] = (x[73]);
  assign t[413] = (x[76]);
  assign t[414] = (x[76]);
  assign t[415] = (x[79]);
  assign t[416] = (x[79]);
  assign t[417] = (x[82]);
  assign t[418] = (x[82]);
  assign t[419] = (x[85]);
  assign t[41] = t[152] ^ t[164];
  assign t[420] = (x[85]);
  assign t[421] = (x[88]);
  assign t[422] = (x[88]);
  assign t[423] = (x[91]);
  assign t[424] = (x[91]);
  assign t[425] = (x[94]);
  assign t[426] = (x[94]);
  assign t[427] = (x[97]);
  assign t[428] = (x[97]);
  assign t[429] = (x[100]);
  assign t[42] = ~(t[165]);
  assign t[430] = (x[100]);
  assign t[431] = (x[103]);
  assign t[432] = (x[103]);
  assign t[433] = (x[106]);
  assign t[434] = (x[106]);
  assign t[435] = (x[109]);
  assign t[436] = (x[109]);
  assign t[437] = (x[112]);
  assign t[438] = (x[112]);
  assign t[439] = (x[115]);
  assign t[43] = ~(t[166] | t[167]);
  assign t[440] = (x[115]);
  assign t[441] = (x[118]);
  assign t[442] = (x[118]);
  assign t[443] = (x[121]);
  assign t[444] = (x[121]);
  assign t[445] = (x[124]);
  assign t[446] = (x[124]);
  assign t[447] = (x[127]);
  assign t[448] = (x[127]);
  assign t[44] = ~(t[168] | t[169]);
  assign t[45] = t[53] & t[54];
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[53] & t[57];
  assign t[48] = t[58] ^ t[59];
  assign t[49] = t[60] & t[61];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] ^ t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[66] ^ t[67];
  assign t[53] = t[68] ^ t[69];
  assign t[54] = t[70] ^ t[71];
  assign t[55] = t[72] & t[73];
  assign t[56] = t[68] & t[74];
  assign t[57] = t[74] ^ t[75];
  assign t[58] = t[69] & t[76];
  assign t[59] = t[72] & t[77];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[78] ^ t[79];
  assign t[61] = t[74] ^ t[65];
  assign t[62] = t[80] & t[81];
  assign t[63] = t[64] & t[82];
  assign t[64] = t[83] ^ t[84];
  assign t[65] = t[85] ^ t[86];
  assign t[66] = t[87] & t[88];
  assign t[67] = t[89] & t[90];
  assign t[68] = t[60] ^ t[64];
  assign t[69] = t[87] ^ t[89];
  assign t[6] = ~(t[10]);
  assign t[70] = t[25] ? t[170] : t[91];
  assign t[71] = t[25] ? t[171] : t[21];
  assign t[72] = t[60] ^ t[87];
  assign t[73] = t[92] ^ t[75];
  assign t[74] = t[93] ^ t[70];
  assign t[75] = t[94] ^ t[71];
  assign t[76] = t[81] ^ t[85];
  assign t[77] = t[93] ^ t[95];
  assign t[78] = t[96] ^ t[97];
  assign t[79] = t[98] & t[99];
  assign t[7] = ~(t[11]);
  assign t[80] = t[64] ^ t[89];
  assign t[81] = t[74] ^ t[92];
  assign t[82] = t[25] ? t[172] : t[100];
  assign t[83] = t[101] ^ t[102];
  assign t[84] = t[103] & t[104];
  assign t[85] = t[105] ^ t[94];
  assign t[86] = t[70] ^ t[82];
  assign t[87] = t[106] ^ t[107];
  assign t[88] = t[82] ^ t[85];
  assign t[89] = t[108] ^ t[109];
  assign t[8] = ~(t[12]);
  assign t[90] = t[110] ^ t[111];
  assign t[91] = t[173] ^ t[174];
  assign t[92] = t[112] ^ t[95];
  assign t[93] = t[25] ? t[175] : t[113];
  assign t[94] = t[25] ? t[176] : t[114];
  assign t[95] = t[25] ? t[177] : t[115];
  assign t[96] = t[116] ^ t[117];
  assign t[97] = t[118] ^ t[119];
  assign t[98] = t[83] ^ t[120];
  assign t[99] = t[121] ^ t[78];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind541(x, y);
 input [129:0] x;
 output y;

 wire [448:0] t;
  assign t[0] = t[1] ? t[2] : t[148];
  assign t[100] = t[178] ^ t[179];
  assign t[101] = t[122] ^ t[97];
  assign t[102] = t[61] ^ t[123];
  assign t[103] = t[78] ^ t[120];
  assign t[104] = t[124] ^ t[83];
  assign t[105] = t[25] ? t[180] : t[125];
  assign t[106] = t[99] & t[126];
  assign t[107] = t[99] ^ t[120];
  assign t[108] = t[104] & t[127];
  assign t[109] = t[104] ^ t[120];
  assign t[10] = t[150] & t[16];
  assign t[110] = t[93] ^ t[71];
  assign t[111] = t[85] ^ t[128];
  assign t[112] = t[25] ? t[181] : t[129];
  assign t[113] = t[182] ^ t[183];
  assign t[114] = t[184] ^ t[185];
  assign t[115] = t[164] ^ t[186];
  assign t[116] = t[130] ^ t[131];
  assign t[117] = t[110] ^ t[76];
  assign t[118] = t[110] & t[76];
  assign t[119] = t[74] & t[132];
  assign t[11] = ~(t[17]);
  assign t[120] = t[124] & t[121];
  assign t[121] = t[133] ^ t[134];
  assign t[122] = t[135] ^ t[136];
  assign t[123] = t[88] ^ t[73];
  assign t[124] = t[137] ^ t[134];
  assign t[125] = t[187] ^ t[188];
  assign t[126] = t[121] & t[83];
  assign t[127] = t[78] & t[124];
  assign t[128] = t[95] ^ t[82];
  assign t[129] = t[189] ^ t[190];
  assign t[12] = ~(t[150]);
  assign t[130] = t[65] & t[82];
  assign t[131] = t[138] & t[81];
  assign t[132] = t[92] ^ t[139];
  assign t[133] = t[140] ^ t[141];
  assign t[134] = t[142] ^ t[119];
  assign t[135] = t[61] & t[123];
  assign t[136] = t[77] & t[73];
  assign t[137] = t[143] ^ t[144];
  assign t[138] = t[77] ^ t[54];
  assign t[139] = t[105] ^ t[71];
  assign t[13] = ~(t[18]);
  assign t[140] = t[145] ^ t[131];
  assign t[141] = t[90] & t[146];
  assign t[142] = t[54] & t[57];
  assign t[143] = t[147] ^ t[136];
  assign t[144] = t[111] & t[88];
  assign t[145] = t[81] ^ t[139];
  assign t[146] = t[82] ^ t[81];
  assign t[147] = t[77] ^ t[73];
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[19] ? t[151] : t[22];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[150] & t[24]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = (t[225]);
  assign t[183] = (t[226]);
  assign t[184] = (t[227]);
  assign t[185] = (t[228]);
  assign t[186] = (t[229]);
  assign t[187] = (t[230]);
  assign t[188] = (t[231]);
  assign t[189] = (t[232]);
  assign t[18] = ~(t[25]);
  assign t[190] = (t[233]);
  assign t[191] = t[234] ^ x[2];
  assign t[192] = t[235] ^ x[5];
  assign t[193] = t[236] ^ x[9];
  assign t[194] = t[237] ^ x[12];
  assign t[195] = t[238] ^ x[15];
  assign t[196] = t[239] ^ x[18];
  assign t[197] = t[240] ^ x[21];
  assign t[198] = t[241] ^ x[24];
  assign t[199] = t[242] ^ x[27];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[30];
  assign t[201] = t[244] ^ x[33];
  assign t[202] = t[245] ^ x[36];
  assign t[203] = t[246] ^ x[39];
  assign t[204] = t[247] ^ x[42];
  assign t[205] = t[248] ^ x[45];
  assign t[206] = t[249] ^ x[48];
  assign t[207] = t[250] ^ x[51];
  assign t[208] = t[251] ^ x[54];
  assign t[209] = t[252] ^ x[57];
  assign t[20] = t[28] ^ t[29];
  assign t[210] = t[253] ^ x[60];
  assign t[211] = t[254] ^ x[63];
  assign t[212] = t[255] ^ x[66];
  assign t[213] = t[256] ^ x[69];
  assign t[214] = t[257] ^ x[72];
  assign t[215] = t[258] ^ x[75];
  assign t[216] = t[259] ^ x[78];
  assign t[217] = t[260] ^ x[81];
  assign t[218] = t[261] ^ x[84];
  assign t[219] = t[262] ^ x[87];
  assign t[21] = t[152] ^ t[153];
  assign t[220] = t[263] ^ x[90];
  assign t[221] = t[264] ^ x[93];
  assign t[222] = t[265] ^ x[96];
  assign t[223] = t[266] ^ x[99];
  assign t[224] = t[267] ^ x[102];
  assign t[225] = t[268] ^ x[105];
  assign t[226] = t[269] ^ x[108];
  assign t[227] = t[270] ^ x[111];
  assign t[228] = t[271] ^ x[114];
  assign t[229] = t[272] ^ x[117];
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = t[273] ^ x[120];
  assign t[231] = t[274] ^ x[123];
  assign t[232] = t[275] ^ x[126];
  assign t[233] = t[276] ^ x[129];
  assign t[234] = (t[277] & ~t[278]);
  assign t[235] = (t[279] & ~t[280]);
  assign t[236] = (t[281] & ~t[282]);
  assign t[237] = (t[283] & ~t[284]);
  assign t[238] = (t[285] & ~t[286]);
  assign t[239] = (t[287] & ~t[288]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[289] & ~t[290]);
  assign t[241] = (t[291] & ~t[292]);
  assign t[242] = (t[293] & ~t[294]);
  assign t[243] = (t[295] & ~t[296]);
  assign t[244] = (t[297] & ~t[298]);
  assign t[245] = (t[299] & ~t[300]);
  assign t[246] = (t[301] & ~t[302]);
  assign t[247] = (t[303] & ~t[304]);
  assign t[248] = (t[305] & ~t[306]);
  assign t[249] = (t[307] & ~t[308]);
  assign t[24] = ~(t[154] | t[34]);
  assign t[250] = (t[309] & ~t[310]);
  assign t[251] = (t[311] & ~t[312]);
  assign t[252] = (t[313] & ~t[314]);
  assign t[253] = (t[315] & ~t[316]);
  assign t[254] = (t[317] & ~t[318]);
  assign t[255] = (t[319] & ~t[320]);
  assign t[256] = (t[321] & ~t[322]);
  assign t[257] = (t[323] & ~t[324]);
  assign t[258] = (t[325] & ~t[326]);
  assign t[259] = (t[327] & ~t[328]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[329] & ~t[330]);
  assign t[261] = (t[331] & ~t[332]);
  assign t[262] = (t[333] & ~t[334]);
  assign t[263] = (t[335] & ~t[336]);
  assign t[264] = (t[337] & ~t[338]);
  assign t[265] = (t[339] & ~t[340]);
  assign t[266] = (t[341] & ~t[342]);
  assign t[267] = (t[343] & ~t[344]);
  assign t[268] = (t[345] & ~t[346]);
  assign t[269] = (t[347] & ~t[348]);
  assign t[26] = ~(t[155] & t[156]);
  assign t[270] = (t[349] & ~t[350]);
  assign t[271] = (t[351] & ~t[352]);
  assign t[272] = (t[353] & ~t[354]);
  assign t[273] = (t[355] & ~t[356]);
  assign t[274] = (t[357] & ~t[358]);
  assign t[275] = (t[359] & ~t[360]);
  assign t[276] = (t[361] & ~t[362]);
  assign t[277] = t[363] ^ x[2];
  assign t[278] = t[364] ^ x[1];
  assign t[279] = t[365] ^ x[5];
  assign t[27] = ~(t[157] & t[158]);
  assign t[280] = t[366] ^ x[4];
  assign t[281] = t[367] ^ x[9];
  assign t[282] = t[368] ^ x[8];
  assign t[283] = t[369] ^ x[12];
  assign t[284] = t[370] ^ x[11];
  assign t[285] = t[371] ^ x[15];
  assign t[286] = t[372] ^ x[14];
  assign t[287] = t[373] ^ x[18];
  assign t[288] = t[374] ^ x[17];
  assign t[289] = t[375] ^ x[21];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[376] ^ x[20];
  assign t[291] = t[377] ^ x[24];
  assign t[292] = t[378] ^ x[23];
  assign t[293] = t[379] ^ x[27];
  assign t[294] = t[380] ^ x[26];
  assign t[295] = t[381] ^ x[30];
  assign t[296] = t[382] ^ x[29];
  assign t[297] = t[383] ^ x[33];
  assign t[298] = t[384] ^ x[32];
  assign t[299] = t[385] ^ x[36];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[149] : t[5];
  assign t[300] = t[386] ^ x[35];
  assign t[301] = t[387] ^ x[39];
  assign t[302] = t[388] ^ x[38];
  assign t[303] = t[389] ^ x[42];
  assign t[304] = t[390] ^ x[41];
  assign t[305] = t[391] ^ x[45];
  assign t[306] = t[392] ^ x[44];
  assign t[307] = t[393] ^ x[48];
  assign t[308] = t[394] ^ x[47];
  assign t[309] = t[395] ^ x[51];
  assign t[30] = t[159] ^ t[41];
  assign t[310] = t[396] ^ x[50];
  assign t[311] = t[397] ^ x[54];
  assign t[312] = t[398] ^ x[53];
  assign t[313] = t[399] ^ x[57];
  assign t[314] = t[400] ^ x[56];
  assign t[315] = t[401] ^ x[60];
  assign t[316] = t[402] ^ x[59];
  assign t[317] = t[403] ^ x[63];
  assign t[318] = t[404] ^ x[62];
  assign t[319] = t[405] ^ x[66];
  assign t[31] = ~(t[160] ^ t[161]);
  assign t[320] = t[406] ^ x[65];
  assign t[321] = t[407] ^ x[69];
  assign t[322] = t[408] ^ x[68];
  assign t[323] = t[409] ^ x[72];
  assign t[324] = t[410] ^ x[71];
  assign t[325] = t[411] ^ x[75];
  assign t[326] = t[412] ^ x[74];
  assign t[327] = t[413] ^ x[78];
  assign t[328] = t[414] ^ x[77];
  assign t[329] = t[415] ^ x[81];
  assign t[32] = ~(t[24]);
  assign t[330] = t[416] ^ x[80];
  assign t[331] = t[417] ^ x[84];
  assign t[332] = t[418] ^ x[83];
  assign t[333] = t[419] ^ x[87];
  assign t[334] = t[420] ^ x[86];
  assign t[335] = t[421] ^ x[90];
  assign t[336] = t[422] ^ x[89];
  assign t[337] = t[423] ^ x[93];
  assign t[338] = t[424] ^ x[92];
  assign t[339] = t[425] ^ x[96];
  assign t[33] = ~(t[162] & t[42]);
  assign t[340] = t[426] ^ x[95];
  assign t[341] = t[427] ^ x[99];
  assign t[342] = t[428] ^ x[98];
  assign t[343] = t[429] ^ x[102];
  assign t[344] = t[430] ^ x[101];
  assign t[345] = t[431] ^ x[105];
  assign t[346] = t[432] ^ x[104];
  assign t[347] = t[433] ^ x[108];
  assign t[348] = t[434] ^ x[107];
  assign t[349] = t[435] ^ x[111];
  assign t[34] = ~(t[43] & t[44]);
  assign t[350] = t[436] ^ x[110];
  assign t[351] = t[437] ^ x[114];
  assign t[352] = t[438] ^ x[113];
  assign t[353] = t[439] ^ x[117];
  assign t[354] = t[440] ^ x[116];
  assign t[355] = t[441] ^ x[120];
  assign t[356] = t[442] ^ x[119];
  assign t[357] = t[443] ^ x[123];
  assign t[358] = t[444] ^ x[122];
  assign t[359] = t[445] ^ x[126];
  assign t[35] = ~(t[163]);
  assign t[360] = t[446] ^ x[125];
  assign t[361] = t[447] ^ x[129];
  assign t[362] = t[448] ^ x[128];
  assign t[363] = (x[0]);
  assign t[364] = (x[0]);
  assign t[365] = (x[3]);
  assign t[366] = (x[3]);
  assign t[367] = (x[7]);
  assign t[368] = (x[7]);
  assign t[369] = (x[10]);
  assign t[36] = ~(t[150]);
  assign t[370] = (x[10]);
  assign t[371] = (x[13]);
  assign t[372] = (x[13]);
  assign t[373] = (x[16]);
  assign t[374] = (x[16]);
  assign t[375] = (x[19]);
  assign t[376] = (x[19]);
  assign t[377] = (x[22]);
  assign t[378] = (x[22]);
  assign t[379] = (x[25]);
  assign t[37] = t[45] ^ t[46];
  assign t[380] = (x[25]);
  assign t[381] = (x[28]);
  assign t[382] = (x[28]);
  assign t[383] = (x[31]);
  assign t[384] = (x[31]);
  assign t[385] = (x[34]);
  assign t[386] = (x[34]);
  assign t[387] = (x[37]);
  assign t[388] = (x[37]);
  assign t[389] = (x[40]);
  assign t[38] = t[47] ^ t[48];
  assign t[390] = (x[40]);
  assign t[391] = (x[43]);
  assign t[392] = (x[43]);
  assign t[393] = (x[46]);
  assign t[394] = (x[46]);
  assign t[395] = (x[49]);
  assign t[396] = (x[49]);
  assign t[397] = (x[52]);
  assign t[398] = (x[52]);
  assign t[399] = (x[55]);
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[55]);
  assign t[401] = (x[58]);
  assign t[402] = (x[58]);
  assign t[403] = (x[61]);
  assign t[404] = (x[61]);
  assign t[405] = (x[64]);
  assign t[406] = (x[64]);
  assign t[407] = (x[67]);
  assign t[408] = (x[67]);
  assign t[409] = (x[70]);
  assign t[40] = t[51] ^ t[52];
  assign t[410] = (x[70]);
  assign t[411] = (x[73]);
  assign t[412] = (x[73]);
  assign t[413] = (x[76]);
  assign t[414] = (x[76]);
  assign t[415] = (x[79]);
  assign t[416] = (x[79]);
  assign t[417] = (x[82]);
  assign t[418] = (x[82]);
  assign t[419] = (x[85]);
  assign t[41] = t[152] ^ t[164];
  assign t[420] = (x[85]);
  assign t[421] = (x[88]);
  assign t[422] = (x[88]);
  assign t[423] = (x[91]);
  assign t[424] = (x[91]);
  assign t[425] = (x[94]);
  assign t[426] = (x[94]);
  assign t[427] = (x[97]);
  assign t[428] = (x[97]);
  assign t[429] = (x[100]);
  assign t[42] = ~(t[165]);
  assign t[430] = (x[100]);
  assign t[431] = (x[103]);
  assign t[432] = (x[103]);
  assign t[433] = (x[106]);
  assign t[434] = (x[106]);
  assign t[435] = (x[109]);
  assign t[436] = (x[109]);
  assign t[437] = (x[112]);
  assign t[438] = (x[112]);
  assign t[439] = (x[115]);
  assign t[43] = ~(t[166] | t[167]);
  assign t[440] = (x[115]);
  assign t[441] = (x[118]);
  assign t[442] = (x[118]);
  assign t[443] = (x[121]);
  assign t[444] = (x[121]);
  assign t[445] = (x[124]);
  assign t[446] = (x[124]);
  assign t[447] = (x[127]);
  assign t[448] = (x[127]);
  assign t[44] = ~(t[168] | t[169]);
  assign t[45] = t[53] & t[54];
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[53] & t[57];
  assign t[48] = t[58] ^ t[59];
  assign t[49] = t[60] & t[61];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] ^ t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[66] ^ t[67];
  assign t[53] = t[68] ^ t[69];
  assign t[54] = t[70] ^ t[71];
  assign t[55] = t[72] & t[73];
  assign t[56] = t[68] & t[74];
  assign t[57] = t[74] ^ t[75];
  assign t[58] = t[69] & t[76];
  assign t[59] = t[72] & t[77];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[78] ^ t[79];
  assign t[61] = t[74] ^ t[65];
  assign t[62] = t[80] & t[81];
  assign t[63] = t[64] & t[82];
  assign t[64] = t[83] ^ t[84];
  assign t[65] = t[85] ^ t[86];
  assign t[66] = t[87] & t[88];
  assign t[67] = t[89] & t[90];
  assign t[68] = t[60] ^ t[64];
  assign t[69] = t[87] ^ t[89];
  assign t[6] = ~(t[10]);
  assign t[70] = t[25] ? t[170] : t[91];
  assign t[71] = t[25] ? t[171] : t[21];
  assign t[72] = t[60] ^ t[87];
  assign t[73] = t[92] ^ t[75];
  assign t[74] = t[93] ^ t[70];
  assign t[75] = t[94] ^ t[71];
  assign t[76] = t[81] ^ t[85];
  assign t[77] = t[93] ^ t[95];
  assign t[78] = t[96] ^ t[97];
  assign t[79] = t[98] & t[99];
  assign t[7] = ~(t[11]);
  assign t[80] = t[64] ^ t[89];
  assign t[81] = t[74] ^ t[92];
  assign t[82] = t[25] ? t[172] : t[100];
  assign t[83] = t[101] ^ t[102];
  assign t[84] = t[103] & t[104];
  assign t[85] = t[105] ^ t[94];
  assign t[86] = t[70] ^ t[82];
  assign t[87] = t[106] ^ t[107];
  assign t[88] = t[82] ^ t[85];
  assign t[89] = t[108] ^ t[109];
  assign t[8] = ~(t[12]);
  assign t[90] = t[110] ^ t[111];
  assign t[91] = t[173] ^ t[174];
  assign t[92] = t[112] ^ t[95];
  assign t[93] = t[25] ? t[175] : t[113];
  assign t[94] = t[25] ? t[176] : t[114];
  assign t[95] = t[25] ? t[177] : t[115];
  assign t[96] = t[116] ^ t[117];
  assign t[97] = t[118] ^ t[119];
  assign t[98] = t[83] ^ t[120];
  assign t[99] = t[121] ^ t[78];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind542(x, y);
 input [132:0] x;
 output y;

 wire [448:0] t;
  assign t[0] = t[1] ? t[2] : t[141];
  assign t[100] = t[113] ^ t[101];
  assign t[101] = t[25] ? t[177] : t[114];
  assign t[102] = t[115] ^ t[106];
  assign t[103] = t[116] ^ t[69];
  assign t[104] = t[86] ^ t[94];
  assign t[105] = t[117] ^ t[118];
  assign t[106] = t[119] ^ t[120];
  assign t[107] = t[83] ^ t[94];
  assign t[108] = t[96] ^ t[73];
  assign t[109] = t[121] ^ t[122];
  assign t[10] = t[143] & t[16];
  assign t[110] = t[123] ^ t[122];
  assign t[111] = t[178] ^ t[179];
  assign t[112] = t[180] ^ t[181];
  assign t[113] = t[25] ? t[182] : t[21];
  assign t[114] = t[183] ^ t[184];
  assign t[115] = t[124] ^ t[125];
  assign t[116] = t[56] ^ t[126];
  assign t[117] = t[127] ^ t[128];
  assign t[118] = t[79] ^ t[129];
  assign t[119] = t[79] & t[129];
  assign t[11] = ~(t[17]);
  assign t[120] = t[56] & t[130];
  assign t[121] = t[131] ^ t[132];
  assign t[122] = t[133] ^ t[120];
  assign t[123] = t[134] ^ t[135];
  assign t[124] = t[116] & t[69];
  assign t[125] = t[82] & t[88];
  assign t[126] = t[76] ^ t[136];
  assign t[127] = t[126] & t[67];
  assign t[128] = t[65] & t[81];
  assign t[129] = t[81] ^ t[76];
  assign t[12] = ~(t[143]);
  assign t[130] = t[100] ^ t[137];
  assign t[131] = t[138] ^ t[128];
  assign t[132] = t[62] & t[63];
  assign t[133] = t[58] & t[139];
  assign t[134] = t[140] ^ t[125];
  assign t[135] = t[80] & t[60];
  assign t[136] = t[71] ^ t[67];
  assign t[137] = t[95] ^ t[73];
  assign t[138] = t[81] ^ t[137];
  assign t[139] = t[56] ^ t[108];
  assign t[13] = ~(t[18]);
  assign t[140] = t[82] ^ t[88];
  assign t[141] = (t[185]);
  assign t[142] = (t[186]);
  assign t[143] = (t[187]);
  assign t[144] = (t[188]);
  assign t[145] = (t[189]);
  assign t[146] = (t[190]);
  assign t[147] = (t[191]);
  assign t[148] = (t[192]);
  assign t[149] = (t[193]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[194]);
  assign t[151] = (t[195]);
  assign t[152] = (t[196]);
  assign t[153] = (t[197]);
  assign t[154] = (t[198]);
  assign t[155] = (t[199]);
  assign t[156] = (t[200]);
  assign t[157] = (t[201]);
  assign t[158] = (t[202]);
  assign t[159] = (t[203]);
  assign t[15] = t[19] ? t[144] : t[22];
  assign t[160] = (t[204]);
  assign t[161] = (t[205]);
  assign t[162] = (t[206]);
  assign t[163] = (t[207]);
  assign t[164] = (t[208]);
  assign t[165] = (t[209]);
  assign t[166] = (t[210]);
  assign t[167] = (t[211]);
  assign t[168] = (t[212]);
  assign t[169] = (t[213]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[214]);
  assign t[171] = (t[215]);
  assign t[172] = (t[216]);
  assign t[173] = (t[217]);
  assign t[174] = (t[218]);
  assign t[175] = (t[219]);
  assign t[176] = (t[220]);
  assign t[177] = (t[221]);
  assign t[178] = (t[222]);
  assign t[179] = (t[223]);
  assign t[17] = ~(t[143] & t[24]);
  assign t[180] = (t[224]);
  assign t[181] = (t[225]);
  assign t[182] = (t[226]);
  assign t[183] = (t[227]);
  assign t[184] = (t[228]);
  assign t[185] = t[229] ^ x[2];
  assign t[186] = t[230] ^ x[5];
  assign t[187] = t[231] ^ x[9];
  assign t[188] = t[232] ^ x[12];
  assign t[189] = t[233] ^ x[15];
  assign t[18] = ~(t[25]);
  assign t[190] = t[234] ^ x[18];
  assign t[191] = t[235] ^ x[21];
  assign t[192] = t[236] ^ x[24];
  assign t[193] = t[237] ^ x[27];
  assign t[194] = t[238] ^ x[30];
  assign t[195] = t[239] ^ x[33];
  assign t[196] = t[240] ^ x[36];
  assign t[197] = t[241] ^ x[39];
  assign t[198] = t[242] ^ x[42];
  assign t[199] = t[243] ^ x[45];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[244] ^ x[48];
  assign t[201] = t[245] ^ x[51];
  assign t[202] = t[246] ^ x[54];
  assign t[203] = t[247] ^ x[57];
  assign t[204] = t[248] ^ x[60];
  assign t[205] = t[249] ^ x[63];
  assign t[206] = t[250] ^ x[66];
  assign t[207] = t[251] ^ x[69];
  assign t[208] = t[252] ^ x[72];
  assign t[209] = t[253] ^ x[75];
  assign t[20] = t[28] ^ t[29];
  assign t[210] = t[254] ^ x[78];
  assign t[211] = t[255] ^ x[81];
  assign t[212] = t[256] ^ x[84];
  assign t[213] = t[257] ^ x[87];
  assign t[214] = t[258] ^ x[90];
  assign t[215] = t[259] ^ x[93];
  assign t[216] = t[260] ^ x[96];
  assign t[217] = t[261] ^ x[99];
  assign t[218] = t[262] ^ x[102];
  assign t[219] = t[263] ^ x[105];
  assign t[21] = t[145] ^ t[146];
  assign t[220] = t[264] ^ x[108];
  assign t[221] = t[265] ^ x[111];
  assign t[222] = t[266] ^ x[114];
  assign t[223] = t[267] ^ x[117];
  assign t[224] = t[268] ^ x[120];
  assign t[225] = t[269] ^ x[123];
  assign t[226] = t[270] ^ x[126];
  assign t[227] = t[271] ^ x[129];
  assign t[228] = t[272] ^ x[132];
  assign t[229] = (t[273] & ~t[274]);
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[275] & ~t[276]);
  assign t[231] = (t[277] & ~t[278]);
  assign t[232] = (t[279] & ~t[280]);
  assign t[233] = (t[281] & ~t[282]);
  assign t[234] = (t[283] & ~t[284]);
  assign t[235] = (t[285] & ~t[286]);
  assign t[236] = (t[287] & ~t[288]);
  assign t[237] = (t[289] & ~t[290]);
  assign t[238] = (t[291] & ~t[292]);
  assign t[239] = (t[293] & ~t[294]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[295] & ~t[296]);
  assign t[241] = (t[297] & ~t[298]);
  assign t[242] = (t[299] & ~t[300]);
  assign t[243] = (t[301] & ~t[302]);
  assign t[244] = (t[303] & ~t[304]);
  assign t[245] = (t[305] & ~t[306]);
  assign t[246] = (t[307] & ~t[308]);
  assign t[247] = (t[309] & ~t[310]);
  assign t[248] = (t[311] & ~t[312]);
  assign t[249] = (t[313] & ~t[314]);
  assign t[24] = ~(t[147] | t[34]);
  assign t[250] = (t[315] & ~t[316]);
  assign t[251] = (t[317] & ~t[318]);
  assign t[252] = (t[319] & ~t[320]);
  assign t[253] = (t[321] & ~t[322]);
  assign t[254] = (t[323] & ~t[324]);
  assign t[255] = (t[325] & ~t[326]);
  assign t[256] = (t[327] & ~t[328]);
  assign t[257] = (t[329] & ~t[330]);
  assign t[258] = (t[331] & ~t[332]);
  assign t[259] = (t[333] & ~t[334]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[335] & ~t[336]);
  assign t[261] = (t[337] & ~t[338]);
  assign t[262] = (t[339] & ~t[340]);
  assign t[263] = (t[341] & ~t[342]);
  assign t[264] = (t[343] & ~t[344]);
  assign t[265] = (t[345] & ~t[346]);
  assign t[266] = (t[347] & ~t[348]);
  assign t[267] = (t[349] & ~t[350]);
  assign t[268] = (t[351] & ~t[352]);
  assign t[269] = (t[353] & ~t[354]);
  assign t[26] = ~(t[148] & t[149]);
  assign t[270] = (t[355] & ~t[356]);
  assign t[271] = (t[357] & ~t[358]);
  assign t[272] = (t[359] & ~t[360]);
  assign t[273] = t[361] ^ x[2];
  assign t[274] = t[362] ^ x[1];
  assign t[275] = t[363] ^ x[5];
  assign t[276] = t[364] ^ x[4];
  assign t[277] = t[365] ^ x[9];
  assign t[278] = t[366] ^ x[8];
  assign t[279] = t[367] ^ x[12];
  assign t[27] = ~(t[150] & t[151]);
  assign t[280] = t[368] ^ x[11];
  assign t[281] = t[369] ^ x[15];
  assign t[282] = t[370] ^ x[14];
  assign t[283] = t[371] ^ x[18];
  assign t[284] = t[372] ^ x[17];
  assign t[285] = t[373] ^ x[21];
  assign t[286] = t[374] ^ x[20];
  assign t[287] = t[375] ^ x[24];
  assign t[288] = t[376] ^ x[23];
  assign t[289] = t[377] ^ x[27];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[378] ^ x[26];
  assign t[291] = t[379] ^ x[30];
  assign t[292] = t[380] ^ x[29];
  assign t[293] = t[381] ^ x[33];
  assign t[294] = t[382] ^ x[32];
  assign t[295] = t[383] ^ x[36];
  assign t[296] = t[384] ^ x[35];
  assign t[297] = t[385] ^ x[39];
  assign t[298] = t[386] ^ x[38];
  assign t[299] = t[387] ^ x[42];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[142] : t[5];
  assign t[300] = t[388] ^ x[41];
  assign t[301] = t[389] ^ x[45];
  assign t[302] = t[390] ^ x[44];
  assign t[303] = t[391] ^ x[48];
  assign t[304] = t[392] ^ x[47];
  assign t[305] = t[393] ^ x[51];
  assign t[306] = t[394] ^ x[50];
  assign t[307] = t[395] ^ x[54];
  assign t[308] = t[396] ^ x[53];
  assign t[309] = t[397] ^ x[57];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[398] ^ x[56];
  assign t[311] = t[399] ^ x[60];
  assign t[312] = t[400] ^ x[59];
  assign t[313] = t[401] ^ x[63];
  assign t[314] = t[402] ^ x[62];
  assign t[315] = t[403] ^ x[66];
  assign t[316] = t[404] ^ x[65];
  assign t[317] = t[405] ^ x[69];
  assign t[318] = t[406] ^ x[68];
  assign t[319] = t[407] ^ x[72];
  assign t[31] = ~(t[152] ^ t[153]);
  assign t[320] = t[408] ^ x[71];
  assign t[321] = t[409] ^ x[75];
  assign t[322] = t[410] ^ x[74];
  assign t[323] = t[411] ^ x[78];
  assign t[324] = t[412] ^ x[77];
  assign t[325] = t[413] ^ x[81];
  assign t[326] = t[414] ^ x[80];
  assign t[327] = t[415] ^ x[84];
  assign t[328] = t[416] ^ x[83];
  assign t[329] = t[417] ^ x[87];
  assign t[32] = ~(t[24]);
  assign t[330] = t[418] ^ x[86];
  assign t[331] = t[419] ^ x[90];
  assign t[332] = t[420] ^ x[89];
  assign t[333] = t[421] ^ x[93];
  assign t[334] = t[422] ^ x[92];
  assign t[335] = t[423] ^ x[96];
  assign t[336] = t[424] ^ x[95];
  assign t[337] = t[425] ^ x[99];
  assign t[338] = t[426] ^ x[98];
  assign t[339] = t[427] ^ x[102];
  assign t[33] = ~(t[154] & t[43]);
  assign t[340] = t[428] ^ x[101];
  assign t[341] = t[429] ^ x[105];
  assign t[342] = t[430] ^ x[104];
  assign t[343] = t[431] ^ x[108];
  assign t[344] = t[432] ^ x[107];
  assign t[345] = t[433] ^ x[111];
  assign t[346] = t[434] ^ x[110];
  assign t[347] = t[435] ^ x[114];
  assign t[348] = t[436] ^ x[113];
  assign t[349] = t[437] ^ x[117];
  assign t[34] = ~(t[44] & t[45]);
  assign t[350] = t[438] ^ x[116];
  assign t[351] = t[439] ^ x[120];
  assign t[352] = t[440] ^ x[119];
  assign t[353] = t[441] ^ x[123];
  assign t[354] = t[442] ^ x[122];
  assign t[355] = t[443] ^ x[126];
  assign t[356] = t[444] ^ x[125];
  assign t[357] = t[445] ^ x[129];
  assign t[358] = t[446] ^ x[128];
  assign t[359] = t[447] ^ x[132];
  assign t[35] = ~(t[155]);
  assign t[360] = t[448] ^ x[131];
  assign t[361] = (x[0]);
  assign t[362] = (x[0]);
  assign t[363] = (x[3]);
  assign t[364] = (x[3]);
  assign t[365] = (x[7]);
  assign t[366] = (x[7]);
  assign t[367] = (x[10]);
  assign t[368] = (x[10]);
  assign t[369] = (x[13]);
  assign t[36] = ~(t[143]);
  assign t[370] = (x[13]);
  assign t[371] = (x[16]);
  assign t[372] = (x[16]);
  assign t[373] = (x[19]);
  assign t[374] = (x[19]);
  assign t[375] = (x[22]);
  assign t[376] = (x[22]);
  assign t[377] = (x[25]);
  assign t[378] = (x[25]);
  assign t[379] = (x[28]);
  assign t[37] = t[46] ^ t[47];
  assign t[380] = (x[28]);
  assign t[381] = (x[31]);
  assign t[382] = (x[31]);
  assign t[383] = (x[34]);
  assign t[384] = (x[34]);
  assign t[385] = (x[37]);
  assign t[386] = (x[37]);
  assign t[387] = (x[40]);
  assign t[388] = (x[40]);
  assign t[389] = (x[43]);
  assign t[38] = t[48] ^ t[49];
  assign t[390] = (x[43]);
  assign t[391] = (x[46]);
  assign t[392] = (x[46]);
  assign t[393] = (x[49]);
  assign t[394] = (x[49]);
  assign t[395] = (x[52]);
  assign t[396] = (x[52]);
  assign t[397] = (x[55]);
  assign t[398] = (x[55]);
  assign t[399] = (x[58]);
  assign t[39] = t[50] ^ t[51];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[58]);
  assign t[401] = (x[61]);
  assign t[402] = (x[61]);
  assign t[403] = (x[64]);
  assign t[404] = (x[64]);
  assign t[405] = (x[67]);
  assign t[406] = (x[67]);
  assign t[407] = (x[70]);
  assign t[408] = (x[70]);
  assign t[409] = (x[73]);
  assign t[40] = t[52] ^ t[53];
  assign t[410] = (x[73]);
  assign t[411] = (x[76]);
  assign t[412] = (x[76]);
  assign t[413] = (x[79]);
  assign t[414] = (x[79]);
  assign t[415] = (x[82]);
  assign t[416] = (x[82]);
  assign t[417] = (x[85]);
  assign t[418] = (x[85]);
  assign t[419] = (x[88]);
  assign t[41] = t[156] ^ t[157];
  assign t[420] = (x[88]);
  assign t[421] = (x[91]);
  assign t[422] = (x[91]);
  assign t[423] = (x[94]);
  assign t[424] = (x[94]);
  assign t[425] = (x[97]);
  assign t[426] = (x[97]);
  assign t[427] = (x[100]);
  assign t[428] = (x[100]);
  assign t[429] = (x[103]);
  assign t[42] = t[145] ^ t[54];
  assign t[430] = (x[103]);
  assign t[431] = (x[106]);
  assign t[432] = (x[106]);
  assign t[433] = (x[109]);
  assign t[434] = (x[109]);
  assign t[435] = (x[112]);
  assign t[436] = (x[112]);
  assign t[437] = (x[115]);
  assign t[438] = (x[115]);
  assign t[439] = (x[118]);
  assign t[43] = ~(t[158]);
  assign t[440] = (x[118]);
  assign t[441] = (x[121]);
  assign t[442] = (x[121]);
  assign t[443] = (x[124]);
  assign t[444] = (x[124]);
  assign t[445] = (x[127]);
  assign t[446] = (x[127]);
  assign t[447] = (x[130]);
  assign t[448] = (x[130]);
  assign t[44] = ~(t[159] | t[160]);
  assign t[45] = ~(t[161] | t[162]);
  assign t[46] = t[55] & t[56];
  assign t[47] = t[57] & t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[61] & t[62];
  assign t[4] = ~(t[7]);
  assign t[50] = t[61] & t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[66] & t[67];
  assign t[53] = t[68] & t[69];
  assign t[54] = t[163] ^ t[164];
  assign t[55] = t[68] ^ t[66];
  assign t[56] = t[70] ^ t[71];
  assign t[57] = t[55] ^ t[72];
  assign t[58] = t[71] ^ t[73];
  assign t[59] = t[74] ^ t[75];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[67] ^ t[76];
  assign t[61] = t[77] ^ t[78];
  assign t[62] = t[79] ^ t[80];
  assign t[63] = t[67] ^ t[81];
  assign t[64] = t[66] ^ t[61];
  assign t[65] = t[82] ^ t[58];
  assign t[66] = t[83] ^ t[84];
  assign t[67] = t[25] ? t[165] : t[85];
  assign t[68] = t[86] ^ t[87];
  assign t[69] = t[60] ^ t[88];
  assign t[6] = ~(t[10]);
  assign t[70] = t[25] ? t[166] : t[89];
  assign t[71] = t[25] ? t[167] : t[90];
  assign t[72] = t[59] ^ t[61];
  assign t[73] = t[25] ? t[168] : t[91];
  assign t[74] = t[92] & t[93];
  assign t[75] = t[92] ^ t[94];
  assign t[76] = t[95] ^ t[96];
  assign t[77] = t[97] & t[98];
  assign t[78] = t[97] ^ t[94];
  assign t[79] = t[70] ^ t[73];
  assign t[7] = ~(t[11]);
  assign t[80] = t[76] ^ t[99];
  assign t[81] = t[56] ^ t[100];
  assign t[82] = t[70] ^ t[101];
  assign t[83] = t[102] ^ t[103];
  assign t[84] = t[104] & t[97];
  assign t[85] = t[169] ^ t[170];
  assign t[86] = t[105] ^ t[106];
  assign t[87] = t[107] & t[92];
  assign t[88] = t[100] ^ t[108];
  assign t[89] = t[163] ^ t[171];
  assign t[8] = ~(t[12]);
  assign t[90] = t[172] ^ t[173];
  assign t[91] = t[164] ^ t[174];
  assign t[92] = t[109] ^ t[86];
  assign t[93] = t[109] & t[83];
  assign t[94] = t[110] & t[109];
  assign t[95] = t[25] ? t[175] : t[111];
  assign t[96] = t[25] ? t[176] : t[112];
  assign t[97] = t[110] ^ t[83];
  assign t[98] = t[86] & t[110];
  assign t[99] = t[101] ^ t[67];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind543(x, y);
 input [132:0] x;
 output y;

 wire [448:0] t;
  assign t[0] = t[1] ? t[2] : t[141];
  assign t[100] = t[113] ^ t[101];
  assign t[101] = t[25] ? t[177] : t[114];
  assign t[102] = t[115] ^ t[106];
  assign t[103] = t[116] ^ t[69];
  assign t[104] = t[86] ^ t[94];
  assign t[105] = t[117] ^ t[118];
  assign t[106] = t[119] ^ t[120];
  assign t[107] = t[83] ^ t[94];
  assign t[108] = t[96] ^ t[73];
  assign t[109] = t[121] ^ t[122];
  assign t[10] = t[143] & t[16];
  assign t[110] = t[123] ^ t[122];
  assign t[111] = t[178] ^ t[179];
  assign t[112] = t[180] ^ t[181];
  assign t[113] = t[25] ? t[182] : t[21];
  assign t[114] = t[183] ^ t[184];
  assign t[115] = t[124] ^ t[125];
  assign t[116] = t[56] ^ t[126];
  assign t[117] = t[127] ^ t[128];
  assign t[118] = t[79] ^ t[129];
  assign t[119] = t[79] & t[129];
  assign t[11] = ~(t[17]);
  assign t[120] = t[56] & t[130];
  assign t[121] = t[131] ^ t[132];
  assign t[122] = t[133] ^ t[120];
  assign t[123] = t[134] ^ t[135];
  assign t[124] = t[116] & t[69];
  assign t[125] = t[82] & t[88];
  assign t[126] = t[76] ^ t[136];
  assign t[127] = t[126] & t[67];
  assign t[128] = t[65] & t[81];
  assign t[129] = t[81] ^ t[76];
  assign t[12] = ~(t[143]);
  assign t[130] = t[100] ^ t[137];
  assign t[131] = t[138] ^ t[128];
  assign t[132] = t[62] & t[63];
  assign t[133] = t[58] & t[139];
  assign t[134] = t[140] ^ t[125];
  assign t[135] = t[80] & t[60];
  assign t[136] = t[71] ^ t[67];
  assign t[137] = t[95] ^ t[73];
  assign t[138] = t[81] ^ t[137];
  assign t[139] = t[56] ^ t[108];
  assign t[13] = ~(t[18]);
  assign t[140] = t[82] ^ t[88];
  assign t[141] = (t[185]);
  assign t[142] = (t[186]);
  assign t[143] = (t[187]);
  assign t[144] = (t[188]);
  assign t[145] = (t[189]);
  assign t[146] = (t[190]);
  assign t[147] = (t[191]);
  assign t[148] = (t[192]);
  assign t[149] = (t[193]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[194]);
  assign t[151] = (t[195]);
  assign t[152] = (t[196]);
  assign t[153] = (t[197]);
  assign t[154] = (t[198]);
  assign t[155] = (t[199]);
  assign t[156] = (t[200]);
  assign t[157] = (t[201]);
  assign t[158] = (t[202]);
  assign t[159] = (t[203]);
  assign t[15] = t[19] ? t[144] : t[22];
  assign t[160] = (t[204]);
  assign t[161] = (t[205]);
  assign t[162] = (t[206]);
  assign t[163] = (t[207]);
  assign t[164] = (t[208]);
  assign t[165] = (t[209]);
  assign t[166] = (t[210]);
  assign t[167] = (t[211]);
  assign t[168] = (t[212]);
  assign t[169] = (t[213]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[214]);
  assign t[171] = (t[215]);
  assign t[172] = (t[216]);
  assign t[173] = (t[217]);
  assign t[174] = (t[218]);
  assign t[175] = (t[219]);
  assign t[176] = (t[220]);
  assign t[177] = (t[221]);
  assign t[178] = (t[222]);
  assign t[179] = (t[223]);
  assign t[17] = ~(t[143] & t[24]);
  assign t[180] = (t[224]);
  assign t[181] = (t[225]);
  assign t[182] = (t[226]);
  assign t[183] = (t[227]);
  assign t[184] = (t[228]);
  assign t[185] = t[229] ^ x[2];
  assign t[186] = t[230] ^ x[5];
  assign t[187] = t[231] ^ x[9];
  assign t[188] = t[232] ^ x[12];
  assign t[189] = t[233] ^ x[15];
  assign t[18] = ~(t[25]);
  assign t[190] = t[234] ^ x[18];
  assign t[191] = t[235] ^ x[21];
  assign t[192] = t[236] ^ x[24];
  assign t[193] = t[237] ^ x[27];
  assign t[194] = t[238] ^ x[30];
  assign t[195] = t[239] ^ x[33];
  assign t[196] = t[240] ^ x[36];
  assign t[197] = t[241] ^ x[39];
  assign t[198] = t[242] ^ x[42];
  assign t[199] = t[243] ^ x[45];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[244] ^ x[48];
  assign t[201] = t[245] ^ x[51];
  assign t[202] = t[246] ^ x[54];
  assign t[203] = t[247] ^ x[57];
  assign t[204] = t[248] ^ x[60];
  assign t[205] = t[249] ^ x[63];
  assign t[206] = t[250] ^ x[66];
  assign t[207] = t[251] ^ x[69];
  assign t[208] = t[252] ^ x[72];
  assign t[209] = t[253] ^ x[75];
  assign t[20] = t[28] ^ t[29];
  assign t[210] = t[254] ^ x[78];
  assign t[211] = t[255] ^ x[81];
  assign t[212] = t[256] ^ x[84];
  assign t[213] = t[257] ^ x[87];
  assign t[214] = t[258] ^ x[90];
  assign t[215] = t[259] ^ x[93];
  assign t[216] = t[260] ^ x[96];
  assign t[217] = t[261] ^ x[99];
  assign t[218] = t[262] ^ x[102];
  assign t[219] = t[263] ^ x[105];
  assign t[21] = t[145] ^ t[146];
  assign t[220] = t[264] ^ x[108];
  assign t[221] = t[265] ^ x[111];
  assign t[222] = t[266] ^ x[114];
  assign t[223] = t[267] ^ x[117];
  assign t[224] = t[268] ^ x[120];
  assign t[225] = t[269] ^ x[123];
  assign t[226] = t[270] ^ x[126];
  assign t[227] = t[271] ^ x[129];
  assign t[228] = t[272] ^ x[132];
  assign t[229] = (t[273] & ~t[274]);
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[275] & ~t[276]);
  assign t[231] = (t[277] & ~t[278]);
  assign t[232] = (t[279] & ~t[280]);
  assign t[233] = (t[281] & ~t[282]);
  assign t[234] = (t[283] & ~t[284]);
  assign t[235] = (t[285] & ~t[286]);
  assign t[236] = (t[287] & ~t[288]);
  assign t[237] = (t[289] & ~t[290]);
  assign t[238] = (t[291] & ~t[292]);
  assign t[239] = (t[293] & ~t[294]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[295] & ~t[296]);
  assign t[241] = (t[297] & ~t[298]);
  assign t[242] = (t[299] & ~t[300]);
  assign t[243] = (t[301] & ~t[302]);
  assign t[244] = (t[303] & ~t[304]);
  assign t[245] = (t[305] & ~t[306]);
  assign t[246] = (t[307] & ~t[308]);
  assign t[247] = (t[309] & ~t[310]);
  assign t[248] = (t[311] & ~t[312]);
  assign t[249] = (t[313] & ~t[314]);
  assign t[24] = ~(t[147] | t[34]);
  assign t[250] = (t[315] & ~t[316]);
  assign t[251] = (t[317] & ~t[318]);
  assign t[252] = (t[319] & ~t[320]);
  assign t[253] = (t[321] & ~t[322]);
  assign t[254] = (t[323] & ~t[324]);
  assign t[255] = (t[325] & ~t[326]);
  assign t[256] = (t[327] & ~t[328]);
  assign t[257] = (t[329] & ~t[330]);
  assign t[258] = (t[331] & ~t[332]);
  assign t[259] = (t[333] & ~t[334]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[335] & ~t[336]);
  assign t[261] = (t[337] & ~t[338]);
  assign t[262] = (t[339] & ~t[340]);
  assign t[263] = (t[341] & ~t[342]);
  assign t[264] = (t[343] & ~t[344]);
  assign t[265] = (t[345] & ~t[346]);
  assign t[266] = (t[347] & ~t[348]);
  assign t[267] = (t[349] & ~t[350]);
  assign t[268] = (t[351] & ~t[352]);
  assign t[269] = (t[353] & ~t[354]);
  assign t[26] = ~(t[148] & t[149]);
  assign t[270] = (t[355] & ~t[356]);
  assign t[271] = (t[357] & ~t[358]);
  assign t[272] = (t[359] & ~t[360]);
  assign t[273] = t[361] ^ x[2];
  assign t[274] = t[362] ^ x[1];
  assign t[275] = t[363] ^ x[5];
  assign t[276] = t[364] ^ x[4];
  assign t[277] = t[365] ^ x[9];
  assign t[278] = t[366] ^ x[8];
  assign t[279] = t[367] ^ x[12];
  assign t[27] = ~(t[150] & t[151]);
  assign t[280] = t[368] ^ x[11];
  assign t[281] = t[369] ^ x[15];
  assign t[282] = t[370] ^ x[14];
  assign t[283] = t[371] ^ x[18];
  assign t[284] = t[372] ^ x[17];
  assign t[285] = t[373] ^ x[21];
  assign t[286] = t[374] ^ x[20];
  assign t[287] = t[375] ^ x[24];
  assign t[288] = t[376] ^ x[23];
  assign t[289] = t[377] ^ x[27];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[378] ^ x[26];
  assign t[291] = t[379] ^ x[30];
  assign t[292] = t[380] ^ x[29];
  assign t[293] = t[381] ^ x[33];
  assign t[294] = t[382] ^ x[32];
  assign t[295] = t[383] ^ x[36];
  assign t[296] = t[384] ^ x[35];
  assign t[297] = t[385] ^ x[39];
  assign t[298] = t[386] ^ x[38];
  assign t[299] = t[387] ^ x[42];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[142] : t[5];
  assign t[300] = t[388] ^ x[41];
  assign t[301] = t[389] ^ x[45];
  assign t[302] = t[390] ^ x[44];
  assign t[303] = t[391] ^ x[48];
  assign t[304] = t[392] ^ x[47];
  assign t[305] = t[393] ^ x[51];
  assign t[306] = t[394] ^ x[50];
  assign t[307] = t[395] ^ x[54];
  assign t[308] = t[396] ^ x[53];
  assign t[309] = t[397] ^ x[57];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[398] ^ x[56];
  assign t[311] = t[399] ^ x[60];
  assign t[312] = t[400] ^ x[59];
  assign t[313] = t[401] ^ x[63];
  assign t[314] = t[402] ^ x[62];
  assign t[315] = t[403] ^ x[66];
  assign t[316] = t[404] ^ x[65];
  assign t[317] = t[405] ^ x[69];
  assign t[318] = t[406] ^ x[68];
  assign t[319] = t[407] ^ x[72];
  assign t[31] = ~(t[152] ^ t[153]);
  assign t[320] = t[408] ^ x[71];
  assign t[321] = t[409] ^ x[75];
  assign t[322] = t[410] ^ x[74];
  assign t[323] = t[411] ^ x[78];
  assign t[324] = t[412] ^ x[77];
  assign t[325] = t[413] ^ x[81];
  assign t[326] = t[414] ^ x[80];
  assign t[327] = t[415] ^ x[84];
  assign t[328] = t[416] ^ x[83];
  assign t[329] = t[417] ^ x[87];
  assign t[32] = ~(t[24]);
  assign t[330] = t[418] ^ x[86];
  assign t[331] = t[419] ^ x[90];
  assign t[332] = t[420] ^ x[89];
  assign t[333] = t[421] ^ x[93];
  assign t[334] = t[422] ^ x[92];
  assign t[335] = t[423] ^ x[96];
  assign t[336] = t[424] ^ x[95];
  assign t[337] = t[425] ^ x[99];
  assign t[338] = t[426] ^ x[98];
  assign t[339] = t[427] ^ x[102];
  assign t[33] = ~(t[154] & t[43]);
  assign t[340] = t[428] ^ x[101];
  assign t[341] = t[429] ^ x[105];
  assign t[342] = t[430] ^ x[104];
  assign t[343] = t[431] ^ x[108];
  assign t[344] = t[432] ^ x[107];
  assign t[345] = t[433] ^ x[111];
  assign t[346] = t[434] ^ x[110];
  assign t[347] = t[435] ^ x[114];
  assign t[348] = t[436] ^ x[113];
  assign t[349] = t[437] ^ x[117];
  assign t[34] = ~(t[44] & t[45]);
  assign t[350] = t[438] ^ x[116];
  assign t[351] = t[439] ^ x[120];
  assign t[352] = t[440] ^ x[119];
  assign t[353] = t[441] ^ x[123];
  assign t[354] = t[442] ^ x[122];
  assign t[355] = t[443] ^ x[126];
  assign t[356] = t[444] ^ x[125];
  assign t[357] = t[445] ^ x[129];
  assign t[358] = t[446] ^ x[128];
  assign t[359] = t[447] ^ x[132];
  assign t[35] = ~(t[155]);
  assign t[360] = t[448] ^ x[131];
  assign t[361] = (x[0]);
  assign t[362] = (x[0]);
  assign t[363] = (x[3]);
  assign t[364] = (x[3]);
  assign t[365] = (x[7]);
  assign t[366] = (x[7]);
  assign t[367] = (x[10]);
  assign t[368] = (x[10]);
  assign t[369] = (x[13]);
  assign t[36] = ~(t[143]);
  assign t[370] = (x[13]);
  assign t[371] = (x[16]);
  assign t[372] = (x[16]);
  assign t[373] = (x[19]);
  assign t[374] = (x[19]);
  assign t[375] = (x[22]);
  assign t[376] = (x[22]);
  assign t[377] = (x[25]);
  assign t[378] = (x[25]);
  assign t[379] = (x[28]);
  assign t[37] = t[46] ^ t[47];
  assign t[380] = (x[28]);
  assign t[381] = (x[31]);
  assign t[382] = (x[31]);
  assign t[383] = (x[34]);
  assign t[384] = (x[34]);
  assign t[385] = (x[37]);
  assign t[386] = (x[37]);
  assign t[387] = (x[40]);
  assign t[388] = (x[40]);
  assign t[389] = (x[43]);
  assign t[38] = t[48] ^ t[49];
  assign t[390] = (x[43]);
  assign t[391] = (x[46]);
  assign t[392] = (x[46]);
  assign t[393] = (x[49]);
  assign t[394] = (x[49]);
  assign t[395] = (x[52]);
  assign t[396] = (x[52]);
  assign t[397] = (x[55]);
  assign t[398] = (x[55]);
  assign t[399] = (x[58]);
  assign t[39] = t[50] ^ t[51];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[58]);
  assign t[401] = (x[61]);
  assign t[402] = (x[61]);
  assign t[403] = (x[64]);
  assign t[404] = (x[64]);
  assign t[405] = (x[67]);
  assign t[406] = (x[67]);
  assign t[407] = (x[70]);
  assign t[408] = (x[70]);
  assign t[409] = (x[73]);
  assign t[40] = t[52] ^ t[53];
  assign t[410] = (x[73]);
  assign t[411] = (x[76]);
  assign t[412] = (x[76]);
  assign t[413] = (x[79]);
  assign t[414] = (x[79]);
  assign t[415] = (x[82]);
  assign t[416] = (x[82]);
  assign t[417] = (x[85]);
  assign t[418] = (x[85]);
  assign t[419] = (x[88]);
  assign t[41] = t[156] ^ t[157];
  assign t[420] = (x[88]);
  assign t[421] = (x[91]);
  assign t[422] = (x[91]);
  assign t[423] = (x[94]);
  assign t[424] = (x[94]);
  assign t[425] = (x[97]);
  assign t[426] = (x[97]);
  assign t[427] = (x[100]);
  assign t[428] = (x[100]);
  assign t[429] = (x[103]);
  assign t[42] = t[145] ^ t[54];
  assign t[430] = (x[103]);
  assign t[431] = (x[106]);
  assign t[432] = (x[106]);
  assign t[433] = (x[109]);
  assign t[434] = (x[109]);
  assign t[435] = (x[112]);
  assign t[436] = (x[112]);
  assign t[437] = (x[115]);
  assign t[438] = (x[115]);
  assign t[439] = (x[118]);
  assign t[43] = ~(t[158]);
  assign t[440] = (x[118]);
  assign t[441] = (x[121]);
  assign t[442] = (x[121]);
  assign t[443] = (x[124]);
  assign t[444] = (x[124]);
  assign t[445] = (x[127]);
  assign t[446] = (x[127]);
  assign t[447] = (x[130]);
  assign t[448] = (x[130]);
  assign t[44] = ~(t[159] | t[160]);
  assign t[45] = ~(t[161] | t[162]);
  assign t[46] = t[55] & t[56];
  assign t[47] = t[57] & t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[61] & t[62];
  assign t[4] = ~(t[7]);
  assign t[50] = t[61] & t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[66] & t[67];
  assign t[53] = t[68] & t[69];
  assign t[54] = t[163] ^ t[164];
  assign t[55] = t[68] ^ t[66];
  assign t[56] = t[70] ^ t[71];
  assign t[57] = t[55] ^ t[72];
  assign t[58] = t[71] ^ t[73];
  assign t[59] = t[74] ^ t[75];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[67] ^ t[76];
  assign t[61] = t[77] ^ t[78];
  assign t[62] = t[79] ^ t[80];
  assign t[63] = t[67] ^ t[81];
  assign t[64] = t[66] ^ t[61];
  assign t[65] = t[82] ^ t[58];
  assign t[66] = t[83] ^ t[84];
  assign t[67] = t[25] ? t[165] : t[85];
  assign t[68] = t[86] ^ t[87];
  assign t[69] = t[60] ^ t[88];
  assign t[6] = ~(t[10]);
  assign t[70] = t[25] ? t[166] : t[89];
  assign t[71] = t[25] ? t[167] : t[90];
  assign t[72] = t[59] ^ t[61];
  assign t[73] = t[25] ? t[168] : t[91];
  assign t[74] = t[92] & t[93];
  assign t[75] = t[92] ^ t[94];
  assign t[76] = t[95] ^ t[96];
  assign t[77] = t[97] & t[98];
  assign t[78] = t[97] ^ t[94];
  assign t[79] = t[70] ^ t[73];
  assign t[7] = ~(t[11]);
  assign t[80] = t[76] ^ t[99];
  assign t[81] = t[56] ^ t[100];
  assign t[82] = t[70] ^ t[101];
  assign t[83] = t[102] ^ t[103];
  assign t[84] = t[104] & t[97];
  assign t[85] = t[169] ^ t[170];
  assign t[86] = t[105] ^ t[106];
  assign t[87] = t[107] & t[92];
  assign t[88] = t[100] ^ t[108];
  assign t[89] = t[163] ^ t[171];
  assign t[8] = ~(t[12]);
  assign t[90] = t[172] ^ t[173];
  assign t[91] = t[164] ^ t[174];
  assign t[92] = t[109] ^ t[86];
  assign t[93] = t[109] & t[83];
  assign t[94] = t[110] & t[109];
  assign t[95] = t[25] ? t[175] : t[111];
  assign t[96] = t[25] ? t[176] : t[112];
  assign t[97] = t[110] ^ t[83];
  assign t[98] = t[86] & t[110];
  assign t[99] = t[101] ^ t[67];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind544(x, y);
 input [132:0] x;
 output y;

 wire [449:0] t;
  assign t[0] = t[1] ? t[2] : t[142];
  assign t[100] = t[86] & t[113];
  assign t[101] = t[91] ^ t[78];
  assign t[102] = t[75] ^ t[91];
  assign t[103] = t[115] ^ t[116];
  assign t[104] = t[117] ^ t[118];
  assign t[105] = t[88] ^ t[96];
  assign t[106] = t[119] ^ t[104];
  assign t[107] = t[120] ^ t[121];
  assign t[108] = t[86] ^ t[96];
  assign t[109] = t[165] ^ t[179];
  assign t[10] = t[144] & t[16];
  assign t[110] = t[180] ^ t[181];
  assign t[111] = t[182] ^ t[183];
  assign t[112] = t[122] ^ t[123];
  assign t[113] = t[124] ^ t[123];
  assign t[114] = t[184] ^ t[185];
  assign t[115] = t[125] ^ t[126];
  assign t[116] = t[82] ^ t[127];
  assign t[117] = t[82] & t[127];
  assign t[118] = t[61] & t[128];
  assign t[119] = t[129] ^ t[130];
  assign t[11] = ~(t[17]);
  assign t[120] = t[61] ^ t[131];
  assign t[121] = t[63] ^ t[60];
  assign t[122] = t[132] ^ t[133];
  assign t[123] = t[134] ^ t[118];
  assign t[124] = t[135] ^ t[136];
  assign t[125] = t[131] & t[78];
  assign t[126] = t[85] & t[67];
  assign t[127] = t[67] ^ t[79];
  assign t[128] = t[73] ^ t[137];
  assign t[129] = t[120] & t[121];
  assign t[12] = ~(t[144]);
  assign t[130] = t[102] & t[60];
  assign t[131] = t[79] ^ t[138];
  assign t[132] = t[139] ^ t[126];
  assign t[133] = t[65] & t[84];
  assign t[134] = t[47] & t[140];
  assign t[135] = t[141] ^ t[130];
  assign t[136] = t[83] & t[63];
  assign t[137] = t[98] ^ t[58];
  assign t[138] = t[57] ^ t[78];
  assign t[139] = t[67] ^ t[137];
  assign t[13] = ~(t[18]);
  assign t[140] = t[61] ^ t[74];
  assign t[141] = t[102] ^ t[60];
  assign t[142] = (t[186]);
  assign t[143] = (t[187]);
  assign t[144] = (t[188]);
  assign t[145] = (t[189]);
  assign t[146] = (t[190]);
  assign t[147] = (t[191]);
  assign t[148] = (t[192]);
  assign t[149] = (t[193]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[194]);
  assign t[151] = (t[195]);
  assign t[152] = (t[196]);
  assign t[153] = (t[197]);
  assign t[154] = (t[198]);
  assign t[155] = (t[199]);
  assign t[156] = (t[200]);
  assign t[157] = (t[201]);
  assign t[158] = (t[202]);
  assign t[159] = (t[203]);
  assign t[15] = t[19] ? t[145] : t[22];
  assign t[160] = (t[204]);
  assign t[161] = (t[205]);
  assign t[162] = (t[206]);
  assign t[163] = (t[207]);
  assign t[164] = (t[208]);
  assign t[165] = (t[209]);
  assign t[166] = (t[210]);
  assign t[167] = (t[211]);
  assign t[168] = (t[212]);
  assign t[169] = (t[213]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[214]);
  assign t[171] = (t[215]);
  assign t[172] = (t[216]);
  assign t[173] = (t[217]);
  assign t[174] = (t[218]);
  assign t[175] = (t[219]);
  assign t[176] = (t[220]);
  assign t[177] = (t[221]);
  assign t[178] = (t[222]);
  assign t[179] = (t[223]);
  assign t[17] = ~(t[144] & t[24]);
  assign t[180] = (t[224]);
  assign t[181] = (t[225]);
  assign t[182] = (t[226]);
  assign t[183] = (t[227]);
  assign t[184] = (t[228]);
  assign t[185] = (t[229]);
  assign t[186] = t[230] ^ x[2];
  assign t[187] = t[231] ^ x[5];
  assign t[188] = t[232] ^ x[9];
  assign t[189] = t[233] ^ x[12];
  assign t[18] = ~(t[25]);
  assign t[190] = t[234] ^ x[15];
  assign t[191] = t[235] ^ x[18];
  assign t[192] = t[236] ^ x[21];
  assign t[193] = t[237] ^ x[24];
  assign t[194] = t[238] ^ x[27];
  assign t[195] = t[239] ^ x[30];
  assign t[196] = t[240] ^ x[33];
  assign t[197] = t[241] ^ x[36];
  assign t[198] = t[242] ^ x[39];
  assign t[199] = t[243] ^ x[42];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[244] ^ x[45];
  assign t[201] = t[245] ^ x[48];
  assign t[202] = t[246] ^ x[51];
  assign t[203] = t[247] ^ x[54];
  assign t[204] = t[248] ^ x[57];
  assign t[205] = t[249] ^ x[60];
  assign t[206] = t[250] ^ x[63];
  assign t[207] = t[251] ^ x[66];
  assign t[208] = t[252] ^ x[69];
  assign t[209] = t[253] ^ x[72];
  assign t[20] = t[28] ^ t[29];
  assign t[210] = t[254] ^ x[75];
  assign t[211] = t[255] ^ x[78];
  assign t[212] = t[256] ^ x[81];
  assign t[213] = t[257] ^ x[84];
  assign t[214] = t[258] ^ x[87];
  assign t[215] = t[259] ^ x[90];
  assign t[216] = t[260] ^ x[93];
  assign t[217] = t[261] ^ x[96];
  assign t[218] = t[262] ^ x[99];
  assign t[219] = t[263] ^ x[102];
  assign t[21] = t[146] ^ t[147];
  assign t[220] = t[264] ^ x[105];
  assign t[221] = t[265] ^ x[108];
  assign t[222] = t[266] ^ x[111];
  assign t[223] = t[267] ^ x[114];
  assign t[224] = t[268] ^ x[117];
  assign t[225] = t[269] ^ x[120];
  assign t[226] = t[270] ^ x[123];
  assign t[227] = t[271] ^ x[126];
  assign t[228] = t[272] ^ x[129];
  assign t[229] = t[273] ^ x[132];
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[274] & ~t[275]);
  assign t[231] = (t[276] & ~t[277]);
  assign t[232] = (t[278] & ~t[279]);
  assign t[233] = (t[280] & ~t[281]);
  assign t[234] = (t[282] & ~t[283]);
  assign t[235] = (t[284] & ~t[285]);
  assign t[236] = (t[286] & ~t[287]);
  assign t[237] = (t[288] & ~t[289]);
  assign t[238] = (t[290] & ~t[291]);
  assign t[239] = (t[292] & ~t[293]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[294] & ~t[295]);
  assign t[241] = (t[296] & ~t[297]);
  assign t[242] = (t[298] & ~t[299]);
  assign t[243] = (t[300] & ~t[301]);
  assign t[244] = (t[302] & ~t[303]);
  assign t[245] = (t[304] & ~t[305]);
  assign t[246] = (t[306] & ~t[307]);
  assign t[247] = (t[308] & ~t[309]);
  assign t[248] = (t[310] & ~t[311]);
  assign t[249] = (t[312] & ~t[313]);
  assign t[24] = ~(t[148] | t[34]);
  assign t[250] = (t[314] & ~t[315]);
  assign t[251] = (t[316] & ~t[317]);
  assign t[252] = (t[318] & ~t[319]);
  assign t[253] = (t[320] & ~t[321]);
  assign t[254] = (t[322] & ~t[323]);
  assign t[255] = (t[324] & ~t[325]);
  assign t[256] = (t[326] & ~t[327]);
  assign t[257] = (t[328] & ~t[329]);
  assign t[258] = (t[330] & ~t[331]);
  assign t[259] = (t[332] & ~t[333]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[334] & ~t[335]);
  assign t[261] = (t[336] & ~t[337]);
  assign t[262] = (t[338] & ~t[339]);
  assign t[263] = (t[340] & ~t[341]);
  assign t[264] = (t[342] & ~t[343]);
  assign t[265] = (t[344] & ~t[345]);
  assign t[266] = (t[346] & ~t[347]);
  assign t[267] = (t[348] & ~t[349]);
  assign t[268] = (t[350] & ~t[351]);
  assign t[269] = (t[352] & ~t[353]);
  assign t[26] = ~(t[149] & t[150]);
  assign t[270] = (t[354] & ~t[355]);
  assign t[271] = (t[356] & ~t[357]);
  assign t[272] = (t[358] & ~t[359]);
  assign t[273] = (t[360] & ~t[361]);
  assign t[274] = t[362] ^ x[2];
  assign t[275] = t[363] ^ x[1];
  assign t[276] = t[364] ^ x[5];
  assign t[277] = t[365] ^ x[4];
  assign t[278] = t[366] ^ x[9];
  assign t[279] = t[367] ^ x[8];
  assign t[27] = ~(t[151] & t[152]);
  assign t[280] = t[368] ^ x[12];
  assign t[281] = t[369] ^ x[11];
  assign t[282] = t[370] ^ x[15];
  assign t[283] = t[371] ^ x[14];
  assign t[284] = t[372] ^ x[18];
  assign t[285] = t[373] ^ x[17];
  assign t[286] = t[374] ^ x[21];
  assign t[287] = t[375] ^ x[20];
  assign t[288] = t[376] ^ x[24];
  assign t[289] = t[377] ^ x[23];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[378] ^ x[27];
  assign t[291] = t[379] ^ x[26];
  assign t[292] = t[380] ^ x[30];
  assign t[293] = t[381] ^ x[29];
  assign t[294] = t[382] ^ x[33];
  assign t[295] = t[383] ^ x[32];
  assign t[296] = t[384] ^ x[36];
  assign t[297] = t[385] ^ x[35];
  assign t[298] = t[386] ^ x[39];
  assign t[299] = t[387] ^ x[38];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[143] : t[5];
  assign t[300] = t[388] ^ x[42];
  assign t[301] = t[389] ^ x[41];
  assign t[302] = t[390] ^ x[45];
  assign t[303] = t[391] ^ x[44];
  assign t[304] = t[392] ^ x[48];
  assign t[305] = t[393] ^ x[47];
  assign t[306] = t[394] ^ x[51];
  assign t[307] = t[395] ^ x[50];
  assign t[308] = t[396] ^ x[54];
  assign t[309] = t[397] ^ x[53];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[398] ^ x[57];
  assign t[311] = t[399] ^ x[56];
  assign t[312] = t[400] ^ x[60];
  assign t[313] = t[401] ^ x[59];
  assign t[314] = t[402] ^ x[63];
  assign t[315] = t[403] ^ x[62];
  assign t[316] = t[404] ^ x[66];
  assign t[317] = t[405] ^ x[65];
  assign t[318] = t[406] ^ x[69];
  assign t[319] = t[407] ^ x[68];
  assign t[31] = ~(t[153] ^ t[154]);
  assign t[320] = t[408] ^ x[72];
  assign t[321] = t[409] ^ x[71];
  assign t[322] = t[410] ^ x[75];
  assign t[323] = t[411] ^ x[74];
  assign t[324] = t[412] ^ x[78];
  assign t[325] = t[413] ^ x[77];
  assign t[326] = t[414] ^ x[81];
  assign t[327] = t[415] ^ x[80];
  assign t[328] = t[416] ^ x[84];
  assign t[329] = t[417] ^ x[83];
  assign t[32] = ~(t[24]);
  assign t[330] = t[418] ^ x[87];
  assign t[331] = t[419] ^ x[86];
  assign t[332] = t[420] ^ x[90];
  assign t[333] = t[421] ^ x[89];
  assign t[334] = t[422] ^ x[93];
  assign t[335] = t[423] ^ x[92];
  assign t[336] = t[424] ^ x[96];
  assign t[337] = t[425] ^ x[95];
  assign t[338] = t[426] ^ x[99];
  assign t[339] = t[427] ^ x[98];
  assign t[33] = ~(t[155] & t[43]);
  assign t[340] = t[428] ^ x[102];
  assign t[341] = t[429] ^ x[101];
  assign t[342] = t[430] ^ x[105];
  assign t[343] = t[431] ^ x[104];
  assign t[344] = t[432] ^ x[108];
  assign t[345] = t[433] ^ x[107];
  assign t[346] = t[434] ^ x[111];
  assign t[347] = t[435] ^ x[110];
  assign t[348] = t[436] ^ x[114];
  assign t[349] = t[437] ^ x[113];
  assign t[34] = ~(t[44] & t[45]);
  assign t[350] = t[438] ^ x[117];
  assign t[351] = t[439] ^ x[116];
  assign t[352] = t[440] ^ x[120];
  assign t[353] = t[441] ^ x[119];
  assign t[354] = t[442] ^ x[123];
  assign t[355] = t[443] ^ x[122];
  assign t[356] = t[444] ^ x[126];
  assign t[357] = t[445] ^ x[125];
  assign t[358] = t[446] ^ x[129];
  assign t[359] = t[447] ^ x[128];
  assign t[35] = ~(t[156]);
  assign t[360] = t[448] ^ x[132];
  assign t[361] = t[449] ^ x[131];
  assign t[362] = (x[0]);
  assign t[363] = (x[0]);
  assign t[364] = (x[3]);
  assign t[365] = (x[3]);
  assign t[366] = (x[7]);
  assign t[367] = (x[7]);
  assign t[368] = (x[10]);
  assign t[369] = (x[10]);
  assign t[36] = ~(t[144]);
  assign t[370] = (x[13]);
  assign t[371] = (x[13]);
  assign t[372] = (x[16]);
  assign t[373] = (x[16]);
  assign t[374] = (x[19]);
  assign t[375] = (x[19]);
  assign t[376] = (x[22]);
  assign t[377] = (x[22]);
  assign t[378] = (x[25]);
  assign t[379] = (x[25]);
  assign t[37] = t[46] & t[47];
  assign t[380] = (x[28]);
  assign t[381] = (x[28]);
  assign t[382] = (x[31]);
  assign t[383] = (x[31]);
  assign t[384] = (x[34]);
  assign t[385] = (x[34]);
  assign t[386] = (x[37]);
  assign t[387] = (x[37]);
  assign t[388] = (x[40]);
  assign t[389] = (x[40]);
  assign t[38] = t[48] ^ t[49];
  assign t[390] = (x[43]);
  assign t[391] = (x[43]);
  assign t[392] = (x[46]);
  assign t[393] = (x[46]);
  assign t[394] = (x[49]);
  assign t[395] = (x[49]);
  assign t[396] = (x[52]);
  assign t[397] = (x[52]);
  assign t[398] = (x[55]);
  assign t[399] = (x[55]);
  assign t[39] = t[50] ^ t[51];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[58]);
  assign t[401] = (x[58]);
  assign t[402] = (x[61]);
  assign t[403] = (x[61]);
  assign t[404] = (x[64]);
  assign t[405] = (x[64]);
  assign t[406] = (x[67]);
  assign t[407] = (x[67]);
  assign t[408] = (x[70]);
  assign t[409] = (x[70]);
  assign t[40] = t[52] ^ t[53];
  assign t[410] = (x[73]);
  assign t[411] = (x[73]);
  assign t[412] = (x[76]);
  assign t[413] = (x[76]);
  assign t[414] = (x[79]);
  assign t[415] = (x[79]);
  assign t[416] = (x[82]);
  assign t[417] = (x[82]);
  assign t[418] = (x[85]);
  assign t[419] = (x[85]);
  assign t[41] = t[157] ^ t[158];
  assign t[420] = (x[88]);
  assign t[421] = (x[88]);
  assign t[422] = (x[91]);
  assign t[423] = (x[91]);
  assign t[424] = (x[94]);
  assign t[425] = (x[94]);
  assign t[426] = (x[97]);
  assign t[427] = (x[97]);
  assign t[428] = (x[100]);
  assign t[429] = (x[100]);
  assign t[42] = t[146] ^ t[54];
  assign t[430] = (x[103]);
  assign t[431] = (x[103]);
  assign t[432] = (x[106]);
  assign t[433] = (x[106]);
  assign t[434] = (x[109]);
  assign t[435] = (x[109]);
  assign t[436] = (x[112]);
  assign t[437] = (x[112]);
  assign t[438] = (x[115]);
  assign t[439] = (x[115]);
  assign t[43] = ~(t[159]);
  assign t[440] = (x[118]);
  assign t[441] = (x[118]);
  assign t[442] = (x[121]);
  assign t[443] = (x[121]);
  assign t[444] = (x[124]);
  assign t[445] = (x[124]);
  assign t[446] = (x[127]);
  assign t[447] = (x[127]);
  assign t[448] = (x[130]);
  assign t[449] = (x[130]);
  assign t[44] = ~(t[160] | t[161]);
  assign t[45] = ~(t[162] | t[163]);
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[57] ^ t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[55] & t[61];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] & t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[66] & t[67];
  assign t[53] = t[68] ^ t[69];
  assign t[54] = t[164] ^ t[165];
  assign t[55] = t[70] ^ t[71];
  assign t[56] = t[62] ^ t[64];
  assign t[57] = t[25] ? t[166] : t[21];
  assign t[58] = t[25] ? t[167] : t[72];
  assign t[59] = t[70] ^ t[62];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[73] ^ t[74];
  assign t[61] = t[75] ^ t[57];
  assign t[62] = t[76] ^ t[77];
  assign t[63] = t[78] ^ t[79];
  assign t[64] = t[80] ^ t[81];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[71] ^ t[64];
  assign t[67] = t[61] ^ t[73];
  assign t[68] = t[64] & t[84];
  assign t[69] = t[66] & t[85];
  assign t[6] = ~(t[10]);
  assign t[70] = t[86] ^ t[87];
  assign t[71] = t[88] ^ t[89];
  assign t[72] = t[168] ^ t[169];
  assign t[73] = t[90] ^ t[91];
  assign t[74] = t[92] ^ t[58];
  assign t[75] = t[25] ? t[170] : t[93];
  assign t[76] = t[94] & t[95];
  assign t[77] = t[94] ^ t[96];
  assign t[78] = t[25] ? t[171] : t[97];
  assign t[79] = t[98] ^ t[92];
  assign t[7] = ~(t[11]);
  assign t[80] = t[99] & t[100];
  assign t[81] = t[99] ^ t[96];
  assign t[82] = t[75] ^ t[58];
  assign t[83] = t[79] ^ t[101];
  assign t[84] = t[78] ^ t[67];
  assign t[85] = t[102] ^ t[47];
  assign t[86] = t[103] ^ t[104];
  assign t[87] = t[105] & t[94];
  assign t[88] = t[106] ^ t[107];
  assign t[89] = t[108] & t[99];
  assign t[8] = ~(t[12]);
  assign t[90] = t[25] ? t[172] : t[109];
  assign t[91] = t[25] ? t[173] : t[110];
  assign t[92] = t[25] ? t[174] : t[111];
  assign t[93] = t[164] ^ t[175];
  assign t[94] = t[112] ^ t[86];
  assign t[95] = t[112] & t[88];
  assign t[96] = t[113] & t[112];
  assign t[97] = t[176] ^ t[177];
  assign t[98] = t[25] ? t[178] : t[114];
  assign t[99] = t[113] ^ t[88];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind545(x, y);
 input [132:0] x;
 output y;

 wire [449:0] t;
  assign t[0] = t[1] ? t[2] : t[142];
  assign t[100] = t[86] & t[113];
  assign t[101] = t[91] ^ t[78];
  assign t[102] = t[75] ^ t[91];
  assign t[103] = t[115] ^ t[116];
  assign t[104] = t[117] ^ t[118];
  assign t[105] = t[88] ^ t[96];
  assign t[106] = t[119] ^ t[104];
  assign t[107] = t[120] ^ t[121];
  assign t[108] = t[86] ^ t[96];
  assign t[109] = t[165] ^ t[179];
  assign t[10] = t[144] & t[16];
  assign t[110] = t[180] ^ t[181];
  assign t[111] = t[182] ^ t[183];
  assign t[112] = t[122] ^ t[123];
  assign t[113] = t[124] ^ t[123];
  assign t[114] = t[184] ^ t[185];
  assign t[115] = t[125] ^ t[126];
  assign t[116] = t[82] ^ t[127];
  assign t[117] = t[82] & t[127];
  assign t[118] = t[61] & t[128];
  assign t[119] = t[129] ^ t[130];
  assign t[11] = ~(t[17]);
  assign t[120] = t[61] ^ t[131];
  assign t[121] = t[63] ^ t[60];
  assign t[122] = t[132] ^ t[133];
  assign t[123] = t[134] ^ t[118];
  assign t[124] = t[135] ^ t[136];
  assign t[125] = t[131] & t[78];
  assign t[126] = t[85] & t[67];
  assign t[127] = t[67] ^ t[79];
  assign t[128] = t[73] ^ t[137];
  assign t[129] = t[120] & t[121];
  assign t[12] = ~(t[144]);
  assign t[130] = t[102] & t[60];
  assign t[131] = t[79] ^ t[138];
  assign t[132] = t[139] ^ t[126];
  assign t[133] = t[65] & t[84];
  assign t[134] = t[47] & t[140];
  assign t[135] = t[141] ^ t[130];
  assign t[136] = t[83] & t[63];
  assign t[137] = t[98] ^ t[58];
  assign t[138] = t[57] ^ t[78];
  assign t[139] = t[67] ^ t[137];
  assign t[13] = ~(t[18]);
  assign t[140] = t[61] ^ t[74];
  assign t[141] = t[102] ^ t[60];
  assign t[142] = (t[186]);
  assign t[143] = (t[187]);
  assign t[144] = (t[188]);
  assign t[145] = (t[189]);
  assign t[146] = (t[190]);
  assign t[147] = (t[191]);
  assign t[148] = (t[192]);
  assign t[149] = (t[193]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[194]);
  assign t[151] = (t[195]);
  assign t[152] = (t[196]);
  assign t[153] = (t[197]);
  assign t[154] = (t[198]);
  assign t[155] = (t[199]);
  assign t[156] = (t[200]);
  assign t[157] = (t[201]);
  assign t[158] = (t[202]);
  assign t[159] = (t[203]);
  assign t[15] = t[19] ? t[145] : t[22];
  assign t[160] = (t[204]);
  assign t[161] = (t[205]);
  assign t[162] = (t[206]);
  assign t[163] = (t[207]);
  assign t[164] = (t[208]);
  assign t[165] = (t[209]);
  assign t[166] = (t[210]);
  assign t[167] = (t[211]);
  assign t[168] = (t[212]);
  assign t[169] = (t[213]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[214]);
  assign t[171] = (t[215]);
  assign t[172] = (t[216]);
  assign t[173] = (t[217]);
  assign t[174] = (t[218]);
  assign t[175] = (t[219]);
  assign t[176] = (t[220]);
  assign t[177] = (t[221]);
  assign t[178] = (t[222]);
  assign t[179] = (t[223]);
  assign t[17] = ~(t[144] & t[24]);
  assign t[180] = (t[224]);
  assign t[181] = (t[225]);
  assign t[182] = (t[226]);
  assign t[183] = (t[227]);
  assign t[184] = (t[228]);
  assign t[185] = (t[229]);
  assign t[186] = t[230] ^ x[2];
  assign t[187] = t[231] ^ x[5];
  assign t[188] = t[232] ^ x[9];
  assign t[189] = t[233] ^ x[12];
  assign t[18] = ~(t[25]);
  assign t[190] = t[234] ^ x[15];
  assign t[191] = t[235] ^ x[18];
  assign t[192] = t[236] ^ x[21];
  assign t[193] = t[237] ^ x[24];
  assign t[194] = t[238] ^ x[27];
  assign t[195] = t[239] ^ x[30];
  assign t[196] = t[240] ^ x[33];
  assign t[197] = t[241] ^ x[36];
  assign t[198] = t[242] ^ x[39];
  assign t[199] = t[243] ^ x[42];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[244] ^ x[45];
  assign t[201] = t[245] ^ x[48];
  assign t[202] = t[246] ^ x[51];
  assign t[203] = t[247] ^ x[54];
  assign t[204] = t[248] ^ x[57];
  assign t[205] = t[249] ^ x[60];
  assign t[206] = t[250] ^ x[63];
  assign t[207] = t[251] ^ x[66];
  assign t[208] = t[252] ^ x[69];
  assign t[209] = t[253] ^ x[72];
  assign t[20] = t[28] ^ t[29];
  assign t[210] = t[254] ^ x[75];
  assign t[211] = t[255] ^ x[78];
  assign t[212] = t[256] ^ x[81];
  assign t[213] = t[257] ^ x[84];
  assign t[214] = t[258] ^ x[87];
  assign t[215] = t[259] ^ x[90];
  assign t[216] = t[260] ^ x[93];
  assign t[217] = t[261] ^ x[96];
  assign t[218] = t[262] ^ x[99];
  assign t[219] = t[263] ^ x[102];
  assign t[21] = t[146] ^ t[147];
  assign t[220] = t[264] ^ x[105];
  assign t[221] = t[265] ^ x[108];
  assign t[222] = t[266] ^ x[111];
  assign t[223] = t[267] ^ x[114];
  assign t[224] = t[268] ^ x[117];
  assign t[225] = t[269] ^ x[120];
  assign t[226] = t[270] ^ x[123];
  assign t[227] = t[271] ^ x[126];
  assign t[228] = t[272] ^ x[129];
  assign t[229] = t[273] ^ x[132];
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[274] & ~t[275]);
  assign t[231] = (t[276] & ~t[277]);
  assign t[232] = (t[278] & ~t[279]);
  assign t[233] = (t[280] & ~t[281]);
  assign t[234] = (t[282] & ~t[283]);
  assign t[235] = (t[284] & ~t[285]);
  assign t[236] = (t[286] & ~t[287]);
  assign t[237] = (t[288] & ~t[289]);
  assign t[238] = (t[290] & ~t[291]);
  assign t[239] = (t[292] & ~t[293]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[294] & ~t[295]);
  assign t[241] = (t[296] & ~t[297]);
  assign t[242] = (t[298] & ~t[299]);
  assign t[243] = (t[300] & ~t[301]);
  assign t[244] = (t[302] & ~t[303]);
  assign t[245] = (t[304] & ~t[305]);
  assign t[246] = (t[306] & ~t[307]);
  assign t[247] = (t[308] & ~t[309]);
  assign t[248] = (t[310] & ~t[311]);
  assign t[249] = (t[312] & ~t[313]);
  assign t[24] = ~(t[148] | t[34]);
  assign t[250] = (t[314] & ~t[315]);
  assign t[251] = (t[316] & ~t[317]);
  assign t[252] = (t[318] & ~t[319]);
  assign t[253] = (t[320] & ~t[321]);
  assign t[254] = (t[322] & ~t[323]);
  assign t[255] = (t[324] & ~t[325]);
  assign t[256] = (t[326] & ~t[327]);
  assign t[257] = (t[328] & ~t[329]);
  assign t[258] = (t[330] & ~t[331]);
  assign t[259] = (t[332] & ~t[333]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[334] & ~t[335]);
  assign t[261] = (t[336] & ~t[337]);
  assign t[262] = (t[338] & ~t[339]);
  assign t[263] = (t[340] & ~t[341]);
  assign t[264] = (t[342] & ~t[343]);
  assign t[265] = (t[344] & ~t[345]);
  assign t[266] = (t[346] & ~t[347]);
  assign t[267] = (t[348] & ~t[349]);
  assign t[268] = (t[350] & ~t[351]);
  assign t[269] = (t[352] & ~t[353]);
  assign t[26] = ~(t[149] & t[150]);
  assign t[270] = (t[354] & ~t[355]);
  assign t[271] = (t[356] & ~t[357]);
  assign t[272] = (t[358] & ~t[359]);
  assign t[273] = (t[360] & ~t[361]);
  assign t[274] = t[362] ^ x[2];
  assign t[275] = t[363] ^ x[1];
  assign t[276] = t[364] ^ x[5];
  assign t[277] = t[365] ^ x[4];
  assign t[278] = t[366] ^ x[9];
  assign t[279] = t[367] ^ x[8];
  assign t[27] = ~(t[151] & t[152]);
  assign t[280] = t[368] ^ x[12];
  assign t[281] = t[369] ^ x[11];
  assign t[282] = t[370] ^ x[15];
  assign t[283] = t[371] ^ x[14];
  assign t[284] = t[372] ^ x[18];
  assign t[285] = t[373] ^ x[17];
  assign t[286] = t[374] ^ x[21];
  assign t[287] = t[375] ^ x[20];
  assign t[288] = t[376] ^ x[24];
  assign t[289] = t[377] ^ x[23];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[378] ^ x[27];
  assign t[291] = t[379] ^ x[26];
  assign t[292] = t[380] ^ x[30];
  assign t[293] = t[381] ^ x[29];
  assign t[294] = t[382] ^ x[33];
  assign t[295] = t[383] ^ x[32];
  assign t[296] = t[384] ^ x[36];
  assign t[297] = t[385] ^ x[35];
  assign t[298] = t[386] ^ x[39];
  assign t[299] = t[387] ^ x[38];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[143] : t[5];
  assign t[300] = t[388] ^ x[42];
  assign t[301] = t[389] ^ x[41];
  assign t[302] = t[390] ^ x[45];
  assign t[303] = t[391] ^ x[44];
  assign t[304] = t[392] ^ x[48];
  assign t[305] = t[393] ^ x[47];
  assign t[306] = t[394] ^ x[51];
  assign t[307] = t[395] ^ x[50];
  assign t[308] = t[396] ^ x[54];
  assign t[309] = t[397] ^ x[53];
  assign t[30] = t[41] ^ t[42];
  assign t[310] = t[398] ^ x[57];
  assign t[311] = t[399] ^ x[56];
  assign t[312] = t[400] ^ x[60];
  assign t[313] = t[401] ^ x[59];
  assign t[314] = t[402] ^ x[63];
  assign t[315] = t[403] ^ x[62];
  assign t[316] = t[404] ^ x[66];
  assign t[317] = t[405] ^ x[65];
  assign t[318] = t[406] ^ x[69];
  assign t[319] = t[407] ^ x[68];
  assign t[31] = ~(t[153] ^ t[154]);
  assign t[320] = t[408] ^ x[72];
  assign t[321] = t[409] ^ x[71];
  assign t[322] = t[410] ^ x[75];
  assign t[323] = t[411] ^ x[74];
  assign t[324] = t[412] ^ x[78];
  assign t[325] = t[413] ^ x[77];
  assign t[326] = t[414] ^ x[81];
  assign t[327] = t[415] ^ x[80];
  assign t[328] = t[416] ^ x[84];
  assign t[329] = t[417] ^ x[83];
  assign t[32] = ~(t[24]);
  assign t[330] = t[418] ^ x[87];
  assign t[331] = t[419] ^ x[86];
  assign t[332] = t[420] ^ x[90];
  assign t[333] = t[421] ^ x[89];
  assign t[334] = t[422] ^ x[93];
  assign t[335] = t[423] ^ x[92];
  assign t[336] = t[424] ^ x[96];
  assign t[337] = t[425] ^ x[95];
  assign t[338] = t[426] ^ x[99];
  assign t[339] = t[427] ^ x[98];
  assign t[33] = ~(t[155] & t[43]);
  assign t[340] = t[428] ^ x[102];
  assign t[341] = t[429] ^ x[101];
  assign t[342] = t[430] ^ x[105];
  assign t[343] = t[431] ^ x[104];
  assign t[344] = t[432] ^ x[108];
  assign t[345] = t[433] ^ x[107];
  assign t[346] = t[434] ^ x[111];
  assign t[347] = t[435] ^ x[110];
  assign t[348] = t[436] ^ x[114];
  assign t[349] = t[437] ^ x[113];
  assign t[34] = ~(t[44] & t[45]);
  assign t[350] = t[438] ^ x[117];
  assign t[351] = t[439] ^ x[116];
  assign t[352] = t[440] ^ x[120];
  assign t[353] = t[441] ^ x[119];
  assign t[354] = t[442] ^ x[123];
  assign t[355] = t[443] ^ x[122];
  assign t[356] = t[444] ^ x[126];
  assign t[357] = t[445] ^ x[125];
  assign t[358] = t[446] ^ x[129];
  assign t[359] = t[447] ^ x[128];
  assign t[35] = ~(t[156]);
  assign t[360] = t[448] ^ x[132];
  assign t[361] = t[449] ^ x[131];
  assign t[362] = (x[0]);
  assign t[363] = (x[0]);
  assign t[364] = (x[3]);
  assign t[365] = (x[3]);
  assign t[366] = (x[7]);
  assign t[367] = (x[7]);
  assign t[368] = (x[10]);
  assign t[369] = (x[10]);
  assign t[36] = ~(t[144]);
  assign t[370] = (x[13]);
  assign t[371] = (x[13]);
  assign t[372] = (x[16]);
  assign t[373] = (x[16]);
  assign t[374] = (x[19]);
  assign t[375] = (x[19]);
  assign t[376] = (x[22]);
  assign t[377] = (x[22]);
  assign t[378] = (x[25]);
  assign t[379] = (x[25]);
  assign t[37] = t[46] & t[47];
  assign t[380] = (x[28]);
  assign t[381] = (x[28]);
  assign t[382] = (x[31]);
  assign t[383] = (x[31]);
  assign t[384] = (x[34]);
  assign t[385] = (x[34]);
  assign t[386] = (x[37]);
  assign t[387] = (x[37]);
  assign t[388] = (x[40]);
  assign t[389] = (x[40]);
  assign t[38] = t[48] ^ t[49];
  assign t[390] = (x[43]);
  assign t[391] = (x[43]);
  assign t[392] = (x[46]);
  assign t[393] = (x[46]);
  assign t[394] = (x[49]);
  assign t[395] = (x[49]);
  assign t[396] = (x[52]);
  assign t[397] = (x[52]);
  assign t[398] = (x[55]);
  assign t[399] = (x[55]);
  assign t[39] = t[50] ^ t[51];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[58]);
  assign t[401] = (x[58]);
  assign t[402] = (x[61]);
  assign t[403] = (x[61]);
  assign t[404] = (x[64]);
  assign t[405] = (x[64]);
  assign t[406] = (x[67]);
  assign t[407] = (x[67]);
  assign t[408] = (x[70]);
  assign t[409] = (x[70]);
  assign t[40] = t[52] ^ t[53];
  assign t[410] = (x[73]);
  assign t[411] = (x[73]);
  assign t[412] = (x[76]);
  assign t[413] = (x[76]);
  assign t[414] = (x[79]);
  assign t[415] = (x[79]);
  assign t[416] = (x[82]);
  assign t[417] = (x[82]);
  assign t[418] = (x[85]);
  assign t[419] = (x[85]);
  assign t[41] = t[157] ^ t[158];
  assign t[420] = (x[88]);
  assign t[421] = (x[88]);
  assign t[422] = (x[91]);
  assign t[423] = (x[91]);
  assign t[424] = (x[94]);
  assign t[425] = (x[94]);
  assign t[426] = (x[97]);
  assign t[427] = (x[97]);
  assign t[428] = (x[100]);
  assign t[429] = (x[100]);
  assign t[42] = t[146] ^ t[54];
  assign t[430] = (x[103]);
  assign t[431] = (x[103]);
  assign t[432] = (x[106]);
  assign t[433] = (x[106]);
  assign t[434] = (x[109]);
  assign t[435] = (x[109]);
  assign t[436] = (x[112]);
  assign t[437] = (x[112]);
  assign t[438] = (x[115]);
  assign t[439] = (x[115]);
  assign t[43] = ~(t[159]);
  assign t[440] = (x[118]);
  assign t[441] = (x[118]);
  assign t[442] = (x[121]);
  assign t[443] = (x[121]);
  assign t[444] = (x[124]);
  assign t[445] = (x[124]);
  assign t[446] = (x[127]);
  assign t[447] = (x[127]);
  assign t[448] = (x[130]);
  assign t[449] = (x[130]);
  assign t[44] = ~(t[160] | t[161]);
  assign t[45] = ~(t[162] | t[163]);
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[57] ^ t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[55] & t[61];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] & t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[66] & t[67];
  assign t[53] = t[68] ^ t[69];
  assign t[54] = t[164] ^ t[165];
  assign t[55] = t[70] ^ t[71];
  assign t[56] = t[62] ^ t[64];
  assign t[57] = t[25] ? t[166] : t[21];
  assign t[58] = t[25] ? t[167] : t[72];
  assign t[59] = t[70] ^ t[62];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[73] ^ t[74];
  assign t[61] = t[75] ^ t[57];
  assign t[62] = t[76] ^ t[77];
  assign t[63] = t[78] ^ t[79];
  assign t[64] = t[80] ^ t[81];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[71] ^ t[64];
  assign t[67] = t[61] ^ t[73];
  assign t[68] = t[64] & t[84];
  assign t[69] = t[66] & t[85];
  assign t[6] = ~(t[10]);
  assign t[70] = t[86] ^ t[87];
  assign t[71] = t[88] ^ t[89];
  assign t[72] = t[168] ^ t[169];
  assign t[73] = t[90] ^ t[91];
  assign t[74] = t[92] ^ t[58];
  assign t[75] = t[25] ? t[170] : t[93];
  assign t[76] = t[94] & t[95];
  assign t[77] = t[94] ^ t[96];
  assign t[78] = t[25] ? t[171] : t[97];
  assign t[79] = t[98] ^ t[92];
  assign t[7] = ~(t[11]);
  assign t[80] = t[99] & t[100];
  assign t[81] = t[99] ^ t[96];
  assign t[82] = t[75] ^ t[58];
  assign t[83] = t[79] ^ t[101];
  assign t[84] = t[78] ^ t[67];
  assign t[85] = t[102] ^ t[47];
  assign t[86] = t[103] ^ t[104];
  assign t[87] = t[105] & t[94];
  assign t[88] = t[106] ^ t[107];
  assign t[89] = t[108] & t[99];
  assign t[8] = ~(t[12]);
  assign t[90] = t[25] ? t[172] : t[109];
  assign t[91] = t[25] ? t[173] : t[110];
  assign t[92] = t[25] ? t[174] : t[111];
  assign t[93] = t[164] ^ t[175];
  assign t[94] = t[112] ^ t[86];
  assign t[95] = t[112] & t[88];
  assign t[96] = t[113] & t[112];
  assign t[97] = t[176] ^ t[177];
  assign t[98] = t[25] ? t[178] : t[114];
  assign t[99] = t[113] ^ t[88];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind546(x, y);
 input [129:0] x;
 output y;

 wire [439:0] t;
  assign t[0] = t[1] ? t[2] : t[139];
  assign t[100] = t[25] ? t[176] : t[112];
  assign t[101] = t[155] ^ t[177];
  assign t[102] = t[113] ^ t[114];
  assign t[103] = t[115] ^ t[114];
  assign t[104] = t[178] ^ t[179];
  assign t[105] = t[116] ^ t[117];
  assign t[106] = t[46] ^ t[57];
  assign t[107] = t[46] & t[57];
  assign t[108] = t[66] & t[65];
  assign t[109] = t[118] ^ t[94];
  assign t[10] = t[141] & t[16];
  assign t[110] = t[61] ^ t[119];
  assign t[111] = t[76] ^ t[87];
  assign t[112] = t[180] ^ t[181];
  assign t[113] = t[120] ^ t[121];
  assign t[114] = t[122] ^ t[108];
  assign t[115] = t[123] ^ t[124];
  assign t[116] = t[78] & t[81];
  assign t[117] = t[125] & t[73];
  assign t[118] = t[126] ^ t[127];
  assign t[119] = t[128] ^ t[129];
  assign t[11] = ~(t[17]);
  assign t[120] = t[130] ^ t[117];
  assign t[121] = t[131] & t[132];
  assign t[122] = t[133] & t[134];
  assign t[123] = t[135] ^ t[127];
  assign t[124] = t[136] & t[128];
  assign t[125] = t[59] ^ t[133];
  assign t[126] = t[61] & t[119];
  assign t[127] = t[59] & t[129];
  assign t[128] = t[81] ^ t[74];
  assign t[129] = t[82] ^ t[137];
  assign t[12] = ~(t[141]);
  assign t[130] = t[73] ^ t[83];
  assign t[131] = t[46] ^ t[136];
  assign t[132] = t[81] ^ t[73];
  assign t[133] = t[84] ^ t[56];
  assign t[134] = t[66] ^ t[137];
  assign t[135] = t[59] ^ t[129];
  assign t[136] = t[74] ^ t[138];
  assign t[137] = t[91] ^ t[56];
  assign t[138] = t[75] ^ t[81];
  assign t[139] = (t[182]);
  assign t[13] = ~(t[18]);
  assign t[140] = (t[183]);
  assign t[141] = (t[184]);
  assign t[142] = (t[185]);
  assign t[143] = (t[186]);
  assign t[144] = (t[187]);
  assign t[145] = (t[188]);
  assign t[146] = (t[189]);
  assign t[147] = (t[190]);
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[19] ? t[142] : t[22];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[141] & t[24]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = t[225] ^ x[2];
  assign t[183] = t[226] ^ x[5];
  assign t[184] = t[227] ^ x[9];
  assign t[185] = t[228] ^ x[12];
  assign t[186] = t[229] ^ x[15];
  assign t[187] = t[230] ^ x[18];
  assign t[188] = t[231] ^ x[21];
  assign t[189] = t[232] ^ x[24];
  assign t[18] = ~(t[25]);
  assign t[190] = t[233] ^ x[27];
  assign t[191] = t[234] ^ x[30];
  assign t[192] = t[235] ^ x[33];
  assign t[193] = t[236] ^ x[36];
  assign t[194] = t[237] ^ x[39];
  assign t[195] = t[238] ^ x[42];
  assign t[196] = t[239] ^ x[45];
  assign t[197] = t[240] ^ x[48];
  assign t[198] = t[241] ^ x[51];
  assign t[199] = t[242] ^ x[54];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[57];
  assign t[201] = t[244] ^ x[60];
  assign t[202] = t[245] ^ x[63];
  assign t[203] = t[246] ^ x[66];
  assign t[204] = t[247] ^ x[69];
  assign t[205] = t[248] ^ x[72];
  assign t[206] = t[249] ^ x[75];
  assign t[207] = t[250] ^ x[78];
  assign t[208] = t[251] ^ x[81];
  assign t[209] = t[252] ^ x[84];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[253] ^ x[87];
  assign t[211] = t[254] ^ x[90];
  assign t[212] = t[255] ^ x[93];
  assign t[213] = t[256] ^ x[96];
  assign t[214] = t[257] ^ x[99];
  assign t[215] = t[258] ^ x[102];
  assign t[216] = t[259] ^ x[105];
  assign t[217] = t[260] ^ x[108];
  assign t[218] = t[261] ^ x[111];
  assign t[219] = t[262] ^ x[114];
  assign t[21] = t[143] ^ t[144];
  assign t[220] = t[263] ^ x[117];
  assign t[221] = t[264] ^ x[120];
  assign t[222] = t[265] ^ x[123];
  assign t[223] = t[266] ^ x[126];
  assign t[224] = t[267] ^ x[129];
  assign t[225] = (t[268] & ~t[269]);
  assign t[226] = (t[270] & ~t[271]);
  assign t[227] = (t[272] & ~t[273]);
  assign t[228] = (t[274] & ~t[275]);
  assign t[229] = (t[276] & ~t[277]);
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[278] & ~t[279]);
  assign t[231] = (t[280] & ~t[281]);
  assign t[232] = (t[282] & ~t[283]);
  assign t[233] = (t[284] & ~t[285]);
  assign t[234] = (t[286] & ~t[287]);
  assign t[235] = (t[288] & ~t[289]);
  assign t[236] = (t[290] & ~t[291]);
  assign t[237] = (t[292] & ~t[293]);
  assign t[238] = (t[294] & ~t[295]);
  assign t[239] = (t[296] & ~t[297]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[298] & ~t[299]);
  assign t[241] = (t[300] & ~t[301]);
  assign t[242] = (t[302] & ~t[303]);
  assign t[243] = (t[304] & ~t[305]);
  assign t[244] = (t[306] & ~t[307]);
  assign t[245] = (t[308] & ~t[309]);
  assign t[246] = (t[310] & ~t[311]);
  assign t[247] = (t[312] & ~t[313]);
  assign t[248] = (t[314] & ~t[315]);
  assign t[249] = (t[316] & ~t[317]);
  assign t[24] = ~(t[145] | t[34]);
  assign t[250] = (t[318] & ~t[319]);
  assign t[251] = (t[320] & ~t[321]);
  assign t[252] = (t[322] & ~t[323]);
  assign t[253] = (t[324] & ~t[325]);
  assign t[254] = (t[326] & ~t[327]);
  assign t[255] = (t[328] & ~t[329]);
  assign t[256] = (t[330] & ~t[331]);
  assign t[257] = (t[332] & ~t[333]);
  assign t[258] = (t[334] & ~t[335]);
  assign t[259] = (t[336] & ~t[337]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[338] & ~t[339]);
  assign t[261] = (t[340] & ~t[341]);
  assign t[262] = (t[342] & ~t[343]);
  assign t[263] = (t[344] & ~t[345]);
  assign t[264] = (t[346] & ~t[347]);
  assign t[265] = (t[348] & ~t[349]);
  assign t[266] = (t[350] & ~t[351]);
  assign t[267] = (t[352] & ~t[353]);
  assign t[268] = t[354] ^ x[2];
  assign t[269] = t[355] ^ x[1];
  assign t[26] = ~(t[146] & t[147]);
  assign t[270] = t[356] ^ x[5];
  assign t[271] = t[357] ^ x[4];
  assign t[272] = t[358] ^ x[9];
  assign t[273] = t[359] ^ x[8];
  assign t[274] = t[360] ^ x[12];
  assign t[275] = t[361] ^ x[11];
  assign t[276] = t[362] ^ x[15];
  assign t[277] = t[363] ^ x[14];
  assign t[278] = t[364] ^ x[18];
  assign t[279] = t[365] ^ x[17];
  assign t[27] = ~(t[148] & t[149]);
  assign t[280] = t[366] ^ x[21];
  assign t[281] = t[367] ^ x[20];
  assign t[282] = t[368] ^ x[24];
  assign t[283] = t[369] ^ x[23];
  assign t[284] = t[370] ^ x[27];
  assign t[285] = t[371] ^ x[26];
  assign t[286] = t[372] ^ x[30];
  assign t[287] = t[373] ^ x[29];
  assign t[288] = t[374] ^ x[33];
  assign t[289] = t[375] ^ x[32];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[376] ^ x[36];
  assign t[291] = t[377] ^ x[35];
  assign t[292] = t[378] ^ x[39];
  assign t[293] = t[379] ^ x[38];
  assign t[294] = t[380] ^ x[42];
  assign t[295] = t[381] ^ x[41];
  assign t[296] = t[382] ^ x[45];
  assign t[297] = t[383] ^ x[44];
  assign t[298] = t[384] ^ x[48];
  assign t[299] = t[385] ^ x[47];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[140] : t[5];
  assign t[300] = t[386] ^ x[51];
  assign t[301] = t[387] ^ x[50];
  assign t[302] = t[388] ^ x[54];
  assign t[303] = t[389] ^ x[53];
  assign t[304] = t[390] ^ x[57];
  assign t[305] = t[391] ^ x[56];
  assign t[306] = t[392] ^ x[60];
  assign t[307] = t[393] ^ x[59];
  assign t[308] = t[394] ^ x[63];
  assign t[309] = t[395] ^ x[62];
  assign t[30] = t[150] ^ t[41];
  assign t[310] = t[396] ^ x[66];
  assign t[311] = t[397] ^ x[65];
  assign t[312] = t[398] ^ x[69];
  assign t[313] = t[399] ^ x[68];
  assign t[314] = t[400] ^ x[72];
  assign t[315] = t[401] ^ x[71];
  assign t[316] = t[402] ^ x[75];
  assign t[317] = t[403] ^ x[74];
  assign t[318] = t[404] ^ x[78];
  assign t[319] = t[405] ^ x[77];
  assign t[31] = ~(t[151] ^ t[152]);
  assign t[320] = t[406] ^ x[81];
  assign t[321] = t[407] ^ x[80];
  assign t[322] = t[408] ^ x[84];
  assign t[323] = t[409] ^ x[83];
  assign t[324] = t[410] ^ x[87];
  assign t[325] = t[411] ^ x[86];
  assign t[326] = t[412] ^ x[90];
  assign t[327] = t[413] ^ x[89];
  assign t[328] = t[414] ^ x[93];
  assign t[329] = t[415] ^ x[92];
  assign t[32] = ~(t[24]);
  assign t[330] = t[416] ^ x[96];
  assign t[331] = t[417] ^ x[95];
  assign t[332] = t[418] ^ x[99];
  assign t[333] = t[419] ^ x[98];
  assign t[334] = t[420] ^ x[102];
  assign t[335] = t[421] ^ x[101];
  assign t[336] = t[422] ^ x[105];
  assign t[337] = t[423] ^ x[104];
  assign t[338] = t[424] ^ x[108];
  assign t[339] = t[425] ^ x[107];
  assign t[33] = ~(t[153] & t[42]);
  assign t[340] = t[426] ^ x[111];
  assign t[341] = t[427] ^ x[110];
  assign t[342] = t[428] ^ x[114];
  assign t[343] = t[429] ^ x[113];
  assign t[344] = t[430] ^ x[117];
  assign t[345] = t[431] ^ x[116];
  assign t[346] = t[432] ^ x[120];
  assign t[347] = t[433] ^ x[119];
  assign t[348] = t[434] ^ x[123];
  assign t[349] = t[435] ^ x[122];
  assign t[34] = ~(t[43] & t[44]);
  assign t[350] = t[436] ^ x[126];
  assign t[351] = t[437] ^ x[125];
  assign t[352] = t[438] ^ x[129];
  assign t[353] = t[439] ^ x[128];
  assign t[354] = (x[0]);
  assign t[355] = (x[0]);
  assign t[356] = (x[3]);
  assign t[357] = (x[3]);
  assign t[358] = (x[7]);
  assign t[359] = (x[7]);
  assign t[35] = ~(t[154]);
  assign t[360] = (x[10]);
  assign t[361] = (x[10]);
  assign t[362] = (x[13]);
  assign t[363] = (x[13]);
  assign t[364] = (x[16]);
  assign t[365] = (x[16]);
  assign t[366] = (x[19]);
  assign t[367] = (x[19]);
  assign t[368] = (x[22]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[141]);
  assign t[370] = (x[25]);
  assign t[371] = (x[25]);
  assign t[372] = (x[28]);
  assign t[373] = (x[28]);
  assign t[374] = (x[31]);
  assign t[375] = (x[31]);
  assign t[376] = (x[34]);
  assign t[377] = (x[34]);
  assign t[378] = (x[37]);
  assign t[379] = (x[37]);
  assign t[37] = t[45] & t[46];
  assign t[380] = (x[40]);
  assign t[381] = (x[40]);
  assign t[382] = (x[43]);
  assign t[383] = (x[43]);
  assign t[384] = (x[46]);
  assign t[385] = (x[46]);
  assign t[386] = (x[49]);
  assign t[387] = (x[49]);
  assign t[388] = (x[52]);
  assign t[389] = (x[52]);
  assign t[38] = t[47] ^ t[48];
  assign t[390] = (x[55]);
  assign t[391] = (x[55]);
  assign t[392] = (x[58]);
  assign t[393] = (x[58]);
  assign t[394] = (x[61]);
  assign t[395] = (x[61]);
  assign t[396] = (x[64]);
  assign t[397] = (x[64]);
  assign t[398] = (x[67]);
  assign t[399] = (x[67]);
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[70]);
  assign t[401] = (x[70]);
  assign t[402] = (x[73]);
  assign t[403] = (x[73]);
  assign t[404] = (x[76]);
  assign t[405] = (x[76]);
  assign t[406] = (x[79]);
  assign t[407] = (x[79]);
  assign t[408] = (x[82]);
  assign t[409] = (x[82]);
  assign t[40] = t[51] ^ t[52];
  assign t[410] = (x[85]);
  assign t[411] = (x[85]);
  assign t[412] = (x[88]);
  assign t[413] = (x[88]);
  assign t[414] = (x[91]);
  assign t[415] = (x[91]);
  assign t[416] = (x[94]);
  assign t[417] = (x[94]);
  assign t[418] = (x[97]);
  assign t[419] = (x[97]);
  assign t[41] = t[143] ^ t[155];
  assign t[420] = (x[100]);
  assign t[421] = (x[100]);
  assign t[422] = (x[103]);
  assign t[423] = (x[103]);
  assign t[424] = (x[106]);
  assign t[425] = (x[106]);
  assign t[426] = (x[109]);
  assign t[427] = (x[109]);
  assign t[428] = (x[112]);
  assign t[429] = (x[112]);
  assign t[42] = ~(t[156]);
  assign t[430] = (x[115]);
  assign t[431] = (x[115]);
  assign t[432] = (x[118]);
  assign t[433] = (x[118]);
  assign t[434] = (x[121]);
  assign t[435] = (x[121]);
  assign t[436] = (x[124]);
  assign t[437] = (x[124]);
  assign t[438] = (x[127]);
  assign t[439] = (x[127]);
  assign t[43] = ~(t[157] | t[158]);
  assign t[44] = ~(t[159] | t[160]);
  assign t[45] = t[53] ^ t[54];
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[45] & t[57];
  assign t[48] = t[58] & t[59];
  assign t[49] = t[60] & t[61];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] ^ t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[64] & t[66];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[69] ^ t[70];
  assign t[55] = t[25] ? t[161] : t[71];
  assign t[56] = t[25] ? t[162] : t[72];
  assign t[57] = t[73] ^ t[74];
  assign t[58] = t[60] ^ t[53];
  assign t[59] = t[55] ^ t[75];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[76] ^ t[77];
  assign t[61] = t[66] ^ t[78];
  assign t[62] = t[79] & t[73];
  assign t[63] = t[80] & t[81];
  assign t[64] = t[60] ^ t[80];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[55] ^ t[84];
  assign t[67] = t[85] & t[86];
  assign t[68] = t[85] ^ t[87];
  assign t[69] = t[88] & t[89];
  assign t[6] = ~(t[10]);
  assign t[70] = t[88] ^ t[87];
  assign t[71] = t[163] ^ t[164];
  assign t[72] = t[165] ^ t[166];
  assign t[73] = t[66] ^ t[82];
  assign t[74] = t[90] ^ t[91];
  assign t[75] = t[25] ? t[167] : t[92];
  assign t[76] = t[93] ^ t[94];
  assign t[77] = t[95] & t[85];
  assign t[78] = t[74] ^ t[96];
  assign t[79] = t[80] ^ t[54];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ t[98];
  assign t[81] = t[25] ? t[168] : t[99];
  assign t[82] = t[100] ^ t[75];
  assign t[83] = t[90] ^ t[56];
  assign t[84] = t[25] ? t[169] : t[101];
  assign t[85] = t[102] ^ t[76];
  assign t[86] = t[102] & t[97];
  assign t[87] = t[103] & t[102];
  assign t[88] = t[103] ^ t[97];
  assign t[89] = t[76] & t[103];
  assign t[8] = ~(t[12]);
  assign t[90] = t[25] ? t[170] : t[104];
  assign t[91] = t[25] ? t[171] : t[21];
  assign t[92] = t[172] ^ t[173];
  assign t[93] = t[105] ^ t[106];
  assign t[94] = t[107] ^ t[108];
  assign t[95] = t[97] ^ t[87];
  assign t[96] = t[84] ^ t[81];
  assign t[97] = t[109] ^ t[110];
  assign t[98] = t[111] & t[88];
  assign t[99] = t[174] ^ t[175];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind547(x, y);
 input [129:0] x;
 output y;

 wire [439:0] t;
  assign t[0] = t[1] ? t[2] : t[139];
  assign t[100] = t[25] ? t[176] : t[112];
  assign t[101] = t[155] ^ t[177];
  assign t[102] = t[113] ^ t[114];
  assign t[103] = t[115] ^ t[114];
  assign t[104] = t[178] ^ t[179];
  assign t[105] = t[116] ^ t[117];
  assign t[106] = t[46] ^ t[57];
  assign t[107] = t[46] & t[57];
  assign t[108] = t[66] & t[65];
  assign t[109] = t[118] ^ t[94];
  assign t[10] = t[141] & t[16];
  assign t[110] = t[61] ^ t[119];
  assign t[111] = t[76] ^ t[87];
  assign t[112] = t[180] ^ t[181];
  assign t[113] = t[120] ^ t[121];
  assign t[114] = t[122] ^ t[108];
  assign t[115] = t[123] ^ t[124];
  assign t[116] = t[78] & t[81];
  assign t[117] = t[125] & t[73];
  assign t[118] = t[126] ^ t[127];
  assign t[119] = t[128] ^ t[129];
  assign t[11] = ~(t[17]);
  assign t[120] = t[130] ^ t[117];
  assign t[121] = t[131] & t[132];
  assign t[122] = t[133] & t[134];
  assign t[123] = t[135] ^ t[127];
  assign t[124] = t[136] & t[128];
  assign t[125] = t[59] ^ t[133];
  assign t[126] = t[61] & t[119];
  assign t[127] = t[59] & t[129];
  assign t[128] = t[81] ^ t[74];
  assign t[129] = t[82] ^ t[137];
  assign t[12] = ~(t[141]);
  assign t[130] = t[73] ^ t[83];
  assign t[131] = t[46] ^ t[136];
  assign t[132] = t[81] ^ t[73];
  assign t[133] = t[84] ^ t[56];
  assign t[134] = t[66] ^ t[137];
  assign t[135] = t[59] ^ t[129];
  assign t[136] = t[74] ^ t[138];
  assign t[137] = t[91] ^ t[56];
  assign t[138] = t[75] ^ t[81];
  assign t[139] = (t[182]);
  assign t[13] = ~(t[18]);
  assign t[140] = (t[183]);
  assign t[141] = (t[184]);
  assign t[142] = (t[185]);
  assign t[143] = (t[186]);
  assign t[144] = (t[187]);
  assign t[145] = (t[188]);
  assign t[146] = (t[189]);
  assign t[147] = (t[190]);
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[19] ? t[142] : t[22];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[141] & t[24]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = t[225] ^ x[2];
  assign t[183] = t[226] ^ x[5];
  assign t[184] = t[227] ^ x[9];
  assign t[185] = t[228] ^ x[12];
  assign t[186] = t[229] ^ x[15];
  assign t[187] = t[230] ^ x[18];
  assign t[188] = t[231] ^ x[21];
  assign t[189] = t[232] ^ x[24];
  assign t[18] = ~(t[25]);
  assign t[190] = t[233] ^ x[27];
  assign t[191] = t[234] ^ x[30];
  assign t[192] = t[235] ^ x[33];
  assign t[193] = t[236] ^ x[36];
  assign t[194] = t[237] ^ x[39];
  assign t[195] = t[238] ^ x[42];
  assign t[196] = t[239] ^ x[45];
  assign t[197] = t[240] ^ x[48];
  assign t[198] = t[241] ^ x[51];
  assign t[199] = t[242] ^ x[54];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[57];
  assign t[201] = t[244] ^ x[60];
  assign t[202] = t[245] ^ x[63];
  assign t[203] = t[246] ^ x[66];
  assign t[204] = t[247] ^ x[69];
  assign t[205] = t[248] ^ x[72];
  assign t[206] = t[249] ^ x[75];
  assign t[207] = t[250] ^ x[78];
  assign t[208] = t[251] ^ x[81];
  assign t[209] = t[252] ^ x[84];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[253] ^ x[87];
  assign t[211] = t[254] ^ x[90];
  assign t[212] = t[255] ^ x[93];
  assign t[213] = t[256] ^ x[96];
  assign t[214] = t[257] ^ x[99];
  assign t[215] = t[258] ^ x[102];
  assign t[216] = t[259] ^ x[105];
  assign t[217] = t[260] ^ x[108];
  assign t[218] = t[261] ^ x[111];
  assign t[219] = t[262] ^ x[114];
  assign t[21] = t[143] ^ t[144];
  assign t[220] = t[263] ^ x[117];
  assign t[221] = t[264] ^ x[120];
  assign t[222] = t[265] ^ x[123];
  assign t[223] = t[266] ^ x[126];
  assign t[224] = t[267] ^ x[129];
  assign t[225] = (t[268] & ~t[269]);
  assign t[226] = (t[270] & ~t[271]);
  assign t[227] = (t[272] & ~t[273]);
  assign t[228] = (t[274] & ~t[275]);
  assign t[229] = (t[276] & ~t[277]);
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[278] & ~t[279]);
  assign t[231] = (t[280] & ~t[281]);
  assign t[232] = (t[282] & ~t[283]);
  assign t[233] = (t[284] & ~t[285]);
  assign t[234] = (t[286] & ~t[287]);
  assign t[235] = (t[288] & ~t[289]);
  assign t[236] = (t[290] & ~t[291]);
  assign t[237] = (t[292] & ~t[293]);
  assign t[238] = (t[294] & ~t[295]);
  assign t[239] = (t[296] & ~t[297]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[298] & ~t[299]);
  assign t[241] = (t[300] & ~t[301]);
  assign t[242] = (t[302] & ~t[303]);
  assign t[243] = (t[304] & ~t[305]);
  assign t[244] = (t[306] & ~t[307]);
  assign t[245] = (t[308] & ~t[309]);
  assign t[246] = (t[310] & ~t[311]);
  assign t[247] = (t[312] & ~t[313]);
  assign t[248] = (t[314] & ~t[315]);
  assign t[249] = (t[316] & ~t[317]);
  assign t[24] = ~(t[145] | t[34]);
  assign t[250] = (t[318] & ~t[319]);
  assign t[251] = (t[320] & ~t[321]);
  assign t[252] = (t[322] & ~t[323]);
  assign t[253] = (t[324] & ~t[325]);
  assign t[254] = (t[326] & ~t[327]);
  assign t[255] = (t[328] & ~t[329]);
  assign t[256] = (t[330] & ~t[331]);
  assign t[257] = (t[332] & ~t[333]);
  assign t[258] = (t[334] & ~t[335]);
  assign t[259] = (t[336] & ~t[337]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[338] & ~t[339]);
  assign t[261] = (t[340] & ~t[341]);
  assign t[262] = (t[342] & ~t[343]);
  assign t[263] = (t[344] & ~t[345]);
  assign t[264] = (t[346] & ~t[347]);
  assign t[265] = (t[348] & ~t[349]);
  assign t[266] = (t[350] & ~t[351]);
  assign t[267] = (t[352] & ~t[353]);
  assign t[268] = t[354] ^ x[2];
  assign t[269] = t[355] ^ x[1];
  assign t[26] = ~(t[146] & t[147]);
  assign t[270] = t[356] ^ x[5];
  assign t[271] = t[357] ^ x[4];
  assign t[272] = t[358] ^ x[9];
  assign t[273] = t[359] ^ x[8];
  assign t[274] = t[360] ^ x[12];
  assign t[275] = t[361] ^ x[11];
  assign t[276] = t[362] ^ x[15];
  assign t[277] = t[363] ^ x[14];
  assign t[278] = t[364] ^ x[18];
  assign t[279] = t[365] ^ x[17];
  assign t[27] = ~(t[148] & t[149]);
  assign t[280] = t[366] ^ x[21];
  assign t[281] = t[367] ^ x[20];
  assign t[282] = t[368] ^ x[24];
  assign t[283] = t[369] ^ x[23];
  assign t[284] = t[370] ^ x[27];
  assign t[285] = t[371] ^ x[26];
  assign t[286] = t[372] ^ x[30];
  assign t[287] = t[373] ^ x[29];
  assign t[288] = t[374] ^ x[33];
  assign t[289] = t[375] ^ x[32];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[376] ^ x[36];
  assign t[291] = t[377] ^ x[35];
  assign t[292] = t[378] ^ x[39];
  assign t[293] = t[379] ^ x[38];
  assign t[294] = t[380] ^ x[42];
  assign t[295] = t[381] ^ x[41];
  assign t[296] = t[382] ^ x[45];
  assign t[297] = t[383] ^ x[44];
  assign t[298] = t[384] ^ x[48];
  assign t[299] = t[385] ^ x[47];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[140] : t[5];
  assign t[300] = t[386] ^ x[51];
  assign t[301] = t[387] ^ x[50];
  assign t[302] = t[388] ^ x[54];
  assign t[303] = t[389] ^ x[53];
  assign t[304] = t[390] ^ x[57];
  assign t[305] = t[391] ^ x[56];
  assign t[306] = t[392] ^ x[60];
  assign t[307] = t[393] ^ x[59];
  assign t[308] = t[394] ^ x[63];
  assign t[309] = t[395] ^ x[62];
  assign t[30] = t[150] ^ t[41];
  assign t[310] = t[396] ^ x[66];
  assign t[311] = t[397] ^ x[65];
  assign t[312] = t[398] ^ x[69];
  assign t[313] = t[399] ^ x[68];
  assign t[314] = t[400] ^ x[72];
  assign t[315] = t[401] ^ x[71];
  assign t[316] = t[402] ^ x[75];
  assign t[317] = t[403] ^ x[74];
  assign t[318] = t[404] ^ x[78];
  assign t[319] = t[405] ^ x[77];
  assign t[31] = ~(t[151] ^ t[152]);
  assign t[320] = t[406] ^ x[81];
  assign t[321] = t[407] ^ x[80];
  assign t[322] = t[408] ^ x[84];
  assign t[323] = t[409] ^ x[83];
  assign t[324] = t[410] ^ x[87];
  assign t[325] = t[411] ^ x[86];
  assign t[326] = t[412] ^ x[90];
  assign t[327] = t[413] ^ x[89];
  assign t[328] = t[414] ^ x[93];
  assign t[329] = t[415] ^ x[92];
  assign t[32] = ~(t[24]);
  assign t[330] = t[416] ^ x[96];
  assign t[331] = t[417] ^ x[95];
  assign t[332] = t[418] ^ x[99];
  assign t[333] = t[419] ^ x[98];
  assign t[334] = t[420] ^ x[102];
  assign t[335] = t[421] ^ x[101];
  assign t[336] = t[422] ^ x[105];
  assign t[337] = t[423] ^ x[104];
  assign t[338] = t[424] ^ x[108];
  assign t[339] = t[425] ^ x[107];
  assign t[33] = ~(t[153] & t[42]);
  assign t[340] = t[426] ^ x[111];
  assign t[341] = t[427] ^ x[110];
  assign t[342] = t[428] ^ x[114];
  assign t[343] = t[429] ^ x[113];
  assign t[344] = t[430] ^ x[117];
  assign t[345] = t[431] ^ x[116];
  assign t[346] = t[432] ^ x[120];
  assign t[347] = t[433] ^ x[119];
  assign t[348] = t[434] ^ x[123];
  assign t[349] = t[435] ^ x[122];
  assign t[34] = ~(t[43] & t[44]);
  assign t[350] = t[436] ^ x[126];
  assign t[351] = t[437] ^ x[125];
  assign t[352] = t[438] ^ x[129];
  assign t[353] = t[439] ^ x[128];
  assign t[354] = (x[0]);
  assign t[355] = (x[0]);
  assign t[356] = (x[3]);
  assign t[357] = (x[3]);
  assign t[358] = (x[7]);
  assign t[359] = (x[7]);
  assign t[35] = ~(t[154]);
  assign t[360] = (x[10]);
  assign t[361] = (x[10]);
  assign t[362] = (x[13]);
  assign t[363] = (x[13]);
  assign t[364] = (x[16]);
  assign t[365] = (x[16]);
  assign t[366] = (x[19]);
  assign t[367] = (x[19]);
  assign t[368] = (x[22]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[141]);
  assign t[370] = (x[25]);
  assign t[371] = (x[25]);
  assign t[372] = (x[28]);
  assign t[373] = (x[28]);
  assign t[374] = (x[31]);
  assign t[375] = (x[31]);
  assign t[376] = (x[34]);
  assign t[377] = (x[34]);
  assign t[378] = (x[37]);
  assign t[379] = (x[37]);
  assign t[37] = t[45] & t[46];
  assign t[380] = (x[40]);
  assign t[381] = (x[40]);
  assign t[382] = (x[43]);
  assign t[383] = (x[43]);
  assign t[384] = (x[46]);
  assign t[385] = (x[46]);
  assign t[386] = (x[49]);
  assign t[387] = (x[49]);
  assign t[388] = (x[52]);
  assign t[389] = (x[52]);
  assign t[38] = t[47] ^ t[48];
  assign t[390] = (x[55]);
  assign t[391] = (x[55]);
  assign t[392] = (x[58]);
  assign t[393] = (x[58]);
  assign t[394] = (x[61]);
  assign t[395] = (x[61]);
  assign t[396] = (x[64]);
  assign t[397] = (x[64]);
  assign t[398] = (x[67]);
  assign t[399] = (x[67]);
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[70]);
  assign t[401] = (x[70]);
  assign t[402] = (x[73]);
  assign t[403] = (x[73]);
  assign t[404] = (x[76]);
  assign t[405] = (x[76]);
  assign t[406] = (x[79]);
  assign t[407] = (x[79]);
  assign t[408] = (x[82]);
  assign t[409] = (x[82]);
  assign t[40] = t[51] ^ t[52];
  assign t[410] = (x[85]);
  assign t[411] = (x[85]);
  assign t[412] = (x[88]);
  assign t[413] = (x[88]);
  assign t[414] = (x[91]);
  assign t[415] = (x[91]);
  assign t[416] = (x[94]);
  assign t[417] = (x[94]);
  assign t[418] = (x[97]);
  assign t[419] = (x[97]);
  assign t[41] = t[143] ^ t[155];
  assign t[420] = (x[100]);
  assign t[421] = (x[100]);
  assign t[422] = (x[103]);
  assign t[423] = (x[103]);
  assign t[424] = (x[106]);
  assign t[425] = (x[106]);
  assign t[426] = (x[109]);
  assign t[427] = (x[109]);
  assign t[428] = (x[112]);
  assign t[429] = (x[112]);
  assign t[42] = ~(t[156]);
  assign t[430] = (x[115]);
  assign t[431] = (x[115]);
  assign t[432] = (x[118]);
  assign t[433] = (x[118]);
  assign t[434] = (x[121]);
  assign t[435] = (x[121]);
  assign t[436] = (x[124]);
  assign t[437] = (x[124]);
  assign t[438] = (x[127]);
  assign t[439] = (x[127]);
  assign t[43] = ~(t[157] | t[158]);
  assign t[44] = ~(t[159] | t[160]);
  assign t[45] = t[53] ^ t[54];
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[45] & t[57];
  assign t[48] = t[58] & t[59];
  assign t[49] = t[60] & t[61];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] ^ t[63];
  assign t[51] = t[64] & t[65];
  assign t[52] = t[64] & t[66];
  assign t[53] = t[67] ^ t[68];
  assign t[54] = t[69] ^ t[70];
  assign t[55] = t[25] ? t[161] : t[71];
  assign t[56] = t[25] ? t[162] : t[72];
  assign t[57] = t[73] ^ t[74];
  assign t[58] = t[60] ^ t[53];
  assign t[59] = t[55] ^ t[75];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[76] ^ t[77];
  assign t[61] = t[66] ^ t[78];
  assign t[62] = t[79] & t[73];
  assign t[63] = t[80] & t[81];
  assign t[64] = t[60] ^ t[80];
  assign t[65] = t[82] ^ t[83];
  assign t[66] = t[55] ^ t[84];
  assign t[67] = t[85] & t[86];
  assign t[68] = t[85] ^ t[87];
  assign t[69] = t[88] & t[89];
  assign t[6] = ~(t[10]);
  assign t[70] = t[88] ^ t[87];
  assign t[71] = t[163] ^ t[164];
  assign t[72] = t[165] ^ t[166];
  assign t[73] = t[66] ^ t[82];
  assign t[74] = t[90] ^ t[91];
  assign t[75] = t[25] ? t[167] : t[92];
  assign t[76] = t[93] ^ t[94];
  assign t[77] = t[95] & t[85];
  assign t[78] = t[74] ^ t[96];
  assign t[79] = t[80] ^ t[54];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] ^ t[98];
  assign t[81] = t[25] ? t[168] : t[99];
  assign t[82] = t[100] ^ t[75];
  assign t[83] = t[90] ^ t[56];
  assign t[84] = t[25] ? t[169] : t[101];
  assign t[85] = t[102] ^ t[76];
  assign t[86] = t[102] & t[97];
  assign t[87] = t[103] & t[102];
  assign t[88] = t[103] ^ t[97];
  assign t[89] = t[76] & t[103];
  assign t[8] = ~(t[12]);
  assign t[90] = t[25] ? t[170] : t[104];
  assign t[91] = t[25] ? t[171] : t[21];
  assign t[92] = t[172] ^ t[173];
  assign t[93] = t[105] ^ t[106];
  assign t[94] = t[107] ^ t[108];
  assign t[95] = t[97] ^ t[87];
  assign t[96] = t[84] ^ t[81];
  assign t[97] = t[109] ^ t[110];
  assign t[98] = t[111] & t[88];
  assign t[99] = t[174] ^ t[175];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind548(x, y);
 input [129:0] x;
 output y;

 wire [439:0] t;
  assign t[0] = t[1] ? t[2] : t[139];
  assign t[100] = t[117] ^ t[118];
  assign t[101] = t[119] ^ t[104];
  assign t[102] = t[120] ^ t[121];
  assign t[103] = t[122] ^ t[123];
  assign t[104] = t[124] ^ t[118];
  assign t[105] = t[125] ^ t[126];
  assign t[106] = t[155] ^ t[175];
  assign t[107] = t[176] ^ t[177];
  assign t[108] = t[178] ^ t[179];
  assign t[109] = t[84] ^ t[69];
  assign t[10] = t[141] & t[16];
  assign t[110] = t[86] ^ t[85];
  assign t[111] = t[85] ^ t[69];
  assign t[112] = t[110] & t[127];
  assign t[113] = t[110] ^ t[69];
  assign t[114] = t[180] ^ t[181];
  assign t[115] = t[128] ^ t[129];
  assign t[116] = t[56] & t[130];
  assign t[117] = t[60] & t[66];
  assign t[118] = t[58] & t[65];
  assign t[119] = t[131] ^ t[129];
  assign t[11] = ~(t[17]);
  assign t[120] = t[58] ^ t[132];
  assign t[121] = t[130] ^ t[133];
  assign t[122] = t[134] ^ t[135];
  assign t[123] = t[55] ^ t[136];
  assign t[124] = t[55] & t[136];
  assign t[125] = t[137] ^ t[135];
  assign t[126] = t[46] & t[79];
  assign t[127] = t[86] & t[84];
  assign t[128] = t[98] ^ t[133];
  assign t[129] = t[98] & t[133];
  assign t[12] = ~(t[141]);
  assign t[130] = t[92] ^ t[72];
  assign t[131] = t[120] & t[121];
  assign t[132] = t[72] ^ t[138];
  assign t[133] = t[78] ^ t[82];
  assign t[134] = t[132] & t[92];
  assign t[135] = t[80] & t[62];
  assign t[136] = t[62] ^ t[72];
  assign t[137] = t[62] ^ t[81];
  assign t[138] = t[76] ^ t[92];
  assign t[139] = (t[182]);
  assign t[13] = ~(t[18]);
  assign t[140] = (t[183]);
  assign t[141] = (t[184]);
  assign t[142] = (t[185]);
  assign t[143] = (t[186]);
  assign t[144] = (t[187]);
  assign t[145] = (t[188]);
  assign t[146] = (t[189]);
  assign t[147] = (t[190]);
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[19] ? t[142] : t[22];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[141] & t[24]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = t[225] ^ x[2];
  assign t[183] = t[226] ^ x[5];
  assign t[184] = t[227] ^ x[9];
  assign t[185] = t[228] ^ x[12];
  assign t[186] = t[229] ^ x[15];
  assign t[187] = t[230] ^ x[18];
  assign t[188] = t[231] ^ x[21];
  assign t[189] = t[232] ^ x[24];
  assign t[18] = ~(t[25]);
  assign t[190] = t[233] ^ x[27];
  assign t[191] = t[234] ^ x[30];
  assign t[192] = t[235] ^ x[33];
  assign t[193] = t[236] ^ x[36];
  assign t[194] = t[237] ^ x[39];
  assign t[195] = t[238] ^ x[42];
  assign t[196] = t[239] ^ x[45];
  assign t[197] = t[240] ^ x[48];
  assign t[198] = t[241] ^ x[51];
  assign t[199] = t[242] ^ x[54];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[57];
  assign t[201] = t[244] ^ x[60];
  assign t[202] = t[245] ^ x[63];
  assign t[203] = t[246] ^ x[66];
  assign t[204] = t[247] ^ x[69];
  assign t[205] = t[248] ^ x[72];
  assign t[206] = t[249] ^ x[75];
  assign t[207] = t[250] ^ x[78];
  assign t[208] = t[251] ^ x[81];
  assign t[209] = t[252] ^ x[84];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[253] ^ x[87];
  assign t[211] = t[254] ^ x[90];
  assign t[212] = t[255] ^ x[93];
  assign t[213] = t[256] ^ x[96];
  assign t[214] = t[257] ^ x[99];
  assign t[215] = t[258] ^ x[102];
  assign t[216] = t[259] ^ x[105];
  assign t[217] = t[260] ^ x[108];
  assign t[218] = t[261] ^ x[111];
  assign t[219] = t[262] ^ x[114];
  assign t[21] = t[143] ^ t[144];
  assign t[220] = t[263] ^ x[117];
  assign t[221] = t[264] ^ x[120];
  assign t[222] = t[265] ^ x[123];
  assign t[223] = t[266] ^ x[126];
  assign t[224] = t[267] ^ x[129];
  assign t[225] = (t[268] & ~t[269]);
  assign t[226] = (t[270] & ~t[271]);
  assign t[227] = (t[272] & ~t[273]);
  assign t[228] = (t[274] & ~t[275]);
  assign t[229] = (t[276] & ~t[277]);
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[278] & ~t[279]);
  assign t[231] = (t[280] & ~t[281]);
  assign t[232] = (t[282] & ~t[283]);
  assign t[233] = (t[284] & ~t[285]);
  assign t[234] = (t[286] & ~t[287]);
  assign t[235] = (t[288] & ~t[289]);
  assign t[236] = (t[290] & ~t[291]);
  assign t[237] = (t[292] & ~t[293]);
  assign t[238] = (t[294] & ~t[295]);
  assign t[239] = (t[296] & ~t[297]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[298] & ~t[299]);
  assign t[241] = (t[300] & ~t[301]);
  assign t[242] = (t[302] & ~t[303]);
  assign t[243] = (t[304] & ~t[305]);
  assign t[244] = (t[306] & ~t[307]);
  assign t[245] = (t[308] & ~t[309]);
  assign t[246] = (t[310] & ~t[311]);
  assign t[247] = (t[312] & ~t[313]);
  assign t[248] = (t[314] & ~t[315]);
  assign t[249] = (t[316] & ~t[317]);
  assign t[24] = ~(t[145] | t[34]);
  assign t[250] = (t[318] & ~t[319]);
  assign t[251] = (t[320] & ~t[321]);
  assign t[252] = (t[322] & ~t[323]);
  assign t[253] = (t[324] & ~t[325]);
  assign t[254] = (t[326] & ~t[327]);
  assign t[255] = (t[328] & ~t[329]);
  assign t[256] = (t[330] & ~t[331]);
  assign t[257] = (t[332] & ~t[333]);
  assign t[258] = (t[334] & ~t[335]);
  assign t[259] = (t[336] & ~t[337]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[338] & ~t[339]);
  assign t[261] = (t[340] & ~t[341]);
  assign t[262] = (t[342] & ~t[343]);
  assign t[263] = (t[344] & ~t[345]);
  assign t[264] = (t[346] & ~t[347]);
  assign t[265] = (t[348] & ~t[349]);
  assign t[266] = (t[350] & ~t[351]);
  assign t[267] = (t[352] & ~t[353]);
  assign t[268] = t[354] ^ x[2];
  assign t[269] = t[355] ^ x[1];
  assign t[26] = ~(t[146] & t[147]);
  assign t[270] = t[356] ^ x[5];
  assign t[271] = t[357] ^ x[4];
  assign t[272] = t[358] ^ x[9];
  assign t[273] = t[359] ^ x[8];
  assign t[274] = t[360] ^ x[12];
  assign t[275] = t[361] ^ x[11];
  assign t[276] = t[362] ^ x[15];
  assign t[277] = t[363] ^ x[14];
  assign t[278] = t[364] ^ x[18];
  assign t[279] = t[365] ^ x[17];
  assign t[27] = ~(t[148] & t[149]);
  assign t[280] = t[366] ^ x[21];
  assign t[281] = t[367] ^ x[20];
  assign t[282] = t[368] ^ x[24];
  assign t[283] = t[369] ^ x[23];
  assign t[284] = t[370] ^ x[27];
  assign t[285] = t[371] ^ x[26];
  assign t[286] = t[372] ^ x[30];
  assign t[287] = t[373] ^ x[29];
  assign t[288] = t[374] ^ x[33];
  assign t[289] = t[375] ^ x[32];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[376] ^ x[36];
  assign t[291] = t[377] ^ x[35];
  assign t[292] = t[378] ^ x[39];
  assign t[293] = t[379] ^ x[38];
  assign t[294] = t[380] ^ x[42];
  assign t[295] = t[381] ^ x[41];
  assign t[296] = t[382] ^ x[45];
  assign t[297] = t[383] ^ x[44];
  assign t[298] = t[384] ^ x[48];
  assign t[299] = t[385] ^ x[47];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[140] : t[5];
  assign t[300] = t[386] ^ x[51];
  assign t[301] = t[387] ^ x[50];
  assign t[302] = t[388] ^ x[54];
  assign t[303] = t[389] ^ x[53];
  assign t[304] = t[390] ^ x[57];
  assign t[305] = t[391] ^ x[56];
  assign t[306] = t[392] ^ x[60];
  assign t[307] = t[393] ^ x[59];
  assign t[308] = t[394] ^ x[63];
  assign t[309] = t[395] ^ x[62];
  assign t[30] = t[150] ^ t[41];
  assign t[310] = t[396] ^ x[66];
  assign t[311] = t[397] ^ x[65];
  assign t[312] = t[398] ^ x[69];
  assign t[313] = t[399] ^ x[68];
  assign t[314] = t[400] ^ x[72];
  assign t[315] = t[401] ^ x[71];
  assign t[316] = t[402] ^ x[75];
  assign t[317] = t[403] ^ x[74];
  assign t[318] = t[404] ^ x[78];
  assign t[319] = t[405] ^ x[77];
  assign t[31] = ~(t[151] ^ t[152]);
  assign t[320] = t[406] ^ x[81];
  assign t[321] = t[407] ^ x[80];
  assign t[322] = t[408] ^ x[84];
  assign t[323] = t[409] ^ x[83];
  assign t[324] = t[410] ^ x[87];
  assign t[325] = t[411] ^ x[86];
  assign t[326] = t[412] ^ x[90];
  assign t[327] = t[413] ^ x[89];
  assign t[328] = t[414] ^ x[93];
  assign t[329] = t[415] ^ x[92];
  assign t[32] = ~(t[24]);
  assign t[330] = t[416] ^ x[96];
  assign t[331] = t[417] ^ x[95];
  assign t[332] = t[418] ^ x[99];
  assign t[333] = t[419] ^ x[98];
  assign t[334] = t[420] ^ x[102];
  assign t[335] = t[421] ^ x[101];
  assign t[336] = t[422] ^ x[105];
  assign t[337] = t[423] ^ x[104];
  assign t[338] = t[424] ^ x[108];
  assign t[339] = t[425] ^ x[107];
  assign t[33] = ~(t[153] & t[42]);
  assign t[340] = t[426] ^ x[111];
  assign t[341] = t[427] ^ x[110];
  assign t[342] = t[428] ^ x[114];
  assign t[343] = t[429] ^ x[113];
  assign t[344] = t[430] ^ x[117];
  assign t[345] = t[431] ^ x[116];
  assign t[346] = t[432] ^ x[120];
  assign t[347] = t[433] ^ x[119];
  assign t[348] = t[434] ^ x[123];
  assign t[349] = t[435] ^ x[122];
  assign t[34] = ~(t[43] & t[44]);
  assign t[350] = t[436] ^ x[126];
  assign t[351] = t[437] ^ x[125];
  assign t[352] = t[438] ^ x[129];
  assign t[353] = t[439] ^ x[128];
  assign t[354] = (x[0]);
  assign t[355] = (x[0]);
  assign t[356] = (x[3]);
  assign t[357] = (x[3]);
  assign t[358] = (x[7]);
  assign t[359] = (x[7]);
  assign t[35] = ~(t[154]);
  assign t[360] = (x[10]);
  assign t[361] = (x[10]);
  assign t[362] = (x[13]);
  assign t[363] = (x[13]);
  assign t[364] = (x[16]);
  assign t[365] = (x[16]);
  assign t[366] = (x[19]);
  assign t[367] = (x[19]);
  assign t[368] = (x[22]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[141]);
  assign t[370] = (x[25]);
  assign t[371] = (x[25]);
  assign t[372] = (x[28]);
  assign t[373] = (x[28]);
  assign t[374] = (x[31]);
  assign t[375] = (x[31]);
  assign t[376] = (x[34]);
  assign t[377] = (x[34]);
  assign t[378] = (x[37]);
  assign t[379] = (x[37]);
  assign t[37] = t[45] & t[46];
  assign t[380] = (x[40]);
  assign t[381] = (x[40]);
  assign t[382] = (x[43]);
  assign t[383] = (x[43]);
  assign t[384] = (x[46]);
  assign t[385] = (x[46]);
  assign t[386] = (x[49]);
  assign t[387] = (x[49]);
  assign t[388] = (x[52]);
  assign t[389] = (x[52]);
  assign t[38] = t[47] ^ t[48];
  assign t[390] = (x[55]);
  assign t[391] = (x[55]);
  assign t[392] = (x[58]);
  assign t[393] = (x[58]);
  assign t[394] = (x[61]);
  assign t[395] = (x[61]);
  assign t[396] = (x[64]);
  assign t[397] = (x[64]);
  assign t[398] = (x[67]);
  assign t[399] = (x[67]);
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[70]);
  assign t[401] = (x[70]);
  assign t[402] = (x[73]);
  assign t[403] = (x[73]);
  assign t[404] = (x[76]);
  assign t[405] = (x[76]);
  assign t[406] = (x[79]);
  assign t[407] = (x[79]);
  assign t[408] = (x[82]);
  assign t[409] = (x[82]);
  assign t[40] = t[51] ^ t[52];
  assign t[410] = (x[85]);
  assign t[411] = (x[85]);
  assign t[412] = (x[88]);
  assign t[413] = (x[88]);
  assign t[414] = (x[91]);
  assign t[415] = (x[91]);
  assign t[416] = (x[94]);
  assign t[417] = (x[94]);
  assign t[418] = (x[97]);
  assign t[419] = (x[97]);
  assign t[41] = t[143] ^ t[155];
  assign t[420] = (x[100]);
  assign t[421] = (x[100]);
  assign t[422] = (x[103]);
  assign t[423] = (x[103]);
  assign t[424] = (x[106]);
  assign t[425] = (x[106]);
  assign t[426] = (x[109]);
  assign t[427] = (x[109]);
  assign t[428] = (x[112]);
  assign t[429] = (x[112]);
  assign t[42] = ~(t[156]);
  assign t[430] = (x[115]);
  assign t[431] = (x[115]);
  assign t[432] = (x[118]);
  assign t[433] = (x[118]);
  assign t[434] = (x[121]);
  assign t[435] = (x[121]);
  assign t[436] = (x[124]);
  assign t[437] = (x[124]);
  assign t[438] = (x[127]);
  assign t[439] = (x[127]);
  assign t[43] = ~(t[157] | t[158]);
  assign t[44] = ~(t[159] | t[160]);
  assign t[45] = t[53] ^ t[54];
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[57] & t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[61] & t[62];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ t[64];
  assign t[51] = t[57] & t[65];
  assign t[52] = t[59] & t[66];
  assign t[53] = t[67] & t[68];
  assign t[54] = t[67] ^ t[69];
  assign t[55] = t[70] ^ t[71];
  assign t[56] = t[72] ^ t[73];
  assign t[57] = t[74] ^ t[75];
  assign t[58] = t[70] ^ t[76];
  assign t[59] = t[57] ^ t[77];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[76] ^ t[71];
  assign t[61] = t[75] ^ t[45];
  assign t[62] = t[58] ^ t[78];
  assign t[63] = t[45] & t[79];
  assign t[64] = t[61] & t[80];
  assign t[65] = t[78] ^ t[81];
  assign t[66] = t[58] ^ t[82];
  assign t[67] = t[83] ^ t[84];
  assign t[68] = t[85] & t[83];
  assign t[69] = t[83] & t[86];
  assign t[6] = ~(t[10]);
  assign t[70] = t[25] ? t[161] : t[87];
  assign t[71] = t[25] ? t[162] : t[88];
  assign t[72] = t[89] ^ t[90];
  assign t[73] = t[91] ^ t[92];
  assign t[74] = t[85] ^ t[93];
  assign t[75] = t[84] ^ t[94];
  assign t[76] = t[25] ? t[163] : t[95];
  assign t[77] = t[96] ^ t[45];
  assign t[78] = t[97] ^ t[91];
  assign t[79] = t[92] ^ t[62];
  assign t[7] = ~(t[11]);
  assign t[80] = t[98] ^ t[60];
  assign t[81] = t[89] ^ t[71];
  assign t[82] = t[90] ^ t[71];
  assign t[83] = t[99] ^ t[100];
  assign t[84] = t[101] ^ t[102];
  assign t[85] = t[103] ^ t[104];
  assign t[86] = t[105] ^ t[100];
  assign t[87] = t[164] ^ t[165];
  assign t[88] = t[166] ^ t[167];
  assign t[89] = t[25] ? t[168] : t[21];
  assign t[8] = ~(t[12]);
  assign t[90] = t[25] ? t[169] : t[106];
  assign t[91] = t[25] ? t[170] : t[107];
  assign t[92] = t[25] ? t[171] : t[108];
  assign t[93] = t[109] & t[110];
  assign t[94] = t[111] & t[67];
  assign t[95] = t[172] ^ t[173];
  assign t[96] = t[112] ^ t[113];
  assign t[97] = t[25] ? t[174] : t[114];
  assign t[98] = t[70] ^ t[91];
  assign t[99] = t[115] ^ t[116];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind549(x, y);
 input [129:0] x;
 output y;

 wire [439:0] t;
  assign t[0] = t[1] ? t[2] : t[139];
  assign t[100] = t[117] ^ t[118];
  assign t[101] = t[119] ^ t[104];
  assign t[102] = t[120] ^ t[121];
  assign t[103] = t[122] ^ t[123];
  assign t[104] = t[124] ^ t[118];
  assign t[105] = t[125] ^ t[126];
  assign t[106] = t[155] ^ t[175];
  assign t[107] = t[176] ^ t[177];
  assign t[108] = t[178] ^ t[179];
  assign t[109] = t[84] ^ t[69];
  assign t[10] = t[141] & t[16];
  assign t[110] = t[86] ^ t[85];
  assign t[111] = t[85] ^ t[69];
  assign t[112] = t[110] & t[127];
  assign t[113] = t[110] ^ t[69];
  assign t[114] = t[180] ^ t[181];
  assign t[115] = t[128] ^ t[129];
  assign t[116] = t[56] & t[130];
  assign t[117] = t[60] & t[66];
  assign t[118] = t[58] & t[65];
  assign t[119] = t[131] ^ t[129];
  assign t[11] = ~(t[17]);
  assign t[120] = t[58] ^ t[132];
  assign t[121] = t[130] ^ t[133];
  assign t[122] = t[134] ^ t[135];
  assign t[123] = t[55] ^ t[136];
  assign t[124] = t[55] & t[136];
  assign t[125] = t[137] ^ t[135];
  assign t[126] = t[46] & t[79];
  assign t[127] = t[86] & t[84];
  assign t[128] = t[98] ^ t[133];
  assign t[129] = t[98] & t[133];
  assign t[12] = ~(t[141]);
  assign t[130] = t[92] ^ t[72];
  assign t[131] = t[120] & t[121];
  assign t[132] = t[72] ^ t[138];
  assign t[133] = t[78] ^ t[82];
  assign t[134] = t[132] & t[92];
  assign t[135] = t[80] & t[62];
  assign t[136] = t[62] ^ t[72];
  assign t[137] = t[62] ^ t[81];
  assign t[138] = t[76] ^ t[92];
  assign t[139] = (t[182]);
  assign t[13] = ~(t[18]);
  assign t[140] = (t[183]);
  assign t[141] = (t[184]);
  assign t[142] = (t[185]);
  assign t[143] = (t[186]);
  assign t[144] = (t[187]);
  assign t[145] = (t[188]);
  assign t[146] = (t[189]);
  assign t[147] = (t[190]);
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[19] ? t[142] : t[22];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[141] & t[24]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = t[225] ^ x[2];
  assign t[183] = t[226] ^ x[5];
  assign t[184] = t[227] ^ x[9];
  assign t[185] = t[228] ^ x[12];
  assign t[186] = t[229] ^ x[15];
  assign t[187] = t[230] ^ x[18];
  assign t[188] = t[231] ^ x[21];
  assign t[189] = t[232] ^ x[24];
  assign t[18] = ~(t[25]);
  assign t[190] = t[233] ^ x[27];
  assign t[191] = t[234] ^ x[30];
  assign t[192] = t[235] ^ x[33];
  assign t[193] = t[236] ^ x[36];
  assign t[194] = t[237] ^ x[39];
  assign t[195] = t[238] ^ x[42];
  assign t[196] = t[239] ^ x[45];
  assign t[197] = t[240] ^ x[48];
  assign t[198] = t[241] ^ x[51];
  assign t[199] = t[242] ^ x[54];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[57];
  assign t[201] = t[244] ^ x[60];
  assign t[202] = t[245] ^ x[63];
  assign t[203] = t[246] ^ x[66];
  assign t[204] = t[247] ^ x[69];
  assign t[205] = t[248] ^ x[72];
  assign t[206] = t[249] ^ x[75];
  assign t[207] = t[250] ^ x[78];
  assign t[208] = t[251] ^ x[81];
  assign t[209] = t[252] ^ x[84];
  assign t[20] = ~(t[28] ^ t[29]);
  assign t[210] = t[253] ^ x[87];
  assign t[211] = t[254] ^ x[90];
  assign t[212] = t[255] ^ x[93];
  assign t[213] = t[256] ^ x[96];
  assign t[214] = t[257] ^ x[99];
  assign t[215] = t[258] ^ x[102];
  assign t[216] = t[259] ^ x[105];
  assign t[217] = t[260] ^ x[108];
  assign t[218] = t[261] ^ x[111];
  assign t[219] = t[262] ^ x[114];
  assign t[21] = t[143] ^ t[144];
  assign t[220] = t[263] ^ x[117];
  assign t[221] = t[264] ^ x[120];
  assign t[222] = t[265] ^ x[123];
  assign t[223] = t[266] ^ x[126];
  assign t[224] = t[267] ^ x[129];
  assign t[225] = (t[268] & ~t[269]);
  assign t[226] = (t[270] & ~t[271]);
  assign t[227] = (t[272] & ~t[273]);
  assign t[228] = (t[274] & ~t[275]);
  assign t[229] = (t[276] & ~t[277]);
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[278] & ~t[279]);
  assign t[231] = (t[280] & ~t[281]);
  assign t[232] = (t[282] & ~t[283]);
  assign t[233] = (t[284] & ~t[285]);
  assign t[234] = (t[286] & ~t[287]);
  assign t[235] = (t[288] & ~t[289]);
  assign t[236] = (t[290] & ~t[291]);
  assign t[237] = (t[292] & ~t[293]);
  assign t[238] = (t[294] & ~t[295]);
  assign t[239] = (t[296] & ~t[297]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[298] & ~t[299]);
  assign t[241] = (t[300] & ~t[301]);
  assign t[242] = (t[302] & ~t[303]);
  assign t[243] = (t[304] & ~t[305]);
  assign t[244] = (t[306] & ~t[307]);
  assign t[245] = (t[308] & ~t[309]);
  assign t[246] = (t[310] & ~t[311]);
  assign t[247] = (t[312] & ~t[313]);
  assign t[248] = (t[314] & ~t[315]);
  assign t[249] = (t[316] & ~t[317]);
  assign t[24] = ~(t[145] | t[34]);
  assign t[250] = (t[318] & ~t[319]);
  assign t[251] = (t[320] & ~t[321]);
  assign t[252] = (t[322] & ~t[323]);
  assign t[253] = (t[324] & ~t[325]);
  assign t[254] = (t[326] & ~t[327]);
  assign t[255] = (t[328] & ~t[329]);
  assign t[256] = (t[330] & ~t[331]);
  assign t[257] = (t[332] & ~t[333]);
  assign t[258] = (t[334] & ~t[335]);
  assign t[259] = (t[336] & ~t[337]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[338] & ~t[339]);
  assign t[261] = (t[340] & ~t[341]);
  assign t[262] = (t[342] & ~t[343]);
  assign t[263] = (t[344] & ~t[345]);
  assign t[264] = (t[346] & ~t[347]);
  assign t[265] = (t[348] & ~t[349]);
  assign t[266] = (t[350] & ~t[351]);
  assign t[267] = (t[352] & ~t[353]);
  assign t[268] = t[354] ^ x[2];
  assign t[269] = t[355] ^ x[1];
  assign t[26] = ~(t[146] & t[147]);
  assign t[270] = t[356] ^ x[5];
  assign t[271] = t[357] ^ x[4];
  assign t[272] = t[358] ^ x[9];
  assign t[273] = t[359] ^ x[8];
  assign t[274] = t[360] ^ x[12];
  assign t[275] = t[361] ^ x[11];
  assign t[276] = t[362] ^ x[15];
  assign t[277] = t[363] ^ x[14];
  assign t[278] = t[364] ^ x[18];
  assign t[279] = t[365] ^ x[17];
  assign t[27] = ~(t[148] & t[149]);
  assign t[280] = t[366] ^ x[21];
  assign t[281] = t[367] ^ x[20];
  assign t[282] = t[368] ^ x[24];
  assign t[283] = t[369] ^ x[23];
  assign t[284] = t[370] ^ x[27];
  assign t[285] = t[371] ^ x[26];
  assign t[286] = t[372] ^ x[30];
  assign t[287] = t[373] ^ x[29];
  assign t[288] = t[374] ^ x[33];
  assign t[289] = t[375] ^ x[32];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[376] ^ x[36];
  assign t[291] = t[377] ^ x[35];
  assign t[292] = t[378] ^ x[39];
  assign t[293] = t[379] ^ x[38];
  assign t[294] = t[380] ^ x[42];
  assign t[295] = t[381] ^ x[41];
  assign t[296] = t[382] ^ x[45];
  assign t[297] = t[383] ^ x[44];
  assign t[298] = t[384] ^ x[48];
  assign t[299] = t[385] ^ x[47];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[140] : t[5];
  assign t[300] = t[386] ^ x[51];
  assign t[301] = t[387] ^ x[50];
  assign t[302] = t[388] ^ x[54];
  assign t[303] = t[389] ^ x[53];
  assign t[304] = t[390] ^ x[57];
  assign t[305] = t[391] ^ x[56];
  assign t[306] = t[392] ^ x[60];
  assign t[307] = t[393] ^ x[59];
  assign t[308] = t[394] ^ x[63];
  assign t[309] = t[395] ^ x[62];
  assign t[30] = t[150] ^ t[41];
  assign t[310] = t[396] ^ x[66];
  assign t[311] = t[397] ^ x[65];
  assign t[312] = t[398] ^ x[69];
  assign t[313] = t[399] ^ x[68];
  assign t[314] = t[400] ^ x[72];
  assign t[315] = t[401] ^ x[71];
  assign t[316] = t[402] ^ x[75];
  assign t[317] = t[403] ^ x[74];
  assign t[318] = t[404] ^ x[78];
  assign t[319] = t[405] ^ x[77];
  assign t[31] = ~(t[151] ^ t[152]);
  assign t[320] = t[406] ^ x[81];
  assign t[321] = t[407] ^ x[80];
  assign t[322] = t[408] ^ x[84];
  assign t[323] = t[409] ^ x[83];
  assign t[324] = t[410] ^ x[87];
  assign t[325] = t[411] ^ x[86];
  assign t[326] = t[412] ^ x[90];
  assign t[327] = t[413] ^ x[89];
  assign t[328] = t[414] ^ x[93];
  assign t[329] = t[415] ^ x[92];
  assign t[32] = ~(t[24]);
  assign t[330] = t[416] ^ x[96];
  assign t[331] = t[417] ^ x[95];
  assign t[332] = t[418] ^ x[99];
  assign t[333] = t[419] ^ x[98];
  assign t[334] = t[420] ^ x[102];
  assign t[335] = t[421] ^ x[101];
  assign t[336] = t[422] ^ x[105];
  assign t[337] = t[423] ^ x[104];
  assign t[338] = t[424] ^ x[108];
  assign t[339] = t[425] ^ x[107];
  assign t[33] = ~(t[153] & t[42]);
  assign t[340] = t[426] ^ x[111];
  assign t[341] = t[427] ^ x[110];
  assign t[342] = t[428] ^ x[114];
  assign t[343] = t[429] ^ x[113];
  assign t[344] = t[430] ^ x[117];
  assign t[345] = t[431] ^ x[116];
  assign t[346] = t[432] ^ x[120];
  assign t[347] = t[433] ^ x[119];
  assign t[348] = t[434] ^ x[123];
  assign t[349] = t[435] ^ x[122];
  assign t[34] = ~(t[43] & t[44]);
  assign t[350] = t[436] ^ x[126];
  assign t[351] = t[437] ^ x[125];
  assign t[352] = t[438] ^ x[129];
  assign t[353] = t[439] ^ x[128];
  assign t[354] = (x[0]);
  assign t[355] = (x[0]);
  assign t[356] = (x[3]);
  assign t[357] = (x[3]);
  assign t[358] = (x[7]);
  assign t[359] = (x[7]);
  assign t[35] = ~(t[154]);
  assign t[360] = (x[10]);
  assign t[361] = (x[10]);
  assign t[362] = (x[13]);
  assign t[363] = (x[13]);
  assign t[364] = (x[16]);
  assign t[365] = (x[16]);
  assign t[366] = (x[19]);
  assign t[367] = (x[19]);
  assign t[368] = (x[22]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[141]);
  assign t[370] = (x[25]);
  assign t[371] = (x[25]);
  assign t[372] = (x[28]);
  assign t[373] = (x[28]);
  assign t[374] = (x[31]);
  assign t[375] = (x[31]);
  assign t[376] = (x[34]);
  assign t[377] = (x[34]);
  assign t[378] = (x[37]);
  assign t[379] = (x[37]);
  assign t[37] = t[45] & t[46];
  assign t[380] = (x[40]);
  assign t[381] = (x[40]);
  assign t[382] = (x[43]);
  assign t[383] = (x[43]);
  assign t[384] = (x[46]);
  assign t[385] = (x[46]);
  assign t[386] = (x[49]);
  assign t[387] = (x[49]);
  assign t[388] = (x[52]);
  assign t[389] = (x[52]);
  assign t[38] = t[47] ^ t[48];
  assign t[390] = (x[55]);
  assign t[391] = (x[55]);
  assign t[392] = (x[58]);
  assign t[393] = (x[58]);
  assign t[394] = (x[61]);
  assign t[395] = (x[61]);
  assign t[396] = (x[64]);
  assign t[397] = (x[64]);
  assign t[398] = (x[67]);
  assign t[399] = (x[67]);
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[70]);
  assign t[401] = (x[70]);
  assign t[402] = (x[73]);
  assign t[403] = (x[73]);
  assign t[404] = (x[76]);
  assign t[405] = (x[76]);
  assign t[406] = (x[79]);
  assign t[407] = (x[79]);
  assign t[408] = (x[82]);
  assign t[409] = (x[82]);
  assign t[40] = t[51] ^ t[52];
  assign t[410] = (x[85]);
  assign t[411] = (x[85]);
  assign t[412] = (x[88]);
  assign t[413] = (x[88]);
  assign t[414] = (x[91]);
  assign t[415] = (x[91]);
  assign t[416] = (x[94]);
  assign t[417] = (x[94]);
  assign t[418] = (x[97]);
  assign t[419] = (x[97]);
  assign t[41] = t[143] ^ t[155];
  assign t[420] = (x[100]);
  assign t[421] = (x[100]);
  assign t[422] = (x[103]);
  assign t[423] = (x[103]);
  assign t[424] = (x[106]);
  assign t[425] = (x[106]);
  assign t[426] = (x[109]);
  assign t[427] = (x[109]);
  assign t[428] = (x[112]);
  assign t[429] = (x[112]);
  assign t[42] = ~(t[156]);
  assign t[430] = (x[115]);
  assign t[431] = (x[115]);
  assign t[432] = (x[118]);
  assign t[433] = (x[118]);
  assign t[434] = (x[121]);
  assign t[435] = (x[121]);
  assign t[436] = (x[124]);
  assign t[437] = (x[124]);
  assign t[438] = (x[127]);
  assign t[439] = (x[127]);
  assign t[43] = ~(t[157] | t[158]);
  assign t[44] = ~(t[159] | t[160]);
  assign t[45] = t[53] ^ t[54];
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[57] & t[58];
  assign t[48] = t[59] & t[60];
  assign t[49] = t[61] & t[62];
  assign t[4] = ~(t[7]);
  assign t[50] = t[63] ^ t[64];
  assign t[51] = t[57] & t[65];
  assign t[52] = t[59] & t[66];
  assign t[53] = t[67] & t[68];
  assign t[54] = t[67] ^ t[69];
  assign t[55] = t[70] ^ t[71];
  assign t[56] = t[72] ^ t[73];
  assign t[57] = t[74] ^ t[75];
  assign t[58] = t[70] ^ t[76];
  assign t[59] = t[57] ^ t[77];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[76] ^ t[71];
  assign t[61] = t[75] ^ t[45];
  assign t[62] = t[58] ^ t[78];
  assign t[63] = t[45] & t[79];
  assign t[64] = t[61] & t[80];
  assign t[65] = t[78] ^ t[81];
  assign t[66] = t[58] ^ t[82];
  assign t[67] = t[83] ^ t[84];
  assign t[68] = t[85] & t[83];
  assign t[69] = t[83] & t[86];
  assign t[6] = ~(t[10]);
  assign t[70] = t[25] ? t[161] : t[87];
  assign t[71] = t[25] ? t[162] : t[88];
  assign t[72] = t[89] ^ t[90];
  assign t[73] = t[91] ^ t[92];
  assign t[74] = t[85] ^ t[93];
  assign t[75] = t[84] ^ t[94];
  assign t[76] = t[25] ? t[163] : t[95];
  assign t[77] = t[96] ^ t[45];
  assign t[78] = t[97] ^ t[91];
  assign t[79] = t[92] ^ t[62];
  assign t[7] = ~(t[11]);
  assign t[80] = t[98] ^ t[60];
  assign t[81] = t[89] ^ t[71];
  assign t[82] = t[90] ^ t[71];
  assign t[83] = t[99] ^ t[100];
  assign t[84] = t[101] ^ t[102];
  assign t[85] = t[103] ^ t[104];
  assign t[86] = t[105] ^ t[100];
  assign t[87] = t[164] ^ t[165];
  assign t[88] = t[166] ^ t[167];
  assign t[89] = t[25] ? t[168] : t[21];
  assign t[8] = ~(t[12]);
  assign t[90] = t[25] ? t[169] : t[106];
  assign t[91] = t[25] ? t[170] : t[107];
  assign t[92] = t[25] ? t[171] : t[108];
  assign t[93] = t[109] & t[110];
  assign t[94] = t[111] & t[67];
  assign t[95] = t[172] ^ t[173];
  assign t[96] = t[112] ^ t[113];
  assign t[97] = t[25] ? t[174] : t[114];
  assign t[98] = t[70] ^ t[91];
  assign t[99] = t[115] ^ t[116];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind550(x, y);
 input [129:0] x;
 output y;

 wire [440:0] t;
  assign t[0] = t[1] ? t[2] : t[140];
  assign t[100] = t[118] ^ t[119];
  assign t[101] = t[79] ^ t[104];
  assign t[102] = t[120] ^ t[81];
  assign t[103] = t[116] & t[81];
  assign t[104] = t[120] & t[116];
  assign t[105] = t[79] & t[120];
  assign t[106] = t[174] ^ t[175];
  assign t[107] = t[176] ^ t[177];
  assign t[108] = t[178] ^ t[179];
  assign t[109] = t[180] ^ t[181];
  assign t[10] = t[142] & t[16];
  assign t[110] = t[88] ^ t[90];
  assign t[111] = t[156] ^ t[182];
  assign t[112] = t[121] ^ t[122];
  assign t[113] = t[92] ^ t[123];
  assign t[114] = t[92] & t[123];
  assign t[115] = t[59] & t[64];
  assign t[116] = t[124] ^ t[125];
  assign t[117] = t[126] ^ t[127];
  assign t[118] = t[59] ^ t[128];
  assign t[119] = t[76] ^ t[58];
  assign t[11] = ~(t[17]);
  assign t[120] = t[129] ^ t[125];
  assign t[121] = t[128] & t[90];
  assign t[122] = t[61] & t[130];
  assign t[123] = t[130] ^ t[91];
  assign t[124] = t[131] ^ t[132];
  assign t[125] = t[133] ^ t[115];
  assign t[126] = t[118] & t[119];
  assign t[127] = t[75] & t[58];
  assign t[128] = t[91] ^ t[134];
  assign t[129] = t[135] ^ t[136];
  assign t[12] = ~(t[142]);
  assign t[130] = t[59] ^ t[72];
  assign t[131] = t[137] ^ t[122];
  assign t[132] = t[77] & t[138];
  assign t[133] = t[46] & t[65];
  assign t[134] = t[55] ^ t[90];
  assign t[135] = t[139] ^ t[127];
  assign t[136] = t[93] & t[76];
  assign t[137] = t[130] ^ t[78];
  assign t[138] = t[90] ^ t[130];
  assign t[139] = t[75] ^ t[58];
  assign t[13] = ~(t[18]);
  assign t[140] = (t[183]);
  assign t[141] = (t[184]);
  assign t[142] = (t[185]);
  assign t[143] = (t[186]);
  assign t[144] = (t[187]);
  assign t[145] = (t[188]);
  assign t[146] = (t[189]);
  assign t[147] = (t[190]);
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[19] ? t[143] : t[22];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[142] & t[24]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = (t[225]);
  assign t[183] = t[226] ^ x[2];
  assign t[184] = t[227] ^ x[5];
  assign t[185] = t[228] ^ x[9];
  assign t[186] = t[229] ^ x[12];
  assign t[187] = t[230] ^ x[15];
  assign t[188] = t[231] ^ x[18];
  assign t[189] = t[232] ^ x[21];
  assign t[18] = ~(t[25]);
  assign t[190] = t[233] ^ x[24];
  assign t[191] = t[234] ^ x[27];
  assign t[192] = t[235] ^ x[30];
  assign t[193] = t[236] ^ x[33];
  assign t[194] = t[237] ^ x[36];
  assign t[195] = t[238] ^ x[39];
  assign t[196] = t[239] ^ x[42];
  assign t[197] = t[240] ^ x[45];
  assign t[198] = t[241] ^ x[48];
  assign t[199] = t[242] ^ x[51];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[54];
  assign t[201] = t[244] ^ x[57];
  assign t[202] = t[245] ^ x[60];
  assign t[203] = t[246] ^ x[63];
  assign t[204] = t[247] ^ x[66];
  assign t[205] = t[248] ^ x[69];
  assign t[206] = t[249] ^ x[72];
  assign t[207] = t[250] ^ x[75];
  assign t[208] = t[251] ^ x[78];
  assign t[209] = t[252] ^ x[81];
  assign t[20] = t[28] ^ t[29];
  assign t[210] = t[253] ^ x[84];
  assign t[211] = t[254] ^ x[87];
  assign t[212] = t[255] ^ x[90];
  assign t[213] = t[256] ^ x[93];
  assign t[214] = t[257] ^ x[96];
  assign t[215] = t[258] ^ x[99];
  assign t[216] = t[259] ^ x[102];
  assign t[217] = t[260] ^ x[105];
  assign t[218] = t[261] ^ x[108];
  assign t[219] = t[262] ^ x[111];
  assign t[21] = t[144] ^ t[145];
  assign t[220] = t[263] ^ x[114];
  assign t[221] = t[264] ^ x[117];
  assign t[222] = t[265] ^ x[120];
  assign t[223] = t[266] ^ x[123];
  assign t[224] = t[267] ^ x[126];
  assign t[225] = t[268] ^ x[129];
  assign t[226] = (t[269] & ~t[270]);
  assign t[227] = (t[271] & ~t[272]);
  assign t[228] = (t[273] & ~t[274]);
  assign t[229] = (t[275] & ~t[276]);
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[277] & ~t[278]);
  assign t[231] = (t[279] & ~t[280]);
  assign t[232] = (t[281] & ~t[282]);
  assign t[233] = (t[283] & ~t[284]);
  assign t[234] = (t[285] & ~t[286]);
  assign t[235] = (t[287] & ~t[288]);
  assign t[236] = (t[289] & ~t[290]);
  assign t[237] = (t[291] & ~t[292]);
  assign t[238] = (t[293] & ~t[294]);
  assign t[239] = (t[295] & ~t[296]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[297] & ~t[298]);
  assign t[241] = (t[299] & ~t[300]);
  assign t[242] = (t[301] & ~t[302]);
  assign t[243] = (t[303] & ~t[304]);
  assign t[244] = (t[305] & ~t[306]);
  assign t[245] = (t[307] & ~t[308]);
  assign t[246] = (t[309] & ~t[310]);
  assign t[247] = (t[311] & ~t[312]);
  assign t[248] = (t[313] & ~t[314]);
  assign t[249] = (t[315] & ~t[316]);
  assign t[24] = ~(t[146] | t[34]);
  assign t[250] = (t[317] & ~t[318]);
  assign t[251] = (t[319] & ~t[320]);
  assign t[252] = (t[321] & ~t[322]);
  assign t[253] = (t[323] & ~t[324]);
  assign t[254] = (t[325] & ~t[326]);
  assign t[255] = (t[327] & ~t[328]);
  assign t[256] = (t[329] & ~t[330]);
  assign t[257] = (t[331] & ~t[332]);
  assign t[258] = (t[333] & ~t[334]);
  assign t[259] = (t[335] & ~t[336]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[337] & ~t[338]);
  assign t[261] = (t[339] & ~t[340]);
  assign t[262] = (t[341] & ~t[342]);
  assign t[263] = (t[343] & ~t[344]);
  assign t[264] = (t[345] & ~t[346]);
  assign t[265] = (t[347] & ~t[348]);
  assign t[266] = (t[349] & ~t[350]);
  assign t[267] = (t[351] & ~t[352]);
  assign t[268] = (t[353] & ~t[354]);
  assign t[269] = t[355] ^ x[2];
  assign t[26] = ~(t[147] & t[148]);
  assign t[270] = t[356] ^ x[1];
  assign t[271] = t[357] ^ x[5];
  assign t[272] = t[358] ^ x[4];
  assign t[273] = t[359] ^ x[9];
  assign t[274] = t[360] ^ x[8];
  assign t[275] = t[361] ^ x[12];
  assign t[276] = t[362] ^ x[11];
  assign t[277] = t[363] ^ x[15];
  assign t[278] = t[364] ^ x[14];
  assign t[279] = t[365] ^ x[18];
  assign t[27] = ~(t[149] & t[150]);
  assign t[280] = t[366] ^ x[17];
  assign t[281] = t[367] ^ x[21];
  assign t[282] = t[368] ^ x[20];
  assign t[283] = t[369] ^ x[24];
  assign t[284] = t[370] ^ x[23];
  assign t[285] = t[371] ^ x[27];
  assign t[286] = t[372] ^ x[26];
  assign t[287] = t[373] ^ x[30];
  assign t[288] = t[374] ^ x[29];
  assign t[289] = t[375] ^ x[33];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[376] ^ x[32];
  assign t[291] = t[377] ^ x[36];
  assign t[292] = t[378] ^ x[35];
  assign t[293] = t[379] ^ x[39];
  assign t[294] = t[380] ^ x[38];
  assign t[295] = t[381] ^ x[42];
  assign t[296] = t[382] ^ x[41];
  assign t[297] = t[383] ^ x[45];
  assign t[298] = t[384] ^ x[44];
  assign t[299] = t[385] ^ x[48];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[141] : t[5];
  assign t[300] = t[386] ^ x[47];
  assign t[301] = t[387] ^ x[51];
  assign t[302] = t[388] ^ x[50];
  assign t[303] = t[389] ^ x[54];
  assign t[304] = t[390] ^ x[53];
  assign t[305] = t[391] ^ x[57];
  assign t[306] = t[392] ^ x[56];
  assign t[307] = t[393] ^ x[60];
  assign t[308] = t[394] ^ x[59];
  assign t[309] = t[395] ^ x[63];
  assign t[30] = t[151] ^ t[41];
  assign t[310] = t[396] ^ x[62];
  assign t[311] = t[397] ^ x[66];
  assign t[312] = t[398] ^ x[65];
  assign t[313] = t[399] ^ x[69];
  assign t[314] = t[400] ^ x[68];
  assign t[315] = t[401] ^ x[72];
  assign t[316] = t[402] ^ x[71];
  assign t[317] = t[403] ^ x[75];
  assign t[318] = t[404] ^ x[74];
  assign t[319] = t[405] ^ x[78];
  assign t[31] = ~(t[152] ^ t[153]);
  assign t[320] = t[406] ^ x[77];
  assign t[321] = t[407] ^ x[81];
  assign t[322] = t[408] ^ x[80];
  assign t[323] = t[409] ^ x[84];
  assign t[324] = t[410] ^ x[83];
  assign t[325] = t[411] ^ x[87];
  assign t[326] = t[412] ^ x[86];
  assign t[327] = t[413] ^ x[90];
  assign t[328] = t[414] ^ x[89];
  assign t[329] = t[415] ^ x[93];
  assign t[32] = ~(t[24]);
  assign t[330] = t[416] ^ x[92];
  assign t[331] = t[417] ^ x[96];
  assign t[332] = t[418] ^ x[95];
  assign t[333] = t[419] ^ x[99];
  assign t[334] = t[420] ^ x[98];
  assign t[335] = t[421] ^ x[102];
  assign t[336] = t[422] ^ x[101];
  assign t[337] = t[423] ^ x[105];
  assign t[338] = t[424] ^ x[104];
  assign t[339] = t[425] ^ x[108];
  assign t[33] = ~(t[154] & t[42]);
  assign t[340] = t[426] ^ x[107];
  assign t[341] = t[427] ^ x[111];
  assign t[342] = t[428] ^ x[110];
  assign t[343] = t[429] ^ x[114];
  assign t[344] = t[430] ^ x[113];
  assign t[345] = t[431] ^ x[117];
  assign t[346] = t[432] ^ x[116];
  assign t[347] = t[433] ^ x[120];
  assign t[348] = t[434] ^ x[119];
  assign t[349] = t[435] ^ x[123];
  assign t[34] = ~(t[43] & t[44]);
  assign t[350] = t[436] ^ x[122];
  assign t[351] = t[437] ^ x[126];
  assign t[352] = t[438] ^ x[125];
  assign t[353] = t[439] ^ x[129];
  assign t[354] = t[440] ^ x[128];
  assign t[355] = (x[0]);
  assign t[356] = (x[0]);
  assign t[357] = (x[3]);
  assign t[358] = (x[3]);
  assign t[359] = (x[7]);
  assign t[35] = ~(t[155]);
  assign t[360] = (x[7]);
  assign t[361] = (x[10]);
  assign t[362] = (x[10]);
  assign t[363] = (x[13]);
  assign t[364] = (x[13]);
  assign t[365] = (x[16]);
  assign t[366] = (x[16]);
  assign t[367] = (x[19]);
  assign t[368] = (x[19]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[142]);
  assign t[370] = (x[22]);
  assign t[371] = (x[25]);
  assign t[372] = (x[25]);
  assign t[373] = (x[28]);
  assign t[374] = (x[28]);
  assign t[375] = (x[31]);
  assign t[376] = (x[31]);
  assign t[377] = (x[34]);
  assign t[378] = (x[34]);
  assign t[379] = (x[37]);
  assign t[37] = t[45] & t[46];
  assign t[380] = (x[37]);
  assign t[381] = (x[40]);
  assign t[382] = (x[40]);
  assign t[383] = (x[43]);
  assign t[384] = (x[43]);
  assign t[385] = (x[46]);
  assign t[386] = (x[46]);
  assign t[387] = (x[49]);
  assign t[388] = (x[49]);
  assign t[389] = (x[52]);
  assign t[38] = t[47] ^ t[48];
  assign t[390] = (x[52]);
  assign t[391] = (x[55]);
  assign t[392] = (x[55]);
  assign t[393] = (x[58]);
  assign t[394] = (x[58]);
  assign t[395] = (x[61]);
  assign t[396] = (x[61]);
  assign t[397] = (x[64]);
  assign t[398] = (x[64]);
  assign t[399] = (x[67]);
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[67]);
  assign t[401] = (x[70]);
  assign t[402] = (x[70]);
  assign t[403] = (x[73]);
  assign t[404] = (x[73]);
  assign t[405] = (x[76]);
  assign t[406] = (x[76]);
  assign t[407] = (x[79]);
  assign t[408] = (x[79]);
  assign t[409] = (x[82]);
  assign t[40] = t[51] ^ t[52];
  assign t[410] = (x[82]);
  assign t[411] = (x[85]);
  assign t[412] = (x[85]);
  assign t[413] = (x[88]);
  assign t[414] = (x[88]);
  assign t[415] = (x[91]);
  assign t[416] = (x[91]);
  assign t[417] = (x[94]);
  assign t[418] = (x[94]);
  assign t[419] = (x[97]);
  assign t[41] = t[144] ^ t[156];
  assign t[420] = (x[97]);
  assign t[421] = (x[100]);
  assign t[422] = (x[100]);
  assign t[423] = (x[103]);
  assign t[424] = (x[103]);
  assign t[425] = (x[106]);
  assign t[426] = (x[106]);
  assign t[427] = (x[109]);
  assign t[428] = (x[109]);
  assign t[429] = (x[112]);
  assign t[42] = ~(t[157]);
  assign t[430] = (x[112]);
  assign t[431] = (x[115]);
  assign t[432] = (x[115]);
  assign t[433] = (x[118]);
  assign t[434] = (x[118]);
  assign t[435] = (x[121]);
  assign t[436] = (x[121]);
  assign t[437] = (x[124]);
  assign t[438] = (x[124]);
  assign t[439] = (x[127]);
  assign t[43] = ~(t[158] | t[159]);
  assign t[440] = (x[127]);
  assign t[44] = ~(t[160] | t[161]);
  assign t[45] = t[53] ^ t[54];
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[57] & t[58];
  assign t[48] = t[53] & t[59];
  assign t[49] = t[60] & t[61];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] ^ t[63];
  assign t[51] = t[53] & t[64];
  assign t[52] = t[45] & t[65];
  assign t[53] = t[66] ^ t[67];
  assign t[54] = t[68] ^ t[69];
  assign t[55] = t[25] ? t[162] : t[70];
  assign t[56] = t[25] ? t[163] : t[71];
  assign t[57] = t[66] ^ t[68];
  assign t[58] = t[72] ^ t[73];
  assign t[59] = t[74] ^ t[55];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[67] ^ t[69];
  assign t[61] = t[75] ^ t[46];
  assign t[62] = t[68] & t[76];
  assign t[63] = t[69] & t[77];
  assign t[64] = t[72] ^ t[78];
  assign t[65] = t[59] ^ t[73];
  assign t[66] = t[79] ^ t[80];
  assign t[67] = t[81] ^ t[82];
  assign t[68] = t[83] ^ t[84];
  assign t[69] = t[85] ^ t[86];
  assign t[6] = ~(t[10]);
  assign t[70] = t[164] ^ t[165];
  assign t[71] = t[166] ^ t[167];
  assign t[72] = t[87] ^ t[88];
  assign t[73] = t[89] ^ t[56];
  assign t[74] = t[25] ? t[168] : t[21];
  assign t[75] = t[74] ^ t[88];
  assign t[76] = t[90] ^ t[91];
  assign t[77] = t[92] ^ t[93];
  assign t[78] = t[94] ^ t[56];
  assign t[79] = t[95] ^ t[96];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] & t[98];
  assign t[81] = t[99] ^ t[100];
  assign t[82] = t[101] & t[102];
  assign t[83] = t[98] & t[103];
  assign t[84] = t[98] ^ t[104];
  assign t[85] = t[102] & t[105];
  assign t[86] = t[102] ^ t[104];
  assign t[87] = t[25] ? t[169] : t[106];
  assign t[88] = t[25] ? t[170] : t[107];
  assign t[89] = t[25] ? t[171] : t[108];
  assign t[8] = ~(t[12]);
  assign t[90] = t[25] ? t[172] : t[109];
  assign t[91] = t[94] ^ t[89];
  assign t[92] = t[74] ^ t[56];
  assign t[93] = t[91] ^ t[110];
  assign t[94] = t[25] ? t[173] : t[111];
  assign t[95] = t[112] ^ t[113];
  assign t[96] = t[114] ^ t[115];
  assign t[97] = t[81] ^ t[104];
  assign t[98] = t[116] ^ t[79];
  assign t[99] = t[117] ^ t[96];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2ind551(x, y);
 input [129:0] x;
 output y;

 wire [440:0] t;
  assign t[0] = t[1] ? t[2] : t[140];
  assign t[100] = t[118] ^ t[119];
  assign t[101] = t[79] ^ t[104];
  assign t[102] = t[120] ^ t[81];
  assign t[103] = t[116] & t[81];
  assign t[104] = t[120] & t[116];
  assign t[105] = t[79] & t[120];
  assign t[106] = t[174] ^ t[175];
  assign t[107] = t[176] ^ t[177];
  assign t[108] = t[178] ^ t[179];
  assign t[109] = t[180] ^ t[181];
  assign t[10] = t[142] & t[16];
  assign t[110] = t[88] ^ t[90];
  assign t[111] = t[156] ^ t[182];
  assign t[112] = t[121] ^ t[122];
  assign t[113] = t[92] ^ t[123];
  assign t[114] = t[92] & t[123];
  assign t[115] = t[59] & t[64];
  assign t[116] = t[124] ^ t[125];
  assign t[117] = t[126] ^ t[127];
  assign t[118] = t[59] ^ t[128];
  assign t[119] = t[76] ^ t[58];
  assign t[11] = ~(t[17]);
  assign t[120] = t[129] ^ t[125];
  assign t[121] = t[128] & t[90];
  assign t[122] = t[61] & t[130];
  assign t[123] = t[130] ^ t[91];
  assign t[124] = t[131] ^ t[132];
  assign t[125] = t[133] ^ t[115];
  assign t[126] = t[118] & t[119];
  assign t[127] = t[75] & t[58];
  assign t[128] = t[91] ^ t[134];
  assign t[129] = t[135] ^ t[136];
  assign t[12] = ~(t[142]);
  assign t[130] = t[59] ^ t[72];
  assign t[131] = t[137] ^ t[122];
  assign t[132] = t[77] & t[138];
  assign t[133] = t[46] & t[65];
  assign t[134] = t[55] ^ t[90];
  assign t[135] = t[139] ^ t[127];
  assign t[136] = t[93] & t[76];
  assign t[137] = t[130] ^ t[78];
  assign t[138] = t[90] ^ t[130];
  assign t[139] = t[75] ^ t[58];
  assign t[13] = ~(t[18]);
  assign t[140] = (t[183]);
  assign t[141] = (t[184]);
  assign t[142] = (t[185]);
  assign t[143] = (t[186]);
  assign t[144] = (t[187]);
  assign t[145] = (t[188]);
  assign t[146] = (t[189]);
  assign t[147] = (t[190]);
  assign t[148] = (t[191]);
  assign t[149] = (t[192]);
  assign t[14] = t[19] ? t[21] : t[20];
  assign t[150] = (t[193]);
  assign t[151] = (t[194]);
  assign t[152] = (t[195]);
  assign t[153] = (t[196]);
  assign t[154] = (t[197]);
  assign t[155] = (t[198]);
  assign t[156] = (t[199]);
  assign t[157] = (t[200]);
  assign t[158] = (t[201]);
  assign t[159] = (t[202]);
  assign t[15] = t[19] ? t[143] : t[22];
  assign t[160] = (t[203]);
  assign t[161] = (t[204]);
  assign t[162] = (t[205]);
  assign t[163] = (t[206]);
  assign t[164] = (t[207]);
  assign t[165] = (t[208]);
  assign t[166] = (t[209]);
  assign t[167] = (t[210]);
  assign t[168] = (t[211]);
  assign t[169] = (t[212]);
  assign t[16] = t[19] & t[23];
  assign t[170] = (t[213]);
  assign t[171] = (t[214]);
  assign t[172] = (t[215]);
  assign t[173] = (t[216]);
  assign t[174] = (t[217]);
  assign t[175] = (t[218]);
  assign t[176] = (t[219]);
  assign t[177] = (t[220]);
  assign t[178] = (t[221]);
  assign t[179] = (t[222]);
  assign t[17] = ~(t[142] & t[24]);
  assign t[180] = (t[223]);
  assign t[181] = (t[224]);
  assign t[182] = (t[225]);
  assign t[183] = t[226] ^ x[2];
  assign t[184] = t[227] ^ x[5];
  assign t[185] = t[228] ^ x[9];
  assign t[186] = t[229] ^ x[12];
  assign t[187] = t[230] ^ x[15];
  assign t[188] = t[231] ^ x[18];
  assign t[189] = t[232] ^ x[21];
  assign t[18] = ~(t[25]);
  assign t[190] = t[233] ^ x[24];
  assign t[191] = t[234] ^ x[27];
  assign t[192] = t[235] ^ x[30];
  assign t[193] = t[236] ^ x[33];
  assign t[194] = t[237] ^ x[36];
  assign t[195] = t[238] ^ x[39];
  assign t[196] = t[239] ^ x[42];
  assign t[197] = t[240] ^ x[45];
  assign t[198] = t[241] ^ x[48];
  assign t[199] = t[242] ^ x[51];
  assign t[19] = ~(t[26] | t[27]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[54];
  assign t[201] = t[244] ^ x[57];
  assign t[202] = t[245] ^ x[60];
  assign t[203] = t[246] ^ x[63];
  assign t[204] = t[247] ^ x[66];
  assign t[205] = t[248] ^ x[69];
  assign t[206] = t[249] ^ x[72];
  assign t[207] = t[250] ^ x[75];
  assign t[208] = t[251] ^ x[78];
  assign t[209] = t[252] ^ x[81];
  assign t[20] = t[28] ^ t[29];
  assign t[210] = t[253] ^ x[84];
  assign t[211] = t[254] ^ x[87];
  assign t[212] = t[255] ^ x[90];
  assign t[213] = t[256] ^ x[93];
  assign t[214] = t[257] ^ x[96];
  assign t[215] = t[258] ^ x[99];
  assign t[216] = t[259] ^ x[102];
  assign t[217] = t[260] ^ x[105];
  assign t[218] = t[261] ^ x[108];
  assign t[219] = t[262] ^ x[111];
  assign t[21] = t[144] ^ t[145];
  assign t[220] = t[263] ^ x[114];
  assign t[221] = t[264] ^ x[117];
  assign t[222] = t[265] ^ x[120];
  assign t[223] = t[266] ^ x[123];
  assign t[224] = t[267] ^ x[126];
  assign t[225] = t[268] ^ x[129];
  assign t[226] = (t[269] & ~t[270]);
  assign t[227] = (t[271] & ~t[272]);
  assign t[228] = (t[273] & ~t[274]);
  assign t[229] = (t[275] & ~t[276]);
  assign t[22] = ~(t[30] ^ t[31]);
  assign t[230] = (t[277] & ~t[278]);
  assign t[231] = (t[279] & ~t[280]);
  assign t[232] = (t[281] & ~t[282]);
  assign t[233] = (t[283] & ~t[284]);
  assign t[234] = (t[285] & ~t[286]);
  assign t[235] = (t[287] & ~t[288]);
  assign t[236] = (t[289] & ~t[290]);
  assign t[237] = (t[291] & ~t[292]);
  assign t[238] = (t[293] & ~t[294]);
  assign t[239] = (t[295] & ~t[296]);
  assign t[23] = ~(t[32] | t[33]);
  assign t[240] = (t[297] & ~t[298]);
  assign t[241] = (t[299] & ~t[300]);
  assign t[242] = (t[301] & ~t[302]);
  assign t[243] = (t[303] & ~t[304]);
  assign t[244] = (t[305] & ~t[306]);
  assign t[245] = (t[307] & ~t[308]);
  assign t[246] = (t[309] & ~t[310]);
  assign t[247] = (t[311] & ~t[312]);
  assign t[248] = (t[313] & ~t[314]);
  assign t[249] = (t[315] & ~t[316]);
  assign t[24] = ~(t[146] | t[34]);
  assign t[250] = (t[317] & ~t[318]);
  assign t[251] = (t[319] & ~t[320]);
  assign t[252] = (t[321] & ~t[322]);
  assign t[253] = (t[323] & ~t[324]);
  assign t[254] = (t[325] & ~t[326]);
  assign t[255] = (t[327] & ~t[328]);
  assign t[256] = (t[329] & ~t[330]);
  assign t[257] = (t[331] & ~t[332]);
  assign t[258] = (t[333] & ~t[334]);
  assign t[259] = (t[335] & ~t[336]);
  assign t[25] = ~(t[35] | t[36]);
  assign t[260] = (t[337] & ~t[338]);
  assign t[261] = (t[339] & ~t[340]);
  assign t[262] = (t[341] & ~t[342]);
  assign t[263] = (t[343] & ~t[344]);
  assign t[264] = (t[345] & ~t[346]);
  assign t[265] = (t[347] & ~t[348]);
  assign t[266] = (t[349] & ~t[350]);
  assign t[267] = (t[351] & ~t[352]);
  assign t[268] = (t[353] & ~t[354]);
  assign t[269] = t[355] ^ x[2];
  assign t[26] = ~(t[147] & t[148]);
  assign t[270] = t[356] ^ x[1];
  assign t[271] = t[357] ^ x[5];
  assign t[272] = t[358] ^ x[4];
  assign t[273] = t[359] ^ x[9];
  assign t[274] = t[360] ^ x[8];
  assign t[275] = t[361] ^ x[12];
  assign t[276] = t[362] ^ x[11];
  assign t[277] = t[363] ^ x[15];
  assign t[278] = t[364] ^ x[14];
  assign t[279] = t[365] ^ x[18];
  assign t[27] = ~(t[149] & t[150]);
  assign t[280] = t[366] ^ x[17];
  assign t[281] = t[367] ^ x[21];
  assign t[282] = t[368] ^ x[20];
  assign t[283] = t[369] ^ x[24];
  assign t[284] = t[370] ^ x[23];
  assign t[285] = t[371] ^ x[27];
  assign t[286] = t[372] ^ x[26];
  assign t[287] = t[373] ^ x[30];
  assign t[288] = t[374] ^ x[29];
  assign t[289] = t[375] ^ x[33];
  assign t[28] = t[37] ^ t[38];
  assign t[290] = t[376] ^ x[32];
  assign t[291] = t[377] ^ x[36];
  assign t[292] = t[378] ^ x[35];
  assign t[293] = t[379] ^ x[39];
  assign t[294] = t[380] ^ x[38];
  assign t[295] = t[381] ^ x[42];
  assign t[296] = t[382] ^ x[41];
  assign t[297] = t[383] ^ x[45];
  assign t[298] = t[384] ^ x[44];
  assign t[299] = t[385] ^ x[48];
  assign t[29] = t[39] ^ t[40];
  assign t[2] = t[4] ? t[141] : t[5];
  assign t[300] = t[386] ^ x[47];
  assign t[301] = t[387] ^ x[51];
  assign t[302] = t[388] ^ x[50];
  assign t[303] = t[389] ^ x[54];
  assign t[304] = t[390] ^ x[53];
  assign t[305] = t[391] ^ x[57];
  assign t[306] = t[392] ^ x[56];
  assign t[307] = t[393] ^ x[60];
  assign t[308] = t[394] ^ x[59];
  assign t[309] = t[395] ^ x[63];
  assign t[30] = t[151] ^ t[41];
  assign t[310] = t[396] ^ x[62];
  assign t[311] = t[397] ^ x[66];
  assign t[312] = t[398] ^ x[65];
  assign t[313] = t[399] ^ x[69];
  assign t[314] = t[400] ^ x[68];
  assign t[315] = t[401] ^ x[72];
  assign t[316] = t[402] ^ x[71];
  assign t[317] = t[403] ^ x[75];
  assign t[318] = t[404] ^ x[74];
  assign t[319] = t[405] ^ x[78];
  assign t[31] = ~(t[152] ^ t[153]);
  assign t[320] = t[406] ^ x[77];
  assign t[321] = t[407] ^ x[81];
  assign t[322] = t[408] ^ x[80];
  assign t[323] = t[409] ^ x[84];
  assign t[324] = t[410] ^ x[83];
  assign t[325] = t[411] ^ x[87];
  assign t[326] = t[412] ^ x[86];
  assign t[327] = t[413] ^ x[90];
  assign t[328] = t[414] ^ x[89];
  assign t[329] = t[415] ^ x[93];
  assign t[32] = ~(t[24]);
  assign t[330] = t[416] ^ x[92];
  assign t[331] = t[417] ^ x[96];
  assign t[332] = t[418] ^ x[95];
  assign t[333] = t[419] ^ x[99];
  assign t[334] = t[420] ^ x[98];
  assign t[335] = t[421] ^ x[102];
  assign t[336] = t[422] ^ x[101];
  assign t[337] = t[423] ^ x[105];
  assign t[338] = t[424] ^ x[104];
  assign t[339] = t[425] ^ x[108];
  assign t[33] = ~(t[154] & t[42]);
  assign t[340] = t[426] ^ x[107];
  assign t[341] = t[427] ^ x[111];
  assign t[342] = t[428] ^ x[110];
  assign t[343] = t[429] ^ x[114];
  assign t[344] = t[430] ^ x[113];
  assign t[345] = t[431] ^ x[117];
  assign t[346] = t[432] ^ x[116];
  assign t[347] = t[433] ^ x[120];
  assign t[348] = t[434] ^ x[119];
  assign t[349] = t[435] ^ x[123];
  assign t[34] = ~(t[43] & t[44]);
  assign t[350] = t[436] ^ x[122];
  assign t[351] = t[437] ^ x[126];
  assign t[352] = t[438] ^ x[125];
  assign t[353] = t[439] ^ x[129];
  assign t[354] = t[440] ^ x[128];
  assign t[355] = (x[0]);
  assign t[356] = (x[0]);
  assign t[357] = (x[3]);
  assign t[358] = (x[3]);
  assign t[359] = (x[7]);
  assign t[35] = ~(t[155]);
  assign t[360] = (x[7]);
  assign t[361] = (x[10]);
  assign t[362] = (x[10]);
  assign t[363] = (x[13]);
  assign t[364] = (x[13]);
  assign t[365] = (x[16]);
  assign t[366] = (x[16]);
  assign t[367] = (x[19]);
  assign t[368] = (x[19]);
  assign t[369] = (x[22]);
  assign t[36] = ~(t[142]);
  assign t[370] = (x[22]);
  assign t[371] = (x[25]);
  assign t[372] = (x[25]);
  assign t[373] = (x[28]);
  assign t[374] = (x[28]);
  assign t[375] = (x[31]);
  assign t[376] = (x[31]);
  assign t[377] = (x[34]);
  assign t[378] = (x[34]);
  assign t[379] = (x[37]);
  assign t[37] = t[45] & t[46];
  assign t[380] = (x[37]);
  assign t[381] = (x[40]);
  assign t[382] = (x[40]);
  assign t[383] = (x[43]);
  assign t[384] = (x[43]);
  assign t[385] = (x[46]);
  assign t[386] = (x[46]);
  assign t[387] = (x[49]);
  assign t[388] = (x[49]);
  assign t[389] = (x[52]);
  assign t[38] = t[47] ^ t[48];
  assign t[390] = (x[52]);
  assign t[391] = (x[55]);
  assign t[392] = (x[55]);
  assign t[393] = (x[58]);
  assign t[394] = (x[58]);
  assign t[395] = (x[61]);
  assign t[396] = (x[61]);
  assign t[397] = (x[64]);
  assign t[398] = (x[64]);
  assign t[399] = (x[67]);
  assign t[39] = t[49] ^ t[50];
  assign t[3] = ~(t[6]);
  assign t[400] = (x[67]);
  assign t[401] = (x[70]);
  assign t[402] = (x[70]);
  assign t[403] = (x[73]);
  assign t[404] = (x[73]);
  assign t[405] = (x[76]);
  assign t[406] = (x[76]);
  assign t[407] = (x[79]);
  assign t[408] = (x[79]);
  assign t[409] = (x[82]);
  assign t[40] = t[51] ^ t[52];
  assign t[410] = (x[82]);
  assign t[411] = (x[85]);
  assign t[412] = (x[85]);
  assign t[413] = (x[88]);
  assign t[414] = (x[88]);
  assign t[415] = (x[91]);
  assign t[416] = (x[91]);
  assign t[417] = (x[94]);
  assign t[418] = (x[94]);
  assign t[419] = (x[97]);
  assign t[41] = t[144] ^ t[156];
  assign t[420] = (x[97]);
  assign t[421] = (x[100]);
  assign t[422] = (x[100]);
  assign t[423] = (x[103]);
  assign t[424] = (x[103]);
  assign t[425] = (x[106]);
  assign t[426] = (x[106]);
  assign t[427] = (x[109]);
  assign t[428] = (x[109]);
  assign t[429] = (x[112]);
  assign t[42] = ~(t[157]);
  assign t[430] = (x[112]);
  assign t[431] = (x[115]);
  assign t[432] = (x[115]);
  assign t[433] = (x[118]);
  assign t[434] = (x[118]);
  assign t[435] = (x[121]);
  assign t[436] = (x[121]);
  assign t[437] = (x[124]);
  assign t[438] = (x[124]);
  assign t[439] = (x[127]);
  assign t[43] = ~(t[158] | t[159]);
  assign t[440] = (x[127]);
  assign t[44] = ~(t[160] | t[161]);
  assign t[45] = t[53] ^ t[54];
  assign t[46] = t[55] ^ t[56];
  assign t[47] = t[57] & t[58];
  assign t[48] = t[53] & t[59];
  assign t[49] = t[60] & t[61];
  assign t[4] = ~(t[7]);
  assign t[50] = t[62] ^ t[63];
  assign t[51] = t[53] & t[64];
  assign t[52] = t[45] & t[65];
  assign t[53] = t[66] ^ t[67];
  assign t[54] = t[68] ^ t[69];
  assign t[55] = t[25] ? t[162] : t[70];
  assign t[56] = t[25] ? t[163] : t[71];
  assign t[57] = t[66] ^ t[68];
  assign t[58] = t[72] ^ t[73];
  assign t[59] = t[74] ^ t[55];
  assign t[5] = t[8] ? t[9] : x[6];
  assign t[60] = t[67] ^ t[69];
  assign t[61] = t[75] ^ t[46];
  assign t[62] = t[68] & t[76];
  assign t[63] = t[69] & t[77];
  assign t[64] = t[72] ^ t[78];
  assign t[65] = t[59] ^ t[73];
  assign t[66] = t[79] ^ t[80];
  assign t[67] = t[81] ^ t[82];
  assign t[68] = t[83] ^ t[84];
  assign t[69] = t[85] ^ t[86];
  assign t[6] = ~(t[10]);
  assign t[70] = t[164] ^ t[165];
  assign t[71] = t[166] ^ t[167];
  assign t[72] = t[87] ^ t[88];
  assign t[73] = t[89] ^ t[56];
  assign t[74] = t[25] ? t[168] : t[21];
  assign t[75] = t[74] ^ t[88];
  assign t[76] = t[90] ^ t[91];
  assign t[77] = t[92] ^ t[93];
  assign t[78] = t[94] ^ t[56];
  assign t[79] = t[95] ^ t[96];
  assign t[7] = ~(t[11]);
  assign t[80] = t[97] & t[98];
  assign t[81] = t[99] ^ t[100];
  assign t[82] = t[101] & t[102];
  assign t[83] = t[98] & t[103];
  assign t[84] = t[98] ^ t[104];
  assign t[85] = t[102] & t[105];
  assign t[86] = t[102] ^ t[104];
  assign t[87] = t[25] ? t[169] : t[106];
  assign t[88] = t[25] ? t[170] : t[107];
  assign t[89] = t[25] ? t[171] : t[108];
  assign t[8] = ~(t[12]);
  assign t[90] = t[25] ? t[172] : t[109];
  assign t[91] = t[94] ^ t[89];
  assign t[92] = t[74] ^ t[56];
  assign t[93] = t[91] ^ t[110];
  assign t[94] = t[25] ? t[173] : t[111];
  assign t[95] = t[112] ^ t[113];
  assign t[96] = t[114] ^ t[115];
  assign t[97] = t[81] ^ t[104];
  assign t[98] = t[116] ^ t[79];
  assign t[99] = t[117] ^ t[96];
  assign t[9] = t[13] ? t[15] : t[14];
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [1081:0] x;
 output [551:0] y;

  R2ind0 R2ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[2], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x(x[39]), .y(y[4]));
  R2ind5 R2ind5_inst(.x(x[39]), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[26], x[25], x[24], x[23], x[22], x[21], x[5], x[4], x[3], x[42], x[41], x[40]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[26], x[25], x[24], x[23], x[22], x[21], x[5], x[4], x[3], x[42], x[41], x[40]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[48], x[47], x[46], x[45], x[44], x[43], x[5], x[4], x[3]}), .y(y[10]));
  R2ind11 R2ind11_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[48], x[47], x[46], x[45], x[44], x[43], x[5], x[4], x[3]}), .y(y[11]));
  R2ind12 R2ind12_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[11], x[10], x[9], x[45], x[44], x[43]}), .y(y[12]));
  R2ind13 R2ind13_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[11], x[10], x[9], x[45], x[44], x[43]}), .y(y[13]));
  R2ind14 R2ind14_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[14], x[13], x[12], x[11], x[10], x[9]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[14], x[13], x[12], x[11], x[10], x[9]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[48], x[47], x[46], x[51], x[50], x[49], x[14], x[13], x[12]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[48], x[47], x[46], x[51], x[50], x[49], x[14], x[13], x[12]}), .y(y[17]));
  R2ind18 R2ind18_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[51], x[50], x[49], x[17], x[16], x[15], x[48], x[47], x[46], x[5], x[4], x[3]}), .y(y[18]));
  R2ind19 R2ind19_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[51], x[50], x[49], x[17], x[16], x[15], x[48], x[47], x[46], x[5], x[4], x[3]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[23], x[22], x[21], x[17], x[16], x[15], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[20]));
  R2ind21 R2ind21_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[23], x[22], x[21], x[17], x[16], x[15], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[23], x[22], x[21], x[5], x[4], x[3], x[48], x[47], x[46], x[54], x[53], x[52], x[8], x[7], x[6]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[23], x[22], x[21], x[5], x[4], x[3], x[48], x[47], x[46], x[54], x[53], x[52], x[8], x[7], x[6]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[54], x[53], x[52], x[48], x[47], x[46], x[5], x[4], x[3]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[54], x[53], x[52], x[48], x[47], x[46], x[5], x[4], x[3]}), .y(y[25]));
  R2ind26 R2ind26_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[26], x[25], x[24], x[5], x[4], x[3], x[20], x[19], x[18]}), .y(y[26]));
  R2ind27 R2ind27_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[26], x[25], x[24], x[5], x[4], x[3], x[20], x[19], x[18]}), .y(y[27]));
  R2ind28 R2ind28_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[20], x[19], x[18], x[26], x[25], x[24]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[20], x[19], x[18], x[26], x[25], x[24]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[35], x[34], x[33], x[32], x[31], x[30], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[5], x[4], x[3], x[29], x[28], x[27]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[35], x[34], x[33], x[32], x[31], x[30], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[5], x[4], x[3], x[29], x[28], x[27]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[29], x[28], x[27], x[5], x[4], x[3], x[23], x[22], x[21]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[29], x[28], x[27], x[5], x[4], x[3], x[23], x[22], x[21]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[38], x[37], x[36], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[35], x[34], x[33]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[38], x[37], x[36], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[35], x[34], x[33]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[38], x[37], x[36], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[35], x[34], x[33], x[5], x[4], x[3], x[32], x[31], x[30]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[38], x[37], x[36], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[35], x[34], x[33], x[5], x[4], x[3], x[32], x[31], x[30]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[35], x[34], x[33], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[32], x[31], x[30], x[5], x[4], x[3], x[38], x[37], x[36]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[35], x[34], x[33], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[32], x[31], x[30], x[5], x[4], x[3], x[38], x[37], x[36]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[85]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[104], x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[124], x[123], x[122], x[121], x[120], x[119], x[118], x[117], x[116], x[115]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[51], x[50], x[49], x[54], x[53], x[52], x[45], x[44], x[43], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[48], x[47], x[46], x[17], x[16], x[15], x[8], x[7], x[6], x[20], x[19], x[18], x[26], x[25], x[24], x[11], x[10], x[9], x[14], x[13], x[12], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[64], x[63], x[62]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[141], x[140], x[139], x[138], x[137], x[136], x[135], x[64], x[63], x[62]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[74], x[73], x[72]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[74], x[73], x[72]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[84], x[83], x[82]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[155], x[154], x[153], x[152], x[151], x[150], x[149], x[84], x[83], x[82]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[94], x[93], x[92]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[94], x[93], x[92]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[104], x[103], x[102]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[104], x[103], x[102]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[114], x[113], x[112]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[176], x[175], x[174], x[173], x[172], x[171], x[170], x[114], x[113], x[112]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[124], x[123], x[122]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[124], x[123], x[122]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[134], x[133], x[132]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[190], x[189], x[188], x[187], x[186], x[185], x[184], x[134], x[133], x[132]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[141], x[140], x[139]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[141], x[140], x[139]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[148], x[147], x[146]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[148], x[147], x[146]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[155], x[154], x[153]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[155], x[154], x[153]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[162], x[161], x[160]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[162], x[161], x[160]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[169], x[168], x[167]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[225], x[224], x[223], x[222], x[221], x[220], x[219], x[169], x[168], x[167]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[176], x[175], x[174]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[176], x[175], x[174]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[183], x[182], x[181]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[183], x[182], x[181]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[190], x[189], x[188]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[190], x[189], x[188]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[60], x[59], x[58], x[250], x[249], x[248], x[247], x[197], x[196], x[195]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[60], x[59], x[58], x[250], x[249], x[248], x[247], x[197], x[196], x[195]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[70], x[69], x[68], x[254], x[253], x[252], x[251], x[204], x[203], x[202]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[70], x[69], x[68], x[254], x[253], x[252], x[251], x[204], x[203], x[202]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[80], x[79], x[78], x[258], x[257], x[256], x[255], x[211], x[210], x[209]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[80], x[79], x[78], x[258], x[257], x[256], x[255], x[211], x[210], x[209]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[90], x[89], x[88], x[262], x[261], x[260], x[259], x[218], x[217], x[216]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[90], x[89], x[88], x[262], x[261], x[260], x[259], x[218], x[217], x[216]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[100], x[99], x[98], x[266], x[265], x[264], x[263], x[225], x[224], x[223]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[100], x[99], x[98], x[266], x[265], x[264], x[263], x[225], x[224], x[223]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[110], x[109], x[108], x[270], x[269], x[268], x[267], x[232], x[231], x[230]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[110], x[109], x[108], x[270], x[269], x[268], x[267], x[232], x[231], x[230]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[120], x[119], x[118], x[274], x[273], x[272], x[271], x[239], x[238], x[237]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[120], x[119], x[118], x[274], x[273], x[272], x[271], x[239], x[238], x[237]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[130], x[129], x[128], x[278], x[277], x[276], x[275], x[246], x[245], x[244]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[130], x[129], x[128], x[278], x[277], x[276], x[275], x[246], x[245], x[244]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[137], x[136], x[135], x[282], x[281], x[280], x[279], x[60], x[59], x[58]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[137], x[136], x[135], x[282], x[281], x[280], x[279], x[60], x[59], x[58]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[144], x[143], x[142], x[286], x[285], x[284], x[283], x[70], x[69], x[68]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[144], x[143], x[142], x[286], x[285], x[284], x[283], x[70], x[69], x[68]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[151], x[150], x[149], x[290], x[289], x[288], x[287], x[80], x[79], x[78]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[151], x[150], x[149], x[290], x[289], x[288], x[287], x[80], x[79], x[78]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[158], x[157], x[156], x[294], x[293], x[292], x[291], x[90], x[89], x[88]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[158], x[157], x[156], x[294], x[293], x[292], x[291], x[90], x[89], x[88]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[165], x[164], x[163], x[298], x[297], x[296], x[295], x[100], x[99], x[98]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[165], x[164], x[163], x[298], x[297], x[296], x[295], x[100], x[99], x[98]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[172], x[171], x[170], x[302], x[301], x[300], x[299], x[110], x[109], x[108]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[172], x[171], x[170], x[302], x[301], x[300], x[299], x[110], x[109], x[108]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[179], x[178], x[177], x[306], x[305], x[304], x[303], x[120], x[119], x[118]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[179], x[178], x[177], x[306], x[305], x[304], x[303], x[120], x[119], x[118]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[186], x[185], x[184], x[310], x[309], x[308], x[307], x[130], x[129], x[128]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[186], x[185], x[184], x[310], x[309], x[308], x[307], x[130], x[129], x[128]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[193], x[192], x[191], x[314], x[313], x[312], x[311], x[137], x[136], x[135]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[193], x[192], x[191], x[314], x[313], x[312], x[311], x[137], x[136], x[135]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[200], x[199], x[198], x[318], x[317], x[316], x[315], x[144], x[143], x[142]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[200], x[199], x[198], x[318], x[317], x[316], x[315], x[144], x[143], x[142]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[207], x[206], x[205], x[322], x[321], x[320], x[319], x[151], x[150], x[149]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[207], x[206], x[205], x[322], x[321], x[320], x[319], x[151], x[150], x[149]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[214], x[213], x[212], x[326], x[325], x[324], x[323], x[158], x[157], x[156]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[214], x[213], x[212], x[326], x[325], x[324], x[323], x[158], x[157], x[156]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[221], x[220], x[219], x[330], x[329], x[328], x[327], x[165], x[164], x[163]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[221], x[220], x[219], x[330], x[329], x[328], x[327], x[165], x[164], x[163]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[228], x[227], x[226], x[334], x[333], x[332], x[331], x[172], x[171], x[170]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[228], x[227], x[226], x[334], x[333], x[332], x[331], x[172], x[171], x[170]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[235], x[234], x[233], x[338], x[337], x[336], x[335], x[179], x[178], x[177]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[235], x[234], x[233], x[338], x[337], x[336], x[335], x[179], x[178], x[177]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[242], x[241], x[240], x[342], x[341], x[340], x[339], x[186], x[185], x[184]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[242], x[241], x[240], x[342], x[341], x[340], x[339], x[186], x[185], x[184]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[249], x[248], x[247], x[346], x[345], x[344], x[343], x[193], x[192], x[191]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[249], x[248], x[247], x[346], x[345], x[344], x[343], x[193], x[192], x[191]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[253], x[252], x[251], x[350], x[349], x[348], x[347], x[200], x[199], x[198]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[253], x[252], x[251], x[350], x[349], x[348], x[347], x[200], x[199], x[198]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[257], x[256], x[255], x[354], x[353], x[352], x[351], x[207], x[206], x[205]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[257], x[256], x[255], x[354], x[353], x[352], x[351], x[207], x[206], x[205]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[261], x[260], x[259], x[358], x[357], x[356], x[355], x[214], x[213], x[212]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[261], x[260], x[259], x[358], x[357], x[356], x[355], x[214], x[213], x[212]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[265], x[264], x[263], x[362], x[361], x[360], x[359], x[221], x[220], x[219]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[265], x[264], x[263], x[362], x[361], x[360], x[359], x[221], x[220], x[219]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[269], x[268], x[267], x[366], x[365], x[364], x[363], x[228], x[227], x[226]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[269], x[268], x[267], x[366], x[365], x[364], x[363], x[228], x[227], x[226]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[273], x[272], x[271], x[370], x[369], x[368], x[367], x[235], x[234], x[233]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[273], x[272], x[271], x[370], x[369], x[368], x[367], x[235], x[234], x[233]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[277], x[276], x[275], x[374], x[373], x[372], x[371], x[242], x[241], x[240]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[277], x[276], x[275], x[374], x[373], x[372], x[371], x[242], x[241], x[240]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[281], x[280], x[279], x[378], x[377], x[376], x[375], x[249], x[248], x[247]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[281], x[280], x[279], x[378], x[377], x[376], x[375], x[249], x[248], x[247]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[285], x[284], x[283], x[382], x[381], x[380], x[379], x[253], x[252], x[251]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[285], x[284], x[283], x[382], x[381], x[380], x[379], x[253], x[252], x[251]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[289], x[288], x[287], x[386], x[385], x[384], x[383], x[257], x[256], x[255]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[289], x[288], x[287], x[386], x[385], x[384], x[383], x[257], x[256], x[255]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[293], x[292], x[291], x[390], x[389], x[388], x[387], x[261], x[260], x[259]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[293], x[292], x[291], x[390], x[389], x[388], x[387], x[261], x[260], x[259]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[297], x[296], x[295], x[394], x[393], x[392], x[391], x[265], x[264], x[263]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[297], x[296], x[295], x[394], x[393], x[392], x[391], x[265], x[264], x[263]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[301], x[300], x[299], x[398], x[397], x[396], x[395], x[269], x[268], x[267]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[301], x[300], x[299], x[398], x[397], x[396], x[395], x[269], x[268], x[267]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[305], x[304], x[303], x[402], x[401], x[400], x[399], x[273], x[272], x[271]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[305], x[304], x[303], x[402], x[401], x[400], x[399], x[273], x[272], x[271]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[309], x[308], x[307], x[406], x[405], x[404], x[403], x[277], x[276], x[275]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[309], x[308], x[307], x[406], x[405], x[404], x[403], x[277], x[276], x[275]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[313], x[312], x[311], x[410], x[409], x[408], x[407], x[281], x[280], x[279]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[313], x[312], x[311], x[410], x[409], x[408], x[407], x[281], x[280], x[279]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[317], x[316], x[315], x[414], x[413], x[412], x[411], x[285], x[284], x[283]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[317], x[316], x[315], x[414], x[413], x[412], x[411], x[285], x[284], x[283]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[321], x[320], x[319], x[418], x[417], x[416], x[415], x[289], x[288], x[287]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[321], x[320], x[319], x[418], x[417], x[416], x[415], x[289], x[288], x[287]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[325], x[324], x[323], x[422], x[421], x[420], x[419], x[293], x[292], x[291]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[325], x[324], x[323], x[422], x[421], x[420], x[419], x[293], x[292], x[291]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[329], x[328], x[327], x[426], x[425], x[424], x[423], x[297], x[296], x[295]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[329], x[328], x[327], x[426], x[425], x[424], x[423], x[297], x[296], x[295]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[333], x[332], x[331], x[430], x[429], x[428], x[427], x[301], x[300], x[299]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[333], x[332], x[331], x[430], x[429], x[428], x[427], x[301], x[300], x[299]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[337], x[336], x[335], x[434], x[433], x[432], x[431], x[305], x[304], x[303]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[337], x[336], x[335], x[434], x[433], x[432], x[431], x[305], x[304], x[303]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[341], x[340], x[339], x[438], x[437], x[436], x[435], x[309], x[308], x[307]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[341], x[340], x[339], x[438], x[437], x[436], x[435], x[309], x[308], x[307]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[345], x[344], x[343], x[442], x[441], x[440], x[439], x[313], x[312], x[311]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[345], x[344], x[343], x[442], x[441], x[440], x[439], x[313], x[312], x[311]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[349], x[348], x[347], x[446], x[445], x[444], x[443], x[317], x[316], x[315]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[349], x[348], x[347], x[446], x[445], x[444], x[443], x[317], x[316], x[315]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[353], x[352], x[351], x[450], x[449], x[448], x[447], x[321], x[320], x[319]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[353], x[352], x[351], x[450], x[449], x[448], x[447], x[321], x[320], x[319]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[357], x[356], x[355], x[454], x[453], x[452], x[451], x[325], x[324], x[323]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[357], x[356], x[355], x[454], x[453], x[452], x[451], x[325], x[324], x[323]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[361], x[360], x[359], x[458], x[457], x[456], x[455], x[329], x[328], x[327]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[361], x[360], x[359], x[458], x[457], x[456], x[455], x[329], x[328], x[327]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[365], x[364], x[363], x[462], x[461], x[460], x[459], x[333], x[332], x[331]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[365], x[364], x[363], x[462], x[461], x[460], x[459], x[333], x[332], x[331]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[369], x[368], x[367], x[466], x[465], x[464], x[463], x[337], x[336], x[335]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[369], x[368], x[367], x[466], x[465], x[464], x[463], x[337], x[336], x[335]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[373], x[372], x[371], x[470], x[469], x[468], x[467], x[341], x[340], x[339]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[373], x[372], x[371], x[470], x[469], x[468], x[467], x[341], x[340], x[339]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[377], x[376], x[375], x[474], x[473], x[472], x[471], x[345], x[344], x[343]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[377], x[376], x[375], x[474], x[473], x[472], x[471], x[345], x[344], x[343]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[381], x[380], x[379], x[478], x[477], x[476], x[475], x[349], x[348], x[347]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[381], x[380], x[379], x[478], x[477], x[476], x[475], x[349], x[348], x[347]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[385], x[384], x[383], x[482], x[481], x[480], x[479], x[353], x[352], x[351]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[385], x[384], x[383], x[482], x[481], x[480], x[479], x[353], x[352], x[351]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[389], x[388], x[387], x[486], x[485], x[484], x[483], x[357], x[356], x[355]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[389], x[388], x[387], x[486], x[485], x[484], x[483], x[357], x[356], x[355]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[393], x[392], x[391], x[490], x[489], x[488], x[487], x[361], x[360], x[359]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[393], x[392], x[391], x[490], x[489], x[488], x[487], x[361], x[360], x[359]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[397], x[396], x[395], x[494], x[493], x[492], x[491], x[365], x[364], x[363]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[397], x[396], x[395], x[494], x[493], x[492], x[491], x[365], x[364], x[363]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[401], x[400], x[399], x[498], x[497], x[496], x[495], x[369], x[368], x[367]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[401], x[400], x[399], x[498], x[497], x[496], x[495], x[369], x[368], x[367]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[405], x[404], x[403], x[502], x[501], x[500], x[499], x[373], x[372], x[371]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[405], x[404], x[403], x[502], x[501], x[500], x[499], x[373], x[372], x[371]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[409], x[408], x[407], x[506], x[505], x[504], x[503], x[377], x[376], x[375]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[409], x[408], x[407], x[506], x[505], x[504], x[503], x[377], x[376], x[375]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[413], x[412], x[411], x[510], x[509], x[508], x[507], x[381], x[380], x[379]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[413], x[412], x[411], x[510], x[509], x[508], x[507], x[381], x[380], x[379]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[417], x[416], x[415], x[514], x[513], x[512], x[511], x[385], x[384], x[383]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[417], x[416], x[415], x[514], x[513], x[512], x[511], x[385], x[384], x[383]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[421], x[420], x[419], x[518], x[517], x[516], x[515], x[389], x[388], x[387]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[421], x[420], x[419], x[518], x[517], x[516], x[515], x[389], x[388], x[387]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[425], x[424], x[423], x[522], x[521], x[520], x[519], x[393], x[392], x[391]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[425], x[424], x[423], x[522], x[521], x[520], x[519], x[393], x[392], x[391]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[429], x[428], x[427], x[526], x[525], x[524], x[523], x[397], x[396], x[395]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[429], x[428], x[427], x[526], x[525], x[524], x[523], x[397], x[396], x[395]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[433], x[432], x[431], x[530], x[529], x[528], x[527], x[401], x[400], x[399]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[433], x[432], x[431], x[530], x[529], x[528], x[527], x[401], x[400], x[399]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[437], x[436], x[435], x[534], x[533], x[532], x[531], x[405], x[404], x[403]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[437], x[436], x[435], x[534], x[533], x[532], x[531], x[405], x[404], x[403]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[273], x[272], x[271], x[107], x[106], x[105], x[559], x[558], x[557], x[87], x[86], x[85], x[556], x[555], x[554], x[67], x[66], x[65], x[553], x[552], x[551], x[127], x[126], x[125], x[550], x[549], x[548], x[269], x[268], x[267], x[261], x[260], x[259], x[547], x[546], x[545], x[253], x[252], x[251], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[54], x[53], x[52], x[42], x[41], x[40], x[5], x[4], x[3], x[57], x[56], x[55], x[441], x[440], x[439], x[535], x[409], x[408], x[407]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[273], x[272], x[271], x[107], x[106], x[105], x[559], x[558], x[557], x[87], x[86], x[85], x[556], x[555], x[554], x[67], x[66], x[65], x[553], x[552], x[551], x[127], x[126], x[125], x[550], x[549], x[548], x[269], x[268], x[267], x[261], x[260], x[259], x[547], x[546], x[545], x[253], x[252], x[251], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[54], x[53], x[52], x[42], x[41], x[40], x[5], x[4], x[3], x[57], x[56], x[55], x[441], x[440], x[439], x[535], x[409], x[408], x[407]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[553], x[552], x[551], x[261], x[260], x[259], x[253], x[252], x[251], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[127], x[126], x[125], x[550], x[549], x[548], x[107], x[106], x[105], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[257], x[256], x[255], x[265], x[264], x[263], x[277], x[276], x[275], x[269], x[268], x[267], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[249], x[248], x[247], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[23], x[22], x[21], x[538], x[537], x[536], x[8], x[7], x[6], x[42], x[41], x[40], x[5], x[4], x[3], x[67], x[66], x[65], x[445], x[444], x[443], x[563], x[413], x[412], x[411]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[553], x[552], x[551], x[261], x[260], x[259], x[253], x[252], x[251], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[127], x[126], x[125], x[550], x[549], x[548], x[107], x[106], x[105], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[257], x[256], x[255], x[265], x[264], x[263], x[277], x[276], x[275], x[269], x[268], x[267], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[249], x[248], x[247], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[23], x[22], x[21], x[538], x[537], x[536], x[8], x[7], x[6], x[42], x[41], x[40], x[5], x[4], x[3], x[67], x[66], x[65], x[445], x[444], x[443], x[563], x[413], x[412], x[411]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[117], x[116], x[115], x[562], x[561], x[560], x[67], x[66], x[65], x[553], x[552], x[551], x[107], x[106], x[105], x[559], x[558], x[557], x[127], x[126], x[125], x[550], x[549], x[548], x[261], x[260], x[259], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[253], x[252], x[251], x[269], x[268], x[267], x[277], x[276], x[275], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[17], x[16], x[15], x[42], x[41], x[40], x[5], x[4], x[3], x[77], x[76], x[75], x[449], x[448], x[447], x[564], x[417], x[416], x[415]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[117], x[116], x[115], x[562], x[561], x[560], x[67], x[66], x[65], x[553], x[552], x[551], x[107], x[106], x[105], x[559], x[558], x[557], x[127], x[126], x[125], x[550], x[549], x[548], x[261], x[260], x[259], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[253], x[252], x[251], x[269], x[268], x[267], x[277], x[276], x[275], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[17], x[16], x[15], x[42], x[41], x[40], x[5], x[4], x[3], x[77], x[76], x[75], x[449], x[448], x[447], x[564], x[417], x[416], x[415]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[556], x[555], x[554], x[67], x[66], x[65], x[553], x[552], x[551], x[261], x[260], x[259], x[107], x[106], x[105], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[253], x[252], x[251], x[269], x[268], x[267], x[273], x[272], x[271], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[127], x[126], x[125], x[550], x[549], x[548], x[57], x[56], x[55], x[547], x[546], x[545], x[257], x[256], x[255], x[265], x[264], x[263], x[277], x[276], x[275], x[249], x[248], x[247], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[51], x[50], x[49], x[42], x[41], x[40], x[5], x[4], x[3], x[87], x[86], x[85], x[453], x[452], x[451], x[565], x[421], x[420], x[419]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[556], x[555], x[554], x[67], x[66], x[65], x[553], x[552], x[551], x[261], x[260], x[259], x[107], x[106], x[105], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[253], x[252], x[251], x[269], x[268], x[267], x[273], x[272], x[271], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[127], x[126], x[125], x[550], x[549], x[548], x[57], x[56], x[55], x[547], x[546], x[545], x[257], x[256], x[255], x[265], x[264], x[263], x[277], x[276], x[275], x[249], x[248], x[247], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[51], x[50], x[49], x[42], x[41], x[40], x[5], x[4], x[3], x[87], x[86], x[85], x[453], x[452], x[451], x[565], x[421], x[420], x[419]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[107], x[106], x[105], x[559], x[558], x[557], x[67], x[66], x[65], x[553], x[552], x[551], x[87], x[86], x[85], x[556], x[555], x[554], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[127], x[126], x[125], x[550], x[549], x[548], x[269], x[268], x[267], x[253], x[252], x[251], x[261], x[260], x[259], x[249], x[248], x[247], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[541], x[540], x[539], x[257], x[256], x[255], x[265], x[264], x[263], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[538], x[537], x[536], x[14], x[13], x[12], x[5], x[4], x[3], x[97], x[96], x[95], x[457], x[456], x[455], x[566], x[425], x[424], x[423]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[107], x[106], x[105], x[559], x[558], x[557], x[67], x[66], x[65], x[553], x[552], x[551], x[87], x[86], x[85], x[556], x[555], x[554], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[127], x[126], x[125], x[550], x[549], x[548], x[269], x[268], x[267], x[253], x[252], x[251], x[261], x[260], x[259], x[249], x[248], x[247], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[541], x[540], x[539], x[257], x[256], x[255], x[265], x[264], x[263], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[538], x[537], x[536], x[14], x[13], x[12], x[5], x[4], x[3], x[97], x[96], x[95], x[457], x[456], x[455], x[566], x[425], x[424], x[423]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[97], x[96], x[95], x[541], x[540], x[539], x[261], x[260], x[259], x[57], x[56], x[55], x[547], x[546], x[545], x[67], x[66], x[65], x[553], x[552], x[551], x[269], x[268], x[267], x[273], x[272], x[271], x[265], x[264], x[263], x[249], x[248], x[247], x[253], x[252], x[251], x[77], x[76], x[75], x[544], x[543], x[542], x[127], x[126], x[125], x[550], x[549], x[548], x[257], x[256], x[255], x[277], x[276], x[275], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[538], x[537], x[536], x[11], x[10], x[9], x[5], x[4], x[3], x[107], x[106], x[105], x[461], x[460], x[459], x[567], x[429], x[428], x[427]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[97], x[96], x[95], x[541], x[540], x[539], x[261], x[260], x[259], x[57], x[56], x[55], x[547], x[546], x[545], x[67], x[66], x[65], x[553], x[552], x[551], x[269], x[268], x[267], x[273], x[272], x[271], x[265], x[264], x[263], x[249], x[248], x[247], x[253], x[252], x[251], x[77], x[76], x[75], x[544], x[543], x[542], x[127], x[126], x[125], x[550], x[549], x[548], x[257], x[256], x[255], x[277], x[276], x[275], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[538], x[537], x[536], x[11], x[10], x[9], x[5], x[4], x[3], x[107], x[106], x[105], x[461], x[460], x[459], x[567], x[429], x[428], x[427]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[57], x[56], x[55], x[547], x[546], x[545], x[67], x[66], x[65], x[553], x[552], x[551], x[107], x[106], x[105], x[559], x[558], x[557], x[562], x[561], x[560], x[261], x[260], x[259], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[253], x[252], x[251], x[269], x[268], x[267], x[273], x[272], x[271], x[77], x[76], x[75], x[544], x[543], x[542], x[127], x[126], x[125], x[550], x[549], x[548], x[265], x[264], x[263], x[257], x[256], x[255], x[277], x[276], x[275], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[45], x[44], x[43], x[42], x[41], x[40], x[5], x[4], x[3], x[117], x[116], x[115], x[465], x[464], x[463], x[568], x[433], x[432], x[431]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[57], x[56], x[55], x[547], x[546], x[545], x[67], x[66], x[65], x[553], x[552], x[551], x[107], x[106], x[105], x[559], x[558], x[557], x[562], x[561], x[560], x[261], x[260], x[259], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[253], x[252], x[251], x[269], x[268], x[267], x[273], x[272], x[271], x[77], x[76], x[75], x[544], x[543], x[542], x[127], x[126], x[125], x[550], x[549], x[548], x[265], x[264], x[263], x[257], x[256], x[255], x[277], x[276], x[275], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[45], x[44], x[43], x[42], x[41], x[40], x[5], x[4], x[3], x[117], x[116], x[115], x[465], x[464], x[463], x[568], x[433], x[432], x[431]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[57], x[56], x[55], x[547], x[546], x[545], x[107], x[106], x[105], x[559], x[558], x[557], x[67], x[66], x[65], x[553], x[552], x[551], x[87], x[86], x[85], x[556], x[555], x[554], x[273], x[272], x[271], x[249], x[248], x[247], x[550], x[549], x[548], x[269], x[268], x[267], x[253], x[252], x[251], x[261], x[260], x[259], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[257], x[256], x[255], x[265], x[264], x[263], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[48], x[47], x[46], x[42], x[41], x[40], x[5], x[4], x[3], x[127], x[126], x[125], x[469], x[468], x[467], x[569], x[437], x[436], x[435]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[57], x[56], x[55], x[547], x[546], x[545], x[107], x[106], x[105], x[559], x[558], x[557], x[67], x[66], x[65], x[553], x[552], x[551], x[87], x[86], x[85], x[556], x[555], x[554], x[273], x[272], x[271], x[249], x[248], x[247], x[550], x[549], x[548], x[269], x[268], x[267], x[253], x[252], x[251], x[261], x[260], x[259], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[257], x[256], x[255], x[265], x[264], x[263], x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[538], x[537], x[536], x[48], x[47], x[46], x[42], x[41], x[40], x[5], x[4], x[3], x[127], x[126], x[125], x[469], x[468], x[467], x[569], x[437], x[436], x[435]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[473], x[472], x[471], x[570], x[64], x[63], x[62], x[441], x[440], x[439]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[473], x[472], x[471], x[570], x[64], x[63], x[62], x[441], x[440], x[439]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[477], x[476], x[475], x[571], x[74], x[73], x[72], x[445], x[444], x[443]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[477], x[476], x[475], x[571], x[74], x[73], x[72], x[445], x[444], x[443]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[481], x[480], x[479], x[572], x[84], x[83], x[82], x[449], x[448], x[447]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[481], x[480], x[479], x[572], x[84], x[83], x[82], x[449], x[448], x[447]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[485], x[484], x[483], x[573], x[94], x[93], x[92], x[453], x[452], x[451]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[485], x[484], x[483], x[573], x[94], x[93], x[92], x[453], x[452], x[451]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[489], x[488], x[487], x[574], x[104], x[103], x[102], x[457], x[456], x[455]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[489], x[488], x[487], x[574], x[104], x[103], x[102], x[457], x[456], x[455]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[493], x[492], x[491], x[575], x[114], x[113], x[112], x[461], x[460], x[459]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[493], x[492], x[491], x[575], x[114], x[113], x[112], x[461], x[460], x[459]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[497], x[496], x[495], x[576], x[124], x[123], x[122], x[465], x[464], x[463]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[497], x[496], x[495], x[576], x[124], x[123], x[122], x[465], x[464], x[463]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[501], x[500], x[499], x[577], x[134], x[133], x[132], x[469], x[468], x[467]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[501], x[500], x[499], x[577], x[134], x[133], x[132], x[469], x[468], x[467]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[505], x[504], x[503], x[578], x[141], x[140], x[139], x[473], x[472], x[471]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[505], x[504], x[503], x[578], x[141], x[140], x[139], x[473], x[472], x[471]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[509], x[508], x[507], x[579], x[148], x[147], x[146], x[477], x[476], x[475]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[509], x[508], x[507], x[579], x[148], x[147], x[146], x[477], x[476], x[475]}), .y(y[267]));
  R2ind268 R2ind268_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[513], x[512], x[511], x[580], x[155], x[154], x[153], x[481], x[480], x[479]}), .y(y[268]));
  R2ind269 R2ind269_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[513], x[512], x[511], x[580], x[155], x[154], x[153], x[481], x[480], x[479]}), .y(y[269]));
  R2ind270 R2ind270_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[517], x[516], x[515], x[581], x[162], x[161], x[160], x[485], x[484], x[483]}), .y(y[270]));
  R2ind271 R2ind271_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[517], x[516], x[515], x[581], x[162], x[161], x[160], x[485], x[484], x[483]}), .y(y[271]));
  R2ind272 R2ind272_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[521], x[520], x[519], x[582], x[169], x[168], x[167], x[489], x[488], x[487]}), .y(y[272]));
  R2ind273 R2ind273_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[521], x[520], x[519], x[582], x[169], x[168], x[167], x[489], x[488], x[487]}), .y(y[273]));
  R2ind274 R2ind274_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[525], x[524], x[523], x[583], x[176], x[175], x[174], x[493], x[492], x[491]}), .y(y[274]));
  R2ind275 R2ind275_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[525], x[524], x[523], x[583], x[176], x[175], x[174], x[493], x[492], x[491]}), .y(y[275]));
  R2ind276 R2ind276_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[529], x[528], x[527], x[584], x[183], x[182], x[181], x[497], x[496], x[495]}), .y(y[276]));
  R2ind277 R2ind277_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[529], x[528], x[527], x[584], x[183], x[182], x[181], x[497], x[496], x[495]}), .y(y[277]));
  R2ind278 R2ind278_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[533], x[532], x[531], x[585], x[190], x[189], x[188], x[501], x[500], x[499]}), .y(y[278]));
  R2ind279 R2ind279_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[533], x[532], x[531], x[585], x[190], x[189], x[188], x[501], x[500], x[499]}), .y(y[279]));
  R2ind280 R2ind280_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[57], x[56], x[55], x[586], x[197], x[196], x[195], x[505], x[504], x[503]}), .y(y[280]));
  R2ind281 R2ind281_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[57], x[56], x[55], x[586], x[197], x[196], x[195], x[505], x[504], x[503]}), .y(y[281]));
  R2ind282 R2ind282_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[67], x[66], x[65], x[587], x[204], x[203], x[202], x[509], x[508], x[507]}), .y(y[282]));
  R2ind283 R2ind283_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[67], x[66], x[65], x[587], x[204], x[203], x[202], x[509], x[508], x[507]}), .y(y[283]));
  R2ind284 R2ind284_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[77], x[76], x[75], x[588], x[211], x[210], x[209], x[513], x[512], x[511]}), .y(y[284]));
  R2ind285 R2ind285_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[77], x[76], x[75], x[588], x[211], x[210], x[209], x[513], x[512], x[511]}), .y(y[285]));
  R2ind286 R2ind286_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[87], x[86], x[85], x[589], x[218], x[217], x[216], x[517], x[516], x[515]}), .y(y[286]));
  R2ind287 R2ind287_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[87], x[86], x[85], x[589], x[218], x[217], x[216], x[517], x[516], x[515]}), .y(y[287]));
  R2ind288 R2ind288_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[97], x[96], x[95], x[590], x[225], x[224], x[223], x[521], x[520], x[519]}), .y(y[288]));
  R2ind289 R2ind289_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[97], x[96], x[95], x[590], x[225], x[224], x[223], x[521], x[520], x[519]}), .y(y[289]));
  R2ind290 R2ind290_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[107], x[106], x[105], x[591], x[232], x[231], x[230], x[525], x[524], x[523]}), .y(y[290]));
  R2ind291 R2ind291_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[107], x[106], x[105], x[591], x[232], x[231], x[230], x[525], x[524], x[523]}), .y(y[291]));
  R2ind292 R2ind292_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[117], x[116], x[115], x[592], x[239], x[238], x[237], x[529], x[528], x[527]}), .y(y[292]));
  R2ind293 R2ind293_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[117], x[116], x[115], x[592], x[239], x[238], x[237], x[529], x[528], x[527]}), .y(y[293]));
  R2ind294 R2ind294_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[127], x[126], x[125], x[593], x[246], x[245], x[244], x[533], x[532], x[531]}), .y(y[294]));
  R2ind295 R2ind295_inst(.x({x[26], x[25], x[24], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[42], x[41], x[40], x[5], x[4], x[3], x[127], x[126], x[125], x[593], x[246], x[245], x[244], x[533], x[532], x[531]}), .y(y[295]));
  R2ind296 R2ind296_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[597], x[596], x[595], x[594], x[547], x[546], x[545]}), .y(y[296]));
  R2ind297 R2ind297_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[597], x[596], x[595], x[594], x[547], x[546], x[545]}), .y(y[297]));
  R2ind298 R2ind298_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[601], x[600], x[599], x[598], x[553], x[552], x[551]}), .y(y[298]));
  R2ind299 R2ind299_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[601], x[600], x[599], x[598], x[553], x[552], x[551]}), .y(y[299]));
  R2ind300 R2ind300_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[605], x[604], x[603], x[602], x[544], x[543], x[542]}), .y(y[300]));
  R2ind301 R2ind301_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[605], x[604], x[603], x[602], x[544], x[543], x[542]}), .y(y[301]));
  R2ind302 R2ind302_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[609], x[608], x[607], x[606], x[556], x[555], x[554]}), .y(y[302]));
  R2ind303 R2ind303_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[609], x[608], x[607], x[606], x[556], x[555], x[554]}), .y(y[303]));
  R2ind304 R2ind304_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[613], x[612], x[611], x[610], x[541], x[540], x[539]}), .y(y[304]));
  R2ind305 R2ind305_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[613], x[612], x[611], x[610], x[541], x[540], x[539]}), .y(y[305]));
  R2ind306 R2ind306_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[617], x[616], x[615], x[614], x[559], x[558], x[557]}), .y(y[306]));
  R2ind307 R2ind307_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[617], x[616], x[615], x[614], x[559], x[558], x[557]}), .y(y[307]));
  R2ind308 R2ind308_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[621], x[620], x[619], x[618], x[562], x[561], x[560]}), .y(y[308]));
  R2ind309 R2ind309_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[621], x[620], x[619], x[618], x[562], x[561], x[560]}), .y(y[309]));
  R2ind310 R2ind310_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[625], x[624], x[623], x[622], x[550], x[549], x[548]}), .y(y[310]));
  R2ind311 R2ind311_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[625], x[624], x[623], x[622], x[550], x[549], x[548]}), .y(y[311]));
  R2ind312 R2ind312_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[629], x[628], x[627], x[626], x[597], x[596], x[595]}), .y(y[312]));
  R2ind313 R2ind313_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[629], x[628], x[627], x[626], x[597], x[596], x[595]}), .y(y[313]));
  R2ind314 R2ind314_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[633], x[632], x[631], x[630], x[601], x[600], x[599]}), .y(y[314]));
  R2ind315 R2ind315_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[633], x[632], x[631], x[630], x[601], x[600], x[599]}), .y(y[315]));
  R2ind316 R2ind316_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[637], x[636], x[635], x[634], x[605], x[604], x[603]}), .y(y[316]));
  R2ind317 R2ind317_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[637], x[636], x[635], x[634], x[605], x[604], x[603]}), .y(y[317]));
  R2ind318 R2ind318_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[641], x[640], x[639], x[638], x[609], x[608], x[607]}), .y(y[318]));
  R2ind319 R2ind319_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[641], x[640], x[639], x[638], x[609], x[608], x[607]}), .y(y[319]));
  R2ind320 R2ind320_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[645], x[644], x[643], x[642], x[613], x[612], x[611]}), .y(y[320]));
  R2ind321 R2ind321_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[645], x[644], x[643], x[642], x[613], x[612], x[611]}), .y(y[321]));
  R2ind322 R2ind322_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[649], x[648], x[647], x[646], x[617], x[616], x[615]}), .y(y[322]));
  R2ind323 R2ind323_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[649], x[648], x[647], x[646], x[617], x[616], x[615]}), .y(y[323]));
  R2ind324 R2ind324_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[653], x[652], x[651], x[650], x[621], x[620], x[619]}), .y(y[324]));
  R2ind325 R2ind325_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[653], x[652], x[651], x[650], x[621], x[620], x[619]}), .y(y[325]));
  R2ind326 R2ind326_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[657], x[656], x[655], x[654], x[625], x[624], x[623]}), .y(y[326]));
  R2ind327 R2ind327_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[657], x[656], x[655], x[654], x[625], x[624], x[623]}), .y(y[327]));
  R2ind328 R2ind328_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[661], x[660], x[659], x[658], x[629], x[628], x[627]}), .y(y[328]));
  R2ind329 R2ind329_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[661], x[660], x[659], x[658], x[629], x[628], x[627]}), .y(y[329]));
  R2ind330 R2ind330_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[665], x[664], x[663], x[662], x[633], x[632], x[631]}), .y(y[330]));
  R2ind331 R2ind331_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[665], x[664], x[663], x[662], x[633], x[632], x[631]}), .y(y[331]));
  R2ind332 R2ind332_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[669], x[668], x[667], x[666], x[637], x[636], x[635]}), .y(y[332]));
  R2ind333 R2ind333_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[669], x[668], x[667], x[666], x[637], x[636], x[635]}), .y(y[333]));
  R2ind334 R2ind334_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[673], x[672], x[671], x[670], x[641], x[640], x[639]}), .y(y[334]));
  R2ind335 R2ind335_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[673], x[672], x[671], x[670], x[641], x[640], x[639]}), .y(y[335]));
  R2ind336 R2ind336_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[677], x[676], x[675], x[674], x[645], x[644], x[643]}), .y(y[336]));
  R2ind337 R2ind337_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[677], x[676], x[675], x[674], x[645], x[644], x[643]}), .y(y[337]));
  R2ind338 R2ind338_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[681], x[680], x[679], x[678], x[649], x[648], x[647]}), .y(y[338]));
  R2ind339 R2ind339_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[681], x[680], x[679], x[678], x[649], x[648], x[647]}), .y(y[339]));
  R2ind340 R2ind340_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[685], x[684], x[683], x[682], x[653], x[652], x[651]}), .y(y[340]));
  R2ind341 R2ind341_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[685], x[684], x[683], x[682], x[653], x[652], x[651]}), .y(y[341]));
  R2ind342 R2ind342_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[689], x[688], x[687], x[686], x[657], x[656], x[655]}), .y(y[342]));
  R2ind343 R2ind343_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[689], x[688], x[687], x[686], x[657], x[656], x[655]}), .y(y[343]));
  R2ind344 R2ind344_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[702], x[701], x[700], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[699], x[698], x[697], x[696], x[695], x[694], x[550], x[549], x[548], x[23], x[22], x[21], x[547], x[546], x[545], x[5], x[4], x[3], x[693], x[692], x[691], x[690], x[661], x[660], x[659]}), .y(y[344]));
  R2ind345 R2ind345_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[702], x[701], x[700], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[699], x[698], x[697], x[696], x[695], x[694], x[550], x[549], x[548], x[23], x[22], x[21], x[547], x[546], x[545], x[5], x[4], x[3], x[693], x[692], x[691], x[690], x[661], x[660], x[659]}), .y(y[345]));
  R2ind346 R2ind346_inst(.x({x[693], x[692], x[691], x[702], x[701], x[700], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[547], x[546], x[545], x[550], x[549], x[548], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[712], x[711], x[710], x[709], x[708], x[707], x[23], x[22], x[21], x[553], x[552], x[551], x[5], x[4], x[3], x[706], x[705], x[704], x[703], x[665], x[664], x[663]}), .y(y[346]));
  R2ind347 R2ind347_inst(.x({x[693], x[692], x[691], x[702], x[701], x[700], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[547], x[546], x[545], x[550], x[549], x[548], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[712], x[711], x[710], x[709], x[708], x[707], x[23], x[22], x[21], x[553], x[552], x[551], x[5], x[4], x[3], x[706], x[705], x[704], x[703], x[665], x[664], x[663]}), .y(y[347]));
  R2ind348 R2ind348_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[706], x[705], x[704], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[722], x[721], x[720], x[719], x[718], x[717], x[553], x[552], x[551], x[23], x[22], x[21], x[544], x[543], x[542], x[5], x[4], x[3], x[716], x[715], x[714], x[713], x[669], x[668], x[667]}), .y(y[348]));
  R2ind349 R2ind349_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[706], x[705], x[704], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[722], x[721], x[720], x[719], x[718], x[717], x[553], x[552], x[551], x[23], x[22], x[21], x[544], x[543], x[542], x[5], x[4], x[3], x[716], x[715], x[714], x[713], x[669], x[668], x[667]}), .y(y[349]));
  R2ind350 R2ind350_inst(.x({x[716], x[715], x[714], x[702], x[701], x[700], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[544], x[543], x[542], x[550], x[549], x[548], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[732], x[731], x[730], x[729], x[728], x[727], x[23], x[22], x[21], x[556], x[555], x[554], x[5], x[4], x[3], x[726], x[725], x[724], x[723], x[673], x[672], x[671]}), .y(y[350]));
  R2ind351 R2ind351_inst(.x({x[716], x[715], x[714], x[702], x[701], x[700], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[544], x[543], x[542], x[550], x[549], x[548], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[732], x[731], x[730], x[729], x[728], x[727], x[23], x[22], x[21], x[556], x[555], x[554], x[5], x[4], x[3], x[726], x[725], x[724], x[723], x[673], x[672], x[671]}), .y(y[351]));
  R2ind352 R2ind352_inst(.x({x[726], x[725], x[724], x[702], x[701], x[700], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[556], x[555], x[554], x[550], x[549], x[548], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[742], x[741], x[740], x[739], x[738], x[737], x[23], x[22], x[21], x[541], x[540], x[539], x[5], x[4], x[3], x[736], x[735], x[734], x[733], x[677], x[676], x[675]}), .y(y[352]));
  R2ind353 R2ind353_inst(.x({x[726], x[725], x[724], x[702], x[701], x[700], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[556], x[555], x[554], x[550], x[549], x[548], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[742], x[741], x[740], x[739], x[738], x[737], x[23], x[22], x[21], x[541], x[540], x[539], x[5], x[4], x[3], x[736], x[735], x[734], x[733], x[677], x[676], x[675]}), .y(y[353]));
  R2ind354 R2ind354_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[736], x[735], x[734], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[752], x[751], x[750], x[749], x[748], x[747], x[541], x[540], x[539], x[23], x[22], x[21], x[559], x[558], x[557], x[5], x[4], x[3], x[746], x[745], x[744], x[743], x[681], x[680], x[679]}), .y(y[354]));
  R2ind355 R2ind355_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[736], x[735], x[734], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[752], x[751], x[750], x[749], x[748], x[747], x[541], x[540], x[539], x[23], x[22], x[21], x[559], x[558], x[557], x[5], x[4], x[3], x[746], x[745], x[744], x[743], x[681], x[680], x[679]}), .y(y[355]));
  R2ind356 R2ind356_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[746], x[745], x[744], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[762], x[761], x[760], x[759], x[758], x[757], x[559], x[558], x[557], x[23], x[22], x[21], x[562], x[561], x[560], x[5], x[4], x[3], x[756], x[755], x[754], x[753], x[685], x[684], x[683]}), .y(y[356]));
  R2ind357 R2ind357_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[746], x[745], x[744], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[762], x[761], x[760], x[759], x[758], x[757], x[559], x[558], x[557], x[23], x[22], x[21], x[562], x[561], x[560], x[5], x[4], x[3], x[756], x[755], x[754], x[753], x[685], x[684], x[683]}), .y(y[357]));
  R2ind358 R2ind358_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[756], x[755], x[754], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[769], x[768], x[767], x[766], x[765], x[764], x[562], x[561], x[560], x[23], x[22], x[21], x[550], x[549], x[548], x[5], x[4], x[3], x[702], x[701], x[700], x[763], x[689], x[688], x[687]}), .y(y[358]));
  R2ind359 R2ind359_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[756], x[755], x[754], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[769], x[768], x[767], x[766], x[765], x[764], x[562], x[561], x[560], x[23], x[22], x[21], x[550], x[549], x[548], x[5], x[4], x[3], x[702], x[701], x[700], x[763], x[689], x[688], x[687]}), .y(y[359]));
  R2ind360 R2ind360_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[773], x[772], x[771], x[770], x[693], x[692], x[691]}), .y(y[360]));
  R2ind361 R2ind361_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[773], x[772], x[771], x[770], x[693], x[692], x[691]}), .y(y[361]));
  R2ind362 R2ind362_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[777], x[776], x[775], x[774], x[706], x[705], x[704]}), .y(y[362]));
  R2ind363 R2ind363_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[777], x[776], x[775], x[774], x[706], x[705], x[704]}), .y(y[363]));
  R2ind364 R2ind364_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[781], x[780], x[779], x[778], x[716], x[715], x[714]}), .y(y[364]));
  R2ind365 R2ind365_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[781], x[780], x[779], x[778], x[716], x[715], x[714]}), .y(y[365]));
  R2ind366 R2ind366_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[785], x[784], x[783], x[782], x[726], x[725], x[724]}), .y(y[366]));
  R2ind367 R2ind367_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[785], x[784], x[783], x[782], x[726], x[725], x[724]}), .y(y[367]));
  R2ind368 R2ind368_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[789], x[788], x[787], x[786], x[736], x[735], x[734]}), .y(y[368]));
  R2ind369 R2ind369_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[789], x[788], x[787], x[786], x[736], x[735], x[734]}), .y(y[369]));
  R2ind370 R2ind370_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[793], x[792], x[791], x[790], x[746], x[745], x[744]}), .y(y[370]));
  R2ind371 R2ind371_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[793], x[792], x[791], x[790], x[746], x[745], x[744]}), .y(y[371]));
  R2ind372 R2ind372_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[797], x[796], x[795], x[794], x[756], x[755], x[754]}), .y(y[372]));
  R2ind373 R2ind373_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[797], x[796], x[795], x[794], x[756], x[755], x[754]}), .y(y[373]));
  R2ind374 R2ind374_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[801], x[800], x[799], x[798], x[702], x[701], x[700]}), .y(y[374]));
  R2ind375 R2ind375_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[801], x[800], x[799], x[798], x[702], x[701], x[700]}), .y(y[375]));
  R2ind376 R2ind376_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[805], x[804], x[803], x[802], x[772], x[771], x[770]}), .y(y[376]));
  R2ind377 R2ind377_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[805], x[804], x[803], x[802], x[772], x[771], x[770]}), .y(y[377]));
  R2ind378 R2ind378_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[809], x[808], x[807], x[806], x[776], x[775], x[774]}), .y(y[378]));
  R2ind379 R2ind379_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[809], x[808], x[807], x[806], x[776], x[775], x[774]}), .y(y[379]));
  R2ind380 R2ind380_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[813], x[812], x[811], x[810], x[780], x[779], x[778]}), .y(y[380]));
  R2ind381 R2ind381_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[813], x[812], x[811], x[810], x[780], x[779], x[778]}), .y(y[381]));
  R2ind382 R2ind382_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[817], x[816], x[815], x[814], x[784], x[783], x[782]}), .y(y[382]));
  R2ind383 R2ind383_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[817], x[816], x[815], x[814], x[784], x[783], x[782]}), .y(y[383]));
  R2ind384 R2ind384_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[821], x[820], x[819], x[818], x[788], x[787], x[786]}), .y(y[384]));
  R2ind385 R2ind385_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[821], x[820], x[819], x[818], x[788], x[787], x[786]}), .y(y[385]));
  R2ind386 R2ind386_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[825], x[824], x[823], x[822], x[792], x[791], x[790]}), .y(y[386]));
  R2ind387 R2ind387_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[825], x[824], x[823], x[822], x[792], x[791], x[790]}), .y(y[387]));
  R2ind388 R2ind388_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[829], x[828], x[827], x[826], x[796], x[795], x[794]}), .y(y[388]));
  R2ind389 R2ind389_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[829], x[828], x[827], x[826], x[796], x[795], x[794]}), .y(y[389]));
  R2ind390 R2ind390_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[833], x[832], x[831], x[830], x[800], x[799], x[798]}), .y(y[390]));
  R2ind391 R2ind391_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[833], x[832], x[831], x[830], x[800], x[799], x[798]}), .y(y[391]));
  R2ind392 R2ind392_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[837], x[836], x[835], x[834], x[804], x[803], x[802]}), .y(y[392]));
  R2ind393 R2ind393_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[837], x[836], x[835], x[834], x[804], x[803], x[802]}), .y(y[393]));
  R2ind394 R2ind394_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[841], x[840], x[839], x[838], x[808], x[807], x[806]}), .y(y[394]));
  R2ind395 R2ind395_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[841], x[840], x[839], x[838], x[808], x[807], x[806]}), .y(y[395]));
  R2ind396 R2ind396_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[845], x[844], x[843], x[842], x[812], x[811], x[810]}), .y(y[396]));
  R2ind397 R2ind397_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[845], x[844], x[843], x[842], x[812], x[811], x[810]}), .y(y[397]));
  R2ind398 R2ind398_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[849], x[848], x[847], x[846], x[816], x[815], x[814]}), .y(y[398]));
  R2ind399 R2ind399_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[849], x[848], x[847], x[846], x[816], x[815], x[814]}), .y(y[399]));
  R2ind400 R2ind400_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[853], x[852], x[851], x[850], x[820], x[819], x[818]}), .y(y[400]));
  R2ind401 R2ind401_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[853], x[852], x[851], x[850], x[820], x[819], x[818]}), .y(y[401]));
  R2ind402 R2ind402_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[857], x[856], x[855], x[854], x[824], x[823], x[822]}), .y(y[402]));
  R2ind403 R2ind403_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[857], x[856], x[855], x[854], x[824], x[823], x[822]}), .y(y[403]));
  R2ind404 R2ind404_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[861], x[860], x[859], x[858], x[828], x[827], x[826]}), .y(y[404]));
  R2ind405 R2ind405_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[861], x[860], x[859], x[858], x[828], x[827], x[826]}), .y(y[405]));
  R2ind406 R2ind406_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[865], x[864], x[863], x[862], x[832], x[831], x[830]}), .y(y[406]));
  R2ind407 R2ind407_inst(.x({x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[5], x[4], x[3], x[865], x[864], x[863], x[862], x[832], x[831], x[830]}), .y(y[407]));
  R2ind408 R2ind408_inst(.x({x[26], x[25], x[24], x[766], x[765], x[764], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[696], x[695], x[694], x[547], x[546], x[545], x[702], x[701], x[700], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[699], x[698], x[697], x[5], x[4], x[3], x[866], x[693], x[692], x[691], x[836], x[835], x[834]}), .y(y[408]));
  R2ind409 R2ind409_inst(.x({x[26], x[25], x[24], x[766], x[765], x[764], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[696], x[695], x[694], x[547], x[546], x[545], x[702], x[701], x[700], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[699], x[698], x[697], x[5], x[4], x[3], x[866], x[693], x[692], x[691], x[836], x[835], x[834]}), .y(y[409]));
  R2ind410 R2ind410_inst(.x({x[699], x[698], x[697], x[766], x[765], x[764], x[26], x[25], x[24], x[693], x[692], x[691], x[702], x[701], x[700], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[709], x[708], x[707], x[553], x[552], x[551], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[712], x[711], x[710], x[5], x[4], x[3], x[867], x[706], x[705], x[704], x[840], x[839], x[838]}), .y(y[410]));
  R2ind411 R2ind411_inst(.x({x[699], x[698], x[697], x[766], x[765], x[764], x[26], x[25], x[24], x[693], x[692], x[691], x[702], x[701], x[700], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[709], x[708], x[707], x[553], x[552], x[551], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[712], x[711], x[710], x[5], x[4], x[3], x[867], x[706], x[705], x[704], x[840], x[839], x[838]}), .y(y[411]));
  R2ind412 R2ind412_inst(.x({x[26], x[25], x[24], x[712], x[711], x[710], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[544], x[543], x[542], x[722], x[721], x[720], x[706], x[705], x[704], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[719], x[718], x[717], x[5], x[4], x[3], x[868], x[716], x[715], x[714], x[844], x[843], x[842]}), .y(y[412]));
  R2ind413 R2ind413_inst(.x({x[26], x[25], x[24], x[712], x[711], x[710], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[544], x[543], x[542], x[722], x[721], x[720], x[706], x[705], x[704], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[719], x[718], x[717], x[5], x[4], x[3], x[868], x[716], x[715], x[714], x[844], x[843], x[842]}), .y(y[413]));
  R2ind414 R2ind414_inst(.x({x[719], x[718], x[717], x[766], x[765], x[764], x[26], x[25], x[24], x[716], x[715], x[714], x[702], x[701], x[700], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[556], x[555], x[554], x[732], x[731], x[730], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[729], x[728], x[727], x[5], x[4], x[3], x[869], x[726], x[725], x[724], x[848], x[847], x[846]}), .y(y[414]));
  R2ind415 R2ind415_inst(.x({x[719], x[718], x[717], x[766], x[765], x[764], x[26], x[25], x[24], x[716], x[715], x[714], x[702], x[701], x[700], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[556], x[555], x[554], x[732], x[731], x[730], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[729], x[728], x[727], x[5], x[4], x[3], x[869], x[726], x[725], x[724], x[848], x[847], x[846]}), .y(y[415]));
  R2ind416 R2ind416_inst(.x({x[729], x[728], x[727], x[766], x[765], x[764], x[26], x[25], x[24], x[726], x[725], x[724], x[702], x[701], x[700], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[541], x[540], x[539], x[742], x[741], x[740], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[739], x[738], x[737], x[5], x[4], x[3], x[870], x[736], x[735], x[734], x[852], x[851], x[850]}), .y(y[416]));
  R2ind417 R2ind417_inst(.x({x[729], x[728], x[727], x[766], x[765], x[764], x[26], x[25], x[24], x[726], x[725], x[724], x[702], x[701], x[700], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[541], x[540], x[539], x[742], x[741], x[740], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[739], x[738], x[737], x[5], x[4], x[3], x[870], x[736], x[735], x[734], x[852], x[851], x[850]}), .y(y[417]));
  R2ind418 R2ind418_inst(.x({x[26], x[25], x[24], x[739], x[738], x[737], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[559], x[558], x[557], x[752], x[751], x[750], x[736], x[735], x[734], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[749], x[748], x[747], x[5], x[4], x[3], x[871], x[746], x[745], x[744], x[856], x[855], x[854]}), .y(y[418]));
  R2ind419 R2ind419_inst(.x({x[26], x[25], x[24], x[739], x[738], x[737], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[559], x[558], x[557], x[752], x[751], x[750], x[736], x[735], x[734], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[749], x[748], x[747], x[5], x[4], x[3], x[871], x[746], x[745], x[744], x[856], x[855], x[854]}), .y(y[419]));
  R2ind420 R2ind420_inst(.x({x[26], x[25], x[24], x[749], x[748], x[747], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[562], x[561], x[560], x[762], x[761], x[760], x[746], x[745], x[744], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[759], x[758], x[757], x[5], x[4], x[3], x[872], x[756], x[755], x[754], x[860], x[859], x[858]}), .y(y[420]));
  R2ind421 R2ind421_inst(.x({x[26], x[25], x[24], x[749], x[748], x[747], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[562], x[561], x[560], x[762], x[761], x[760], x[746], x[745], x[744], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[759], x[758], x[757], x[5], x[4], x[3], x[872], x[756], x[755], x[754], x[860], x[859], x[858]}), .y(y[421]));
  R2ind422 R2ind422_inst(.x({x[26], x[25], x[24], x[759], x[758], x[757], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[550], x[549], x[548], x[769], x[768], x[767], x[756], x[755], x[754], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[766], x[765], x[764], x[5], x[4], x[3], x[873], x[702], x[701], x[700], x[864], x[863], x[862]}), .y(y[422]));
  R2ind423 R2ind423_inst(.x({x[26], x[25], x[24], x[759], x[758], x[757], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[550], x[549], x[548], x[769], x[768], x[767], x[756], x[755], x[754], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[23], x[22], x[21], x[766], x[765], x[764], x[5], x[4], x[3], x[873], x[702], x[701], x[700], x[864], x[863], x[862]}), .y(y[423]));
  R2ind424 R2ind424_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[880], x[879], x[878], x[877], x[876], x[875], x[874], x[699], x[698], x[697]}), .y(y[424]));
  R2ind425 R2ind425_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[880], x[879], x[878], x[877], x[876], x[875], x[874], x[699], x[698], x[697]}), .y(y[425]));
  R2ind426 R2ind426_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[887], x[886], x[885], x[884], x[883], x[882], x[881], x[712], x[711], x[710]}), .y(y[426]));
  R2ind427 R2ind427_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[887], x[886], x[885], x[884], x[883], x[882], x[881], x[712], x[711], x[710]}), .y(y[427]));
  R2ind428 R2ind428_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[894], x[893], x[892], x[891], x[890], x[889], x[888], x[719], x[718], x[717]}), .y(y[428]));
  R2ind429 R2ind429_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[894], x[893], x[892], x[891], x[890], x[889], x[888], x[719], x[718], x[717]}), .y(y[429]));
  R2ind430 R2ind430_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[901], x[900], x[899], x[898], x[897], x[896], x[895], x[729], x[728], x[727]}), .y(y[430]));
  R2ind431 R2ind431_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[901], x[900], x[899], x[898], x[897], x[896], x[895], x[729], x[728], x[727]}), .y(y[431]));
  R2ind432 R2ind432_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[908], x[907], x[906], x[905], x[904], x[903], x[902], x[739], x[738], x[737]}), .y(y[432]));
  R2ind433 R2ind433_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[908], x[907], x[906], x[905], x[904], x[903], x[902], x[739], x[738], x[737]}), .y(y[433]));
  R2ind434 R2ind434_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[915], x[914], x[913], x[912], x[911], x[910], x[909], x[749], x[748], x[747]}), .y(y[434]));
  R2ind435 R2ind435_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[915], x[914], x[913], x[912], x[911], x[910], x[909], x[749], x[748], x[747]}), .y(y[435]));
  R2ind436 R2ind436_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[922], x[921], x[920], x[919], x[918], x[917], x[916], x[759], x[758], x[757]}), .y(y[436]));
  R2ind437 R2ind437_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[922], x[921], x[920], x[919], x[918], x[917], x[916], x[759], x[758], x[757]}), .y(y[437]));
  R2ind438 R2ind438_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[929], x[928], x[927], x[926], x[925], x[924], x[923], x[766], x[765], x[764]}), .y(y[438]));
  R2ind439 R2ind439_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[929], x[928], x[927], x[926], x[925], x[924], x[923], x[766], x[765], x[764]}), .y(y[439]));
  R2ind440 R2ind440_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[876], x[875], x[874], x[933], x[932], x[931], x[930], x[880], x[879], x[878]}), .y(y[440]));
  R2ind441 R2ind441_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[876], x[875], x[874], x[933], x[932], x[931], x[930], x[880], x[879], x[878]}), .y(y[441]));
  R2ind442 R2ind442_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[883], x[882], x[881], x[937], x[936], x[935], x[934], x[887], x[886], x[885]}), .y(y[442]));
  R2ind443 R2ind443_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[883], x[882], x[881], x[937], x[936], x[935], x[934], x[887], x[886], x[885]}), .y(y[443]));
  R2ind444 R2ind444_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[890], x[889], x[888], x[941], x[940], x[939], x[938], x[894], x[893], x[892]}), .y(y[444]));
  R2ind445 R2ind445_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[890], x[889], x[888], x[941], x[940], x[939], x[938], x[894], x[893], x[892]}), .y(y[445]));
  R2ind446 R2ind446_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[897], x[896], x[895], x[945], x[944], x[943], x[942], x[901], x[900], x[899]}), .y(y[446]));
  R2ind447 R2ind447_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[897], x[896], x[895], x[945], x[944], x[943], x[942], x[901], x[900], x[899]}), .y(y[447]));
  R2ind448 R2ind448_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[904], x[903], x[902], x[949], x[948], x[947], x[946], x[908], x[907], x[906]}), .y(y[448]));
  R2ind449 R2ind449_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[904], x[903], x[902], x[949], x[948], x[947], x[946], x[908], x[907], x[906]}), .y(y[449]));
  R2ind450 R2ind450_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[911], x[910], x[909], x[953], x[952], x[951], x[950], x[915], x[914], x[913]}), .y(y[450]));
  R2ind451 R2ind451_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[911], x[910], x[909], x[953], x[952], x[951], x[950], x[915], x[914], x[913]}), .y(y[451]));
  R2ind452 R2ind452_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[918], x[917], x[916], x[957], x[956], x[955], x[954], x[922], x[921], x[920]}), .y(y[452]));
  R2ind453 R2ind453_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[918], x[917], x[916], x[957], x[956], x[955], x[954], x[922], x[921], x[920]}), .y(y[453]));
  R2ind454 R2ind454_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[925], x[924], x[923], x[961], x[960], x[959], x[958], x[929], x[928], x[927]}), .y(y[454]));
  R2ind455 R2ind455_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[925], x[924], x[923], x[961], x[960], x[959], x[958], x[929], x[928], x[927]}), .y(y[455]));
  R2ind456 R2ind456_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[932], x[931], x[930], x[962], x[699], x[698], x[697], x[876], x[875], x[874]}), .y(y[456]));
  R2ind457 R2ind457_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[932], x[931], x[930], x[962], x[699], x[698], x[697], x[876], x[875], x[874]}), .y(y[457]));
  R2ind458 R2ind458_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[936], x[935], x[934], x[963], x[712], x[711], x[710], x[883], x[882], x[881]}), .y(y[458]));
  R2ind459 R2ind459_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[936], x[935], x[934], x[963], x[712], x[711], x[710], x[883], x[882], x[881]}), .y(y[459]));
  R2ind460 R2ind460_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[940], x[939], x[938], x[964], x[719], x[718], x[717], x[890], x[889], x[888]}), .y(y[460]));
  R2ind461 R2ind461_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[940], x[939], x[938], x[964], x[719], x[718], x[717], x[890], x[889], x[888]}), .y(y[461]));
  R2ind462 R2ind462_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[944], x[943], x[942], x[965], x[729], x[728], x[727], x[897], x[896], x[895]}), .y(y[462]));
  R2ind463 R2ind463_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[944], x[943], x[942], x[965], x[729], x[728], x[727], x[897], x[896], x[895]}), .y(y[463]));
  R2ind464 R2ind464_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[948], x[947], x[946], x[966], x[739], x[738], x[737], x[904], x[903], x[902]}), .y(y[464]));
  R2ind465 R2ind465_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[948], x[947], x[946], x[966], x[739], x[738], x[737], x[904], x[903], x[902]}), .y(y[465]));
  R2ind466 R2ind466_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[952], x[951], x[950], x[967], x[749], x[748], x[747], x[911], x[910], x[909]}), .y(y[466]));
  R2ind467 R2ind467_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[952], x[951], x[950], x[967], x[749], x[748], x[747], x[911], x[910], x[909]}), .y(y[467]));
  R2ind468 R2ind468_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[956], x[955], x[954], x[968], x[759], x[758], x[757], x[918], x[917], x[916]}), .y(y[468]));
  R2ind469 R2ind469_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[956], x[955], x[954], x[968], x[759], x[758], x[757], x[918], x[917], x[916]}), .y(y[469]));
  R2ind470 R2ind470_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[960], x[959], x[958], x[969], x[766], x[765], x[764], x[925], x[924], x[923]}), .y(y[470]));
  R2ind471 R2ind471_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[960], x[959], x[958], x[969], x[766], x[765], x[764], x[925], x[924], x[923]}), .y(y[471]));
  R2ind472 R2ind472_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[769], x[768], x[767], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[547], x[546], x[545], x[693], x[692], x[691], x[766], x[765], x[764], x[23], x[22], x[21], x[699], x[698], x[697], x[5], x[4], x[3], x[696], x[695], x[694], x[970], x[880], x[879], x[878], x[932], x[931], x[930]}), .y(y[472]));
  R2ind473 R2ind473_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[769], x[768], x[767], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[547], x[546], x[545], x[693], x[692], x[691], x[766], x[765], x[764], x[23], x[22], x[21], x[699], x[698], x[697], x[5], x[4], x[3], x[696], x[695], x[694], x[970], x[880], x[879], x[878], x[932], x[931], x[930]}), .y(y[473]));
  R2ind474 R2ind474_inst(.x({x[696], x[695], x[694], x[769], x[768], x[767], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[699], x[698], x[697], x[766], x[765], x[764], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[553], x[552], x[551], x[706], x[705], x[704], x[23], x[22], x[21], x[712], x[711], x[710], x[5], x[4], x[3], x[709], x[708], x[707], x[971], x[887], x[886], x[885], x[936], x[935], x[934]}), .y(y[474]));
  R2ind475 R2ind475_inst(.x({x[696], x[695], x[694], x[769], x[768], x[767], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[699], x[698], x[697], x[766], x[765], x[764], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[553], x[552], x[551], x[706], x[705], x[704], x[23], x[22], x[21], x[712], x[711], x[710], x[5], x[4], x[3], x[709], x[708], x[707], x[971], x[887], x[886], x[885], x[936], x[935], x[934]}), .y(y[475]));
  R2ind476 R2ind476_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[709], x[708], x[707], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[716], x[715], x[714], x[544], x[543], x[542], x[712], x[711], x[710], x[23], x[22], x[21], x[719], x[718], x[717], x[5], x[4], x[3], x[722], x[721], x[720], x[972], x[894], x[893], x[892], x[940], x[939], x[938]}), .y(y[476]));
  R2ind477 R2ind477_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[709], x[708], x[707], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[716], x[715], x[714], x[544], x[543], x[542], x[712], x[711], x[710], x[23], x[22], x[21], x[719], x[718], x[717], x[5], x[4], x[3], x[722], x[721], x[720], x[972], x[894], x[893], x[892], x[940], x[939], x[938]}), .y(y[477]));
  R2ind478 R2ind478_inst(.x({x[722], x[721], x[720], x[769], x[768], x[767], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[719], x[718], x[717], x[766], x[765], x[764], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[726], x[725], x[724], x[556], x[555], x[554], x[23], x[22], x[21], x[729], x[728], x[727], x[5], x[4], x[3], x[732], x[731], x[730], x[973], x[901], x[900], x[899], x[944], x[943], x[942]}), .y(y[478]));
  R2ind479 R2ind479_inst(.x({x[722], x[721], x[720], x[769], x[768], x[767], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[719], x[718], x[717], x[766], x[765], x[764], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[726], x[725], x[724], x[556], x[555], x[554], x[23], x[22], x[21], x[729], x[728], x[727], x[5], x[4], x[3], x[732], x[731], x[730], x[973], x[901], x[900], x[899], x[944], x[943], x[942]}), .y(y[479]));
  R2ind480 R2ind480_inst(.x({x[732], x[731], x[730], x[769], x[768], x[767], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[729], x[728], x[727], x[766], x[765], x[764], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[736], x[735], x[734], x[541], x[540], x[539], x[23], x[22], x[21], x[739], x[738], x[737], x[5], x[4], x[3], x[742], x[741], x[740], x[974], x[908], x[907], x[906], x[948], x[947], x[946]}), .y(y[480]));
  R2ind481 R2ind481_inst(.x({x[732], x[731], x[730], x[769], x[768], x[767], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[729], x[728], x[727], x[766], x[765], x[764], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[736], x[735], x[734], x[541], x[540], x[539], x[23], x[22], x[21], x[739], x[738], x[737], x[5], x[4], x[3], x[742], x[741], x[740], x[974], x[908], x[907], x[906], x[948], x[947], x[946]}), .y(y[481]));
  R2ind482 R2ind482_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[742], x[741], x[740], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[746], x[745], x[744], x[559], x[558], x[557], x[739], x[738], x[737], x[23], x[22], x[21], x[749], x[748], x[747], x[5], x[4], x[3], x[752], x[751], x[750], x[975], x[915], x[914], x[913], x[952], x[951], x[950]}), .y(y[482]));
  R2ind483 R2ind483_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[742], x[741], x[740], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[746], x[745], x[744], x[559], x[558], x[557], x[739], x[738], x[737], x[23], x[22], x[21], x[749], x[748], x[747], x[5], x[4], x[3], x[752], x[751], x[750], x[975], x[915], x[914], x[913], x[952], x[951], x[950]}), .y(y[483]));
  R2ind484 R2ind484_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[752], x[751], x[750], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[756], x[755], x[754], x[562], x[561], x[560], x[749], x[748], x[747], x[23], x[22], x[21], x[759], x[758], x[757], x[5], x[4], x[3], x[762], x[761], x[760], x[976], x[922], x[921], x[920], x[956], x[955], x[954]}), .y(y[484]));
  R2ind485 R2ind485_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[752], x[751], x[750], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[756], x[755], x[754], x[562], x[561], x[560], x[749], x[748], x[747], x[23], x[22], x[21], x[759], x[758], x[757], x[5], x[4], x[3], x[762], x[761], x[760], x[976], x[922], x[921], x[920], x[956], x[955], x[954]}), .y(y[485]));
  R2ind486 R2ind486_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[762], x[761], x[760], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[702], x[701], x[700], x[550], x[549], x[548], x[759], x[758], x[757], x[23], x[22], x[21], x[766], x[765], x[764], x[5], x[4], x[3], x[769], x[768], x[767], x[977], x[929], x[928], x[927], x[960], x[959], x[958]}), .y(y[486]));
  R2ind487 R2ind487_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[762], x[761], x[760], x[42], x[41], x[40], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[702], x[701], x[700], x[550], x[549], x[548], x[759], x[758], x[757], x[23], x[22], x[21], x[766], x[765], x[764], x[5], x[4], x[3], x[769], x[768], x[767], x[977], x[929], x[928], x[927], x[960], x[959], x[958]}), .y(y[487]));
  R2ind488 R2ind488_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[984], x[983], x[982], x[981], x[980], x[979], x[978], x[696], x[695], x[694]}), .y(y[488]));
  R2ind489 R2ind489_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[984], x[983], x[982], x[981], x[980], x[979], x[978], x[696], x[695], x[694]}), .y(y[489]));
  R2ind490 R2ind490_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[991], x[990], x[989], x[988], x[987], x[986], x[985], x[709], x[708], x[707]}), .y(y[490]));
  R2ind491 R2ind491_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[991], x[990], x[989], x[988], x[987], x[986], x[985], x[709], x[708], x[707]}), .y(y[491]));
  R2ind492 R2ind492_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[998], x[997], x[996], x[995], x[994], x[993], x[992], x[722], x[721], x[720]}), .y(y[492]));
  R2ind493 R2ind493_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[998], x[997], x[996], x[995], x[994], x[993], x[992], x[722], x[721], x[720]}), .y(y[493]));
  R2ind494 R2ind494_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1005], x[1004], x[1003], x[1002], x[1001], x[1000], x[999], x[732], x[731], x[730]}), .y(y[494]));
  R2ind495 R2ind495_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1005], x[1004], x[1003], x[1002], x[1001], x[1000], x[999], x[732], x[731], x[730]}), .y(y[495]));
  R2ind496 R2ind496_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1012], x[1011], x[1010], x[1009], x[1008], x[1007], x[1006], x[742], x[741], x[740]}), .y(y[496]));
  R2ind497 R2ind497_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1012], x[1011], x[1010], x[1009], x[1008], x[1007], x[1006], x[742], x[741], x[740]}), .y(y[497]));
  R2ind498 R2ind498_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1019], x[1018], x[1017], x[1016], x[1015], x[1014], x[1013], x[752], x[751], x[750]}), .y(y[498]));
  R2ind499 R2ind499_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1019], x[1018], x[1017], x[1016], x[1015], x[1014], x[1013], x[752], x[751], x[750]}), .y(y[499]));
  R2ind500 R2ind500_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1026], x[1025], x[1024], x[1023], x[1022], x[1021], x[1020], x[762], x[761], x[760]}), .y(y[500]));
  R2ind501 R2ind501_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1026], x[1025], x[1024], x[1023], x[1022], x[1021], x[1020], x[762], x[761], x[760]}), .y(y[501]));
  R2ind502 R2ind502_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1033], x[1032], x[1031], x[1030], x[1029], x[1028], x[1027], x[769], x[768], x[767]}), .y(y[502]));
  R2ind503 R2ind503_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1033], x[1032], x[1031], x[1030], x[1029], x[1028], x[1027], x[769], x[768], x[767]}), .y(y[503]));
  R2ind504 R2ind504_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1037], x[1036], x[1035], x[1034], x[696], x[695], x[694], x[984], x[983], x[982]}), .y(y[504]));
  R2ind505 R2ind505_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1037], x[1036], x[1035], x[1034], x[696], x[695], x[694], x[984], x[983], x[982]}), .y(y[505]));
  R2ind506 R2ind506_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1041], x[1040], x[1039], x[1038], x[709], x[708], x[707], x[991], x[990], x[989]}), .y(y[506]));
  R2ind507 R2ind507_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1041], x[1040], x[1039], x[1038], x[709], x[708], x[707], x[991], x[990], x[989]}), .y(y[507]));
  R2ind508 R2ind508_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1045], x[1044], x[1043], x[1042], x[722], x[721], x[720], x[998], x[997], x[996]}), .y(y[508]));
  R2ind509 R2ind509_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1045], x[1044], x[1043], x[1042], x[722], x[721], x[720], x[998], x[997], x[996]}), .y(y[509]));
  R2ind510 R2ind510_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1049], x[1048], x[1047], x[1046], x[732], x[731], x[730], x[1005], x[1004], x[1003]}), .y(y[510]));
  R2ind511 R2ind511_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1049], x[1048], x[1047], x[1046], x[732], x[731], x[730], x[1005], x[1004], x[1003]}), .y(y[511]));
  R2ind512 R2ind512_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1053], x[1052], x[1051], x[1050], x[742], x[741], x[740], x[1012], x[1011], x[1010]}), .y(y[512]));
  R2ind513 R2ind513_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1053], x[1052], x[1051], x[1050], x[742], x[741], x[740], x[1012], x[1011], x[1010]}), .y(y[513]));
  R2ind514 R2ind514_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1057], x[1056], x[1055], x[1054], x[752], x[751], x[750], x[1019], x[1018], x[1017]}), .y(y[514]));
  R2ind515 R2ind515_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1057], x[1056], x[1055], x[1054], x[752], x[751], x[750], x[1019], x[1018], x[1017]}), .y(y[515]));
  R2ind516 R2ind516_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1061], x[1060], x[1059], x[1058], x[762], x[761], x[760], x[1026], x[1025], x[1024]}), .y(y[516]));
  R2ind517 R2ind517_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1061], x[1060], x[1059], x[1058], x[762], x[761], x[760], x[1026], x[1025], x[1024]}), .y(y[517]));
  R2ind518 R2ind518_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1065], x[1064], x[1063], x[1062], x[769], x[768], x[767], x[1033], x[1032], x[1031]}), .y(y[518]));
  R2ind519 R2ind519_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1065], x[1064], x[1063], x[1062], x[769], x[768], x[767], x[1033], x[1032], x[1031]}), .y(y[519]));
  R2ind520 R2ind520_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[980], x[979], x[978], x[1066], x[984], x[983], x[982], x[1037], x[1036], x[1035]}), .y(y[520]));
  R2ind521 R2ind521_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[980], x[979], x[978], x[1066], x[984], x[983], x[982], x[1037], x[1036], x[1035]}), .y(y[521]));
  R2ind522 R2ind522_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[987], x[986], x[985], x[1067], x[991], x[990], x[989], x[1041], x[1040], x[1039]}), .y(y[522]));
  R2ind523 R2ind523_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[987], x[986], x[985], x[1067], x[991], x[990], x[989], x[1041], x[1040], x[1039]}), .y(y[523]));
  R2ind524 R2ind524_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[994], x[993], x[992], x[1068], x[998], x[997], x[996], x[1045], x[1044], x[1043]}), .y(y[524]));
  R2ind525 R2ind525_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[994], x[993], x[992], x[1068], x[998], x[997], x[996], x[1045], x[1044], x[1043]}), .y(y[525]));
  R2ind526 R2ind526_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1001], x[1000], x[999], x[1069], x[1005], x[1004], x[1003], x[1049], x[1048], x[1047]}), .y(y[526]));
  R2ind527 R2ind527_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1001], x[1000], x[999], x[1069], x[1005], x[1004], x[1003], x[1049], x[1048], x[1047]}), .y(y[527]));
  R2ind528 R2ind528_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1008], x[1007], x[1006], x[1070], x[1012], x[1011], x[1010], x[1053], x[1052], x[1051]}), .y(y[528]));
  R2ind529 R2ind529_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1008], x[1007], x[1006], x[1070], x[1012], x[1011], x[1010], x[1053], x[1052], x[1051]}), .y(y[529]));
  R2ind530 R2ind530_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1015], x[1014], x[1013], x[1071], x[1019], x[1018], x[1017], x[1057], x[1056], x[1055]}), .y(y[530]));
  R2ind531 R2ind531_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1015], x[1014], x[1013], x[1071], x[1019], x[1018], x[1017], x[1057], x[1056], x[1055]}), .y(y[531]));
  R2ind532 R2ind532_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1022], x[1021], x[1020], x[1072], x[1026], x[1025], x[1024], x[1061], x[1060], x[1059]}), .y(y[532]));
  R2ind533 R2ind533_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1022], x[1021], x[1020], x[1072], x[1026], x[1025], x[1024], x[1061], x[1060], x[1059]}), .y(y[533]));
  R2ind534 R2ind534_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1029], x[1028], x[1027], x[1073], x[1033], x[1032], x[1031], x[1065], x[1064], x[1063]}), .y(y[534]));
  R2ind535 R2ind535_inst(.x({x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[5], x[4], x[3], x[1029], x[1028], x[1027], x[1073], x[1033], x[1032], x[1031], x[1065], x[1064], x[1063]}), .y(y[535]));
  R2ind536 R2ind536_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[273], x[272], x[271], x[107], x[106], x[105], x[559], x[558], x[557], x[87], x[86], x[85], x[556], x[555], x[554], x[67], x[66], x[65], x[553], x[552], x[551], x[127], x[126], x[125], x[269], x[268], x[267], x[261], x[260], x[259], x[253], x[252], x[251], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[550], x[549], x[548], x[42], x[41], x[40], x[20], x[19], x[18], x[693], x[692], x[691], x[699], x[698], x[697], x[769], x[768], x[767], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[57], x[56], x[55], x[547], x[546], x[545], x[696], x[695], x[694], x[5], x[4], x[3], x[1074], x[1037], x[1036], x[1035], x[980], x[979], x[978]}), .y(y[536]));
  R2ind537 R2ind537_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[273], x[272], x[271], x[107], x[106], x[105], x[559], x[558], x[557], x[87], x[86], x[85], x[556], x[555], x[554], x[67], x[66], x[65], x[553], x[552], x[551], x[127], x[126], x[125], x[269], x[268], x[267], x[261], x[260], x[259], x[253], x[252], x[251], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[550], x[549], x[548], x[42], x[41], x[40], x[20], x[19], x[18], x[693], x[692], x[691], x[699], x[698], x[697], x[769], x[768], x[767], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[57], x[56], x[55], x[547], x[546], x[545], x[696], x[695], x[694], x[5], x[4], x[3], x[1074], x[1037], x[1036], x[1035], x[980], x[979], x[978]}), .y(y[537]));
  R2ind538 R2ind538_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[261], x[260], x[259], x[253], x[252], x[251], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[127], x[126], x[125], x[107], x[106], x[105], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[257], x[256], x[255], x[265], x[264], x[263], x[277], x[276], x[275], x[269], x[268], x[267], x[273], x[272], x[271], x[57], x[56], x[55], x[249], x[248], x[247], x[547], x[546], x[545], x[550], x[549], x[548], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[696], x[695], x[694], x[769], x[768], x[767], x[42], x[41], x[40], x[20], x[19], x[18], x[706], x[705], x[704], x[712], x[711], x[710], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[67], x[66], x[65], x[553], x[552], x[551], x[709], x[708], x[707], x[5], x[4], x[3], x[1075], x[1041], x[1040], x[1039], x[987], x[986], x[985]}), .y(y[538]));
  R2ind539 R2ind539_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[261], x[260], x[259], x[253], x[252], x[251], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[127], x[126], x[125], x[107], x[106], x[105], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[257], x[256], x[255], x[265], x[264], x[263], x[277], x[276], x[275], x[269], x[268], x[267], x[273], x[272], x[271], x[57], x[56], x[55], x[249], x[248], x[247], x[547], x[546], x[545], x[550], x[549], x[548], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[696], x[695], x[694], x[769], x[768], x[767], x[42], x[41], x[40], x[20], x[19], x[18], x[706], x[705], x[704], x[712], x[711], x[710], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[67], x[66], x[65], x[553], x[552], x[551], x[709], x[708], x[707], x[5], x[4], x[3], x[1075], x[1041], x[1040], x[1039], x[987], x[986], x[985]}), .y(y[539]));
  R2ind540 R2ind540_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[117], x[116], x[115], x[562], x[561], x[560], x[67], x[66], x[65], x[107], x[106], x[105], x[559], x[558], x[557], x[127], x[126], x[125], x[550], x[549], x[548], x[261], x[260], x[259], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[253], x[252], x[251], x[269], x[268], x[267], x[277], x[276], x[275], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[553], x[552], x[551], x[42], x[41], x[40], x[20], x[19], x[18], x[719], x[718], x[717], x[716], x[715], x[714], x[709], x[708], x[707], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[77], x[76], x[75], x[544], x[543], x[542], x[722], x[721], x[720], x[5], x[4], x[3], x[1076], x[1045], x[1044], x[1043], x[994], x[993], x[992]}), .y(y[540]));
  R2ind541 R2ind541_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[117], x[116], x[115], x[562], x[561], x[560], x[67], x[66], x[65], x[107], x[106], x[105], x[559], x[558], x[557], x[127], x[126], x[125], x[550], x[549], x[548], x[261], x[260], x[259], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[253], x[252], x[251], x[269], x[268], x[267], x[277], x[276], x[275], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[257], x[256], x[255], x[265], x[264], x[263], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[553], x[552], x[551], x[42], x[41], x[40], x[20], x[19], x[18], x[719], x[718], x[717], x[716], x[715], x[714], x[709], x[708], x[707], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[77], x[76], x[75], x[544], x[543], x[542], x[722], x[721], x[720], x[5], x[4], x[3], x[1076], x[1045], x[1044], x[1043], x[994], x[993], x[992]}), .y(y[541]));
  R2ind542 R2ind542_inst(.x({x[67], x[66], x[65], x[553], x[552], x[551], x[261], x[260], x[259], x[107], x[106], x[105], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[253], x[252], x[251], x[269], x[268], x[267], x[273], x[272], x[271], x[77], x[76], x[75], x[97], x[96], x[95], x[541], x[540], x[539], x[127], x[126], x[125], x[57], x[56], x[55], x[547], x[546], x[545], x[257], x[256], x[255], x[265], x[264], x[263], x[277], x[276], x[275], x[249], x[248], x[247], x[544], x[543], x[542], x[550], x[549], x[548], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[722], x[721], x[720], x[769], x[768], x[767], x[42], x[41], x[40], x[20], x[19], x[18], x[729], x[728], x[727], x[726], x[725], x[724], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[87], x[86], x[85], x[556], x[555], x[554], x[732], x[731], x[730], x[5], x[4], x[3], x[1077], x[1049], x[1048], x[1047], x[1001], x[1000], x[999]}), .y(y[542]));
  R2ind543 R2ind543_inst(.x({x[67], x[66], x[65], x[553], x[552], x[551], x[261], x[260], x[259], x[107], x[106], x[105], x[559], x[558], x[557], x[117], x[116], x[115], x[562], x[561], x[560], x[253], x[252], x[251], x[269], x[268], x[267], x[273], x[272], x[271], x[77], x[76], x[75], x[97], x[96], x[95], x[541], x[540], x[539], x[127], x[126], x[125], x[57], x[56], x[55], x[547], x[546], x[545], x[257], x[256], x[255], x[265], x[264], x[263], x[277], x[276], x[275], x[249], x[248], x[247], x[544], x[543], x[542], x[550], x[549], x[548], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[722], x[721], x[720], x[769], x[768], x[767], x[42], x[41], x[40], x[20], x[19], x[18], x[729], x[728], x[727], x[726], x[725], x[724], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[87], x[86], x[85], x[556], x[555], x[554], x[732], x[731], x[730], x[5], x[4], x[3], x[1077], x[1049], x[1048], x[1047], x[1001], x[1000], x[999]}), .y(y[543]));
  R2ind544 R2ind544_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[107], x[106], x[105], x[559], x[558], x[557], x[67], x[66], x[65], x[553], x[552], x[551], x[87], x[86], x[85], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[127], x[126], x[125], x[269], x[268], x[267], x[253], x[252], x[251], x[261], x[260], x[259], x[249], x[248], x[247], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[257], x[256], x[255], x[265], x[264], x[263], x[556], x[555], x[554], x[550], x[549], x[548], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[732], x[731], x[730], x[769], x[768], x[767], x[42], x[41], x[40], x[20], x[19], x[18], x[739], x[738], x[737], x[736], x[735], x[734], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[97], x[96], x[95], x[541], x[540], x[539], x[742], x[741], x[740], x[5], x[4], x[3], x[1078], x[1053], x[1052], x[1051], x[1008], x[1007], x[1006]}), .y(y[544]));
  R2ind545 R2ind545_inst(.x({x[117], x[116], x[115], x[562], x[561], x[560], x[107], x[106], x[105], x[559], x[558], x[557], x[67], x[66], x[65], x[553], x[552], x[551], x[87], x[86], x[85], x[273], x[272], x[271], x[57], x[56], x[55], x[547], x[546], x[545], x[127], x[126], x[125], x[269], x[268], x[267], x[253], x[252], x[251], x[261], x[260], x[259], x[249], x[248], x[247], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[257], x[256], x[255], x[265], x[264], x[263], x[556], x[555], x[554], x[550], x[549], x[548], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[732], x[731], x[730], x[769], x[768], x[767], x[42], x[41], x[40], x[20], x[19], x[18], x[739], x[738], x[737], x[736], x[735], x[734], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[97], x[96], x[95], x[541], x[540], x[539], x[742], x[741], x[740], x[5], x[4], x[3], x[1078], x[1053], x[1052], x[1051], x[1008], x[1007], x[1006]}), .y(y[545]));
  R2ind546 R2ind546_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[117], x[116], x[115], x[562], x[561], x[560], x[97], x[96], x[95], x[261], x[260], x[259], x[57], x[56], x[55], x[547], x[546], x[545], x[67], x[66], x[65], x[553], x[552], x[551], x[269], x[268], x[267], x[273], x[272], x[271], x[265], x[264], x[263], x[249], x[248], x[247], x[253], x[252], x[251], x[77], x[76], x[75], x[544], x[543], x[542], x[127], x[126], x[125], x[550], x[549], x[548], x[257], x[256], x[255], x[277], x[276], x[275], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[541], x[540], x[539], x[42], x[41], x[40], x[20], x[19], x[18], x[749], x[748], x[747], x[746], x[745], x[744], x[742], x[741], x[740], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[107], x[106], x[105], x[559], x[558], x[557], x[752], x[751], x[750], x[5], x[4], x[3], x[1079], x[1057], x[1056], x[1055], x[1015], x[1014], x[1013]}), .y(y[546]));
  R2ind547 R2ind547_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[117], x[116], x[115], x[562], x[561], x[560], x[97], x[96], x[95], x[261], x[260], x[259], x[57], x[56], x[55], x[547], x[546], x[545], x[67], x[66], x[65], x[553], x[552], x[551], x[269], x[268], x[267], x[273], x[272], x[271], x[265], x[264], x[263], x[249], x[248], x[247], x[253], x[252], x[251], x[77], x[76], x[75], x[544], x[543], x[542], x[127], x[126], x[125], x[550], x[549], x[548], x[257], x[256], x[255], x[277], x[276], x[275], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[541], x[540], x[539], x[42], x[41], x[40], x[20], x[19], x[18], x[749], x[748], x[747], x[746], x[745], x[744], x[742], x[741], x[740], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[107], x[106], x[105], x[559], x[558], x[557], x[752], x[751], x[750], x[5], x[4], x[3], x[1079], x[1057], x[1056], x[1055], x[1015], x[1014], x[1013]}), .y(y[547]));
  R2ind548 R2ind548_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[57], x[56], x[55], x[547], x[546], x[545], x[67], x[66], x[65], x[553], x[552], x[551], x[107], x[106], x[105], x[261], x[260], x[259], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[253], x[252], x[251], x[269], x[268], x[267], x[273], x[272], x[271], x[77], x[76], x[75], x[544], x[543], x[542], x[127], x[126], x[125], x[550], x[549], x[548], x[265], x[264], x[263], x[257], x[256], x[255], x[277], x[276], x[275], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[559], x[558], x[557], x[42], x[41], x[40], x[20], x[19], x[18], x[759], x[758], x[757], x[756], x[755], x[754], x[752], x[751], x[750], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[117], x[116], x[115], x[562], x[561], x[560], x[762], x[761], x[760], x[5], x[4], x[3], x[1080], x[1061], x[1060], x[1059], x[1022], x[1021], x[1020]}), .y(y[548]));
  R2ind549 R2ind549_inst(.x({x[87], x[86], x[85], x[556], x[555], x[554], x[57], x[56], x[55], x[547], x[546], x[545], x[67], x[66], x[65], x[553], x[552], x[551], x[107], x[106], x[105], x[261], x[260], x[259], x[97], x[96], x[95], x[541], x[540], x[539], x[249], x[248], x[247], x[253], x[252], x[251], x[269], x[268], x[267], x[273], x[272], x[271], x[77], x[76], x[75], x[544], x[543], x[542], x[127], x[126], x[125], x[550], x[549], x[548], x[265], x[264], x[263], x[257], x[256], x[255], x[277], x[276], x[275], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[559], x[558], x[557], x[42], x[41], x[40], x[20], x[19], x[18], x[759], x[758], x[757], x[756], x[755], x[754], x[752], x[751], x[750], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[117], x[116], x[115], x[562], x[561], x[560], x[762], x[761], x[760], x[5], x[4], x[3], x[1080], x[1061], x[1060], x[1059], x[1022], x[1021], x[1020]}), .y(y[549]));
  R2ind550 R2ind550_inst(.x({x[117], x[116], x[115], x[57], x[56], x[55], x[547], x[546], x[545], x[107], x[106], x[105], x[559], x[558], x[557], x[67], x[66], x[65], x[553], x[552], x[551], x[87], x[86], x[85], x[556], x[555], x[554], x[273], x[272], x[271], x[249], x[248], x[247], x[269], x[268], x[267], x[253], x[252], x[251], x[261], x[260], x[259], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[257], x[256], x[255], x[265], x[264], x[263], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[562], x[561], x[560], x[42], x[41], x[40], x[20], x[19], x[18], x[766], x[765], x[764], x[702], x[701], x[700], x[762], x[761], x[760], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[127], x[126], x[125], x[550], x[549], x[548], x[769], x[768], x[767], x[5], x[4], x[3], x[1081], x[1065], x[1064], x[1063], x[1029], x[1028], x[1027]}), .y(y[550]));
  R2ind551 R2ind551_inst(.x({x[117], x[116], x[115], x[57], x[56], x[55], x[547], x[546], x[545], x[107], x[106], x[105], x[559], x[558], x[557], x[67], x[66], x[65], x[553], x[552], x[551], x[87], x[86], x[85], x[556], x[555], x[554], x[273], x[272], x[271], x[249], x[248], x[247], x[269], x[268], x[267], x[253], x[252], x[251], x[261], x[260], x[259], x[277], x[276], x[275], x[77], x[76], x[75], x[544], x[543], x[542], x[97], x[96], x[95], x[541], x[540], x[539], x[257], x[256], x[255], x[265], x[264], x[263], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[562], x[561], x[560], x[42], x[41], x[40], x[20], x[19], x[18], x[766], x[765], x[764], x[702], x[701], x[700], x[762], x[761], x[760], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[23], x[22], x[21], x[127], x[126], x[125], x[550], x[549], x[548], x[769], x[768], x[767], x[5], x[4], x[3], x[1081], x[1065], x[1064], x[1063], x[1029], x[1028], x[1027]}), .y(y[551]));
endmodule

