/* modified netlist. Source: module sbox in file Designs/AESSbox//Canright/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 8 time(s)  */

module sbox_HPC2_ClockGating_d2 (X_s0, clk, X_s1, X_s2, Fresh, rst, Y_s0, Y_s1, Y_s2, Synch);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input rst ;
    input [119:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    output Synch ;
    wire sbe_n10 ;
    wire sbe_n9 ;
    wire sbe_n8 ;
    wire sbe_n7 ;
    wire sbe_n6 ;
    wire sbe_n5 ;
    wire sbe_n4 ;
    wire sbe_n3 ;
    wire sbe_n12 ;
    wire sbe_n11 ;
    wire sbe_n2 ;
    wire sbe_n1 ;
    wire sbe_n25 ;
    wire sbe_n24 ;
    wire sbe_n23 ;
    wire sbe_n22 ;
    wire sbe_n21 ;
    wire sbe_n20 ;
    wire sbe_n19 ;
    wire sbe_n18 ;
    wire sbe_n17 ;
    wire sbe_n16 ;
    wire sbe_n15 ;
    wire sbe_n14 ;
    wire sbe_D_0_ ;
    wire sbe_D_2_ ;
    wire sbe_D_3_ ;
    wire sbe_D_5_ ;
    wire sbe_D_6_ ;
    wire sbe_C_0_ ;
    wire sbe_C_1_ ;
    wire sbe_C_2_ ;
    wire sbe_C_3_ ;
    wire sbe_C_4_ ;
    wire sbe_C_5_ ;
    wire sbe_C_6_ ;
    wire sbe_C_7_ ;
    wire sbe_Y_0_ ;
    wire sbe_Y_1_ ;
    wire sbe_Y_2_ ;
    wire sbe_Y_4_ ;
    wire sbe_Y_5_ ;
    wire sbe_Y_6_ ;
    wire sbe_B_3_ ;
    wire sbe_B_6_ ;
    wire sbe_sel_in_m7_n8 ;
    wire sbe_sel_in_m6_n8 ;
    wire sbe_sel_in_m5_n8 ;
    wire sbe_sel_in_m4_n8 ;
    wire sbe_sel_in_m3_n8 ;
    wire sbe_sel_in_m2_n8 ;
    wire sbe_sel_in_m1_n8 ;
    wire sbe_sel_in_m0_n8 ;
    wire sbe_inv_n21 ;
    wire sbe_inv_n20 ;
    wire sbe_inv_n19 ;
    wire sbe_inv_n18 ;
    wire sbe_inv_n17 ;
    wire sbe_inv_n16 ;
    wire sbe_inv_n15 ;
    wire sbe_inv_n14 ;
    wire sbe_inv_n13 ;
    wire sbe_inv_n12 ;
    wire sbe_inv_n11 ;
    wire sbe_inv_n10 ;
    wire sbe_inv_n9 ;
    wire sbe_inv_n8 ;
    wire sbe_inv_n7 ;
    wire sbe_inv_n6 ;
    wire sbe_inv_n5 ;
    wire sbe_inv_n4 ;
    wire sbe_inv_n3 ;
    wire sbe_inv_n2 ;
    wire sbe_inv_dd ;
    wire sbe_inv_dh ;
    wire sbe_inv_dl ;
    wire sbe_inv_sd_0_ ;
    wire sbe_inv_sd_1_ ;
    wire sbe_inv_d_0_ ;
    wire sbe_inv_d_1_ ;
    wire sbe_inv_d_2_ ;
    wire sbe_inv_d_3_ ;
    wire sbe_inv_bb ;
    wire sbe_inv_bh ;
    wire sbe_inv_bl ;
    wire sbe_inv_aa ;
    wire sbe_inv_ah ;
    wire sbe_inv_al ;
    wire sbe_inv_sb_0_ ;
    wire sbe_inv_sb_1_ ;
    wire sbe_inv_sa_0_ ;
    wire sbe_inv_sa_1_ ;
    wire sbe_inv_dinv_n4 ;
    wire sbe_inv_dinv_n3 ;
    wire sbe_inv_dinv_n2 ;
    wire sbe_inv_dinv_n1 ;
    wire sbe_inv_dinv_sd ;
    wire sbe_inv_dinv_d_0_ ;
    wire sbe_inv_dinv_d_1_ ;
    wire sbe_inv_dinv_sb ;
    wire sbe_inv_dinv_sa ;
    wire sbe_inv_dinv_pmul_n9 ;
    wire sbe_inv_dinv_pmul_n8 ;
    wire sbe_inv_dinv_pmul_n7 ;
    wire sbe_inv_dinv_qmul_n9 ;
    wire sbe_inv_dinv_qmul_n8 ;
    wire sbe_inv_dinv_qmul_n7 ;
    wire sbe_inv_pmul_p_0_ ;
    wire sbe_inv_pmul_p_1_ ;
    wire sbe_inv_pmul_himul_n9 ;
    wire sbe_inv_pmul_himul_n8 ;
    wire sbe_inv_pmul_himul_n7 ;
    wire sbe_inv_pmul_lomul_n9 ;
    wire sbe_inv_pmul_lomul_n8 ;
    wire sbe_inv_pmul_lomul_n7 ;
    wire sbe_inv_pmul_summul_n9 ;
    wire sbe_inv_pmul_summul_n8 ;
    wire sbe_inv_pmul_summul_n7 ;
    wire sbe_inv_qmul_p_0_ ;
    wire sbe_inv_qmul_p_1_ ;
    wire sbe_inv_qmul_himul_n9 ;
    wire sbe_inv_qmul_himul_n8 ;
    wire sbe_inv_qmul_himul_n7 ;
    wire sbe_inv_qmul_lomul_n9 ;
    wire sbe_inv_qmul_lomul_n8 ;
    wire sbe_inv_qmul_lomul_n7 ;
    wire sbe_inv_qmul_summul_n9 ;
    wire sbe_inv_qmul_summul_n8 ;
    wire sbe_inv_qmul_summul_n7 ;
    wire sbe_sel_out_m7_n8 ;
    wire sbe_sel_out_m6_n8 ;
    wire sbe_sel_out_m5_n8 ;
    wire sbe_sel_out_m4_n8 ;
    wire sbe_sel_out_m3_n8 ;
    wire sbe_sel_out_m2_n8 ;
    wire sbe_sel_out_m1_n8 ;
    wire sbe_sel_out_m0_n8 ;
    wire [7:0] O ;
    wire [6:3] sbe_X ;
    wire [7:0] sbe_Z ;
    wire [3:0] sbe_inv_c ;
    wire [1:0] sbe_inv_pmul_pl ;
    wire [1:0] sbe_inv_pmul_ph ;
    wire [1:0] sbe_inv_qmul_pl ;
    wire [1:0] sbe_inv_qmul_ph ;
    wire new_AGEMA_signal_196 ;
    wire new_AGEMA_signal_197 ;
    wire new_AGEMA_signal_202 ;
    wire new_AGEMA_signal_203 ;
    wire new_AGEMA_signal_204 ;
    wire new_AGEMA_signal_205 ;
    wire new_AGEMA_signal_208 ;
    wire new_AGEMA_signal_209 ;
    wire new_AGEMA_signal_210 ;
    wire new_AGEMA_signal_211 ;
    wire new_AGEMA_signal_214 ;
    wire new_AGEMA_signal_215 ;
    wire new_AGEMA_signal_216 ;
    wire new_AGEMA_signal_217 ;
    wire new_AGEMA_signal_220 ;
    wire new_AGEMA_signal_221 ;
    wire new_AGEMA_signal_222 ;
    wire new_AGEMA_signal_223 ;
    wire new_AGEMA_signal_226 ;
    wire new_AGEMA_signal_227 ;
    wire new_AGEMA_signal_228 ;
    wire new_AGEMA_signal_229 ;
    wire new_AGEMA_signal_230 ;
    wire new_AGEMA_signal_231 ;
    wire new_AGEMA_signal_232 ;
    wire new_AGEMA_signal_233 ;
    wire new_AGEMA_signal_234 ;
    wire new_AGEMA_signal_235 ;
    wire new_AGEMA_signal_236 ;
    wire new_AGEMA_signal_237 ;
    wire new_AGEMA_signal_238 ;
    wire new_AGEMA_signal_239 ;
    wire new_AGEMA_signal_240 ;
    wire new_AGEMA_signal_241 ;
    wire new_AGEMA_signal_242 ;
    wire new_AGEMA_signal_243 ;
    wire new_AGEMA_signal_244 ;
    wire new_AGEMA_signal_245 ;
    wire new_AGEMA_signal_246 ;
    wire new_AGEMA_signal_247 ;
    wire new_AGEMA_signal_248 ;
    wire new_AGEMA_signal_249 ;
    wire new_AGEMA_signal_250 ;
    wire new_AGEMA_signal_251 ;
    wire new_AGEMA_signal_252 ;
    wire new_AGEMA_signal_253 ;
    wire new_AGEMA_signal_254 ;
    wire new_AGEMA_signal_255 ;
    wire new_AGEMA_signal_256 ;
    wire new_AGEMA_signal_257 ;
    wire new_AGEMA_signal_258 ;
    wire new_AGEMA_signal_259 ;
    wire new_AGEMA_signal_260 ;
    wire new_AGEMA_signal_261 ;
    wire new_AGEMA_signal_262 ;
    wire new_AGEMA_signal_263 ;
    wire new_AGEMA_signal_264 ;
    wire new_AGEMA_signal_265 ;
    wire new_AGEMA_signal_266 ;
    wire new_AGEMA_signal_267 ;
    wire new_AGEMA_signal_268 ;
    wire new_AGEMA_signal_269 ;
    wire new_AGEMA_signal_270 ;
    wire new_AGEMA_signal_271 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;
    wire new_AGEMA_signal_482 ;
    wire new_AGEMA_signal_483 ;
    wire new_AGEMA_signal_484 ;
    wire new_AGEMA_signal_485 ;
    wire new_AGEMA_signal_486 ;
    wire new_AGEMA_signal_487 ;
    wire new_AGEMA_signal_488 ;
    wire new_AGEMA_signal_489 ;
    wire new_AGEMA_signal_490 ;
    wire new_AGEMA_signal_491 ;
    wire new_AGEMA_signal_492 ;
    wire new_AGEMA_signal_493 ;
    wire new_AGEMA_signal_494 ;
    wire new_AGEMA_signal_495 ;
    wire new_AGEMA_signal_496 ;
    wire new_AGEMA_signal_497 ;
    wire new_AGEMA_signal_498 ;
    wire new_AGEMA_signal_499 ;
    wire new_AGEMA_signal_500 ;
    wire new_AGEMA_signal_501 ;
    wire new_AGEMA_signal_502 ;
    wire new_AGEMA_signal_503 ;
    wire new_AGEMA_signal_504 ;
    wire new_AGEMA_signal_505 ;
    wire new_AGEMA_signal_506 ;
    wire new_AGEMA_signal_507 ;
    wire new_AGEMA_signal_508 ;
    wire new_AGEMA_signal_509 ;
    wire new_AGEMA_signal_510 ;
    wire new_AGEMA_signal_511 ;
    wire new_AGEMA_signal_512 ;
    wire new_AGEMA_signal_513 ;
    wire new_AGEMA_signal_514 ;
    wire new_AGEMA_signal_515 ;
    wire new_AGEMA_signal_516 ;
    wire new_AGEMA_signal_517 ;
    wire new_AGEMA_signal_518 ;
    wire new_AGEMA_signal_519 ;
    wire new_AGEMA_signal_520 ;
    wire new_AGEMA_signal_521 ;
    wire new_AGEMA_signal_522 ;
    wire new_AGEMA_signal_523 ;
    wire new_AGEMA_signal_524 ;
    wire new_AGEMA_signal_525 ;
    wire new_AGEMA_signal_526 ;
    wire new_AGEMA_signal_527 ;
    wire new_AGEMA_signal_528 ;
    wire new_AGEMA_signal_529 ;
    wire new_AGEMA_signal_530 ;
    wire new_AGEMA_signal_531 ;
    wire new_AGEMA_signal_532 ;
    wire new_AGEMA_signal_533 ;
    wire new_AGEMA_signal_534 ;
    wire new_AGEMA_signal_535 ;
    wire new_AGEMA_signal_536 ;
    wire new_AGEMA_signal_537 ;
    wire new_AGEMA_signal_538 ;
    wire new_AGEMA_signal_539 ;
    wire new_AGEMA_signal_540 ;
    wire new_AGEMA_signal_541 ;
    wire new_AGEMA_signal_542 ;
    wire new_AGEMA_signal_543 ;
    wire clk_gated ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U39 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_231, new_AGEMA_signal_230, sbe_n25}), .c ({new_AGEMA_signal_237, new_AGEMA_signal_236, sbe_n12}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U38 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_243, new_AGEMA_signal_242, sbe_Y_4_}), .c ({new_AGEMA_signal_253, new_AGEMA_signal_252, sbe_n24}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U37 ( .a ({new_AGEMA_signal_215, new_AGEMA_signal_214, sbe_Y_2_}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, sbe_n10}), .c ({new_AGEMA_signal_239, new_AGEMA_signal_238, sbe_n23}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U36 ( .a ({new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n9}), .b ({new_AGEMA_signal_203, new_AGEMA_signal_202, sbe_n8}), .c ({new_AGEMA_signal_223, new_AGEMA_signal_222, sbe_n22}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U35 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_205, new_AGEMA_signal_204, sbe_n11}), .c ({new_AGEMA_signal_211, new_AGEMA_signal_210, sbe_n21}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U29 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, sbe_n10}), .c ({new_AGEMA_signal_241, new_AGEMA_signal_240, sbe_Y_6_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U28 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[4], X_s1[4], X_s0[4]}), .c ({new_AGEMA_signal_197, new_AGEMA_signal_196, sbe_Y_5_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U27 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_227, new_AGEMA_signal_226, sbe_n10}), .c ({new_AGEMA_signal_243, new_AGEMA_signal_242, sbe_Y_4_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U26 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n9}), .c ({new_AGEMA_signal_227, new_AGEMA_signal_226, sbe_n10}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U25 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({new_AGEMA_signal_203, new_AGEMA_signal_202, sbe_n8}), .c ({new_AGEMA_signal_215, new_AGEMA_signal_214, sbe_Y_2_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U24 ( .a ({X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s2[7], X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_203, new_AGEMA_signal_202, sbe_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U23 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_221, new_AGEMA_signal_220, sbe_n7}), .c ({new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_Y_1_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U22 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_245, new_AGEMA_signal_244, sbe_B_6_}), .c ({new_AGEMA_signal_255, new_AGEMA_signal_254, sbe_Y_0_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U8 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({new_AGEMA_signal_231, new_AGEMA_signal_230, sbe_n25}), .c ({new_AGEMA_signal_245, new_AGEMA_signal_244, sbe_B_6_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U7 ( .a ({X_s2[5], X_s1[5], X_s0[5]}), .b ({new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n9}), .c ({new_AGEMA_signal_231, new_AGEMA_signal_230, sbe_n25}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U6 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({new_AGEMA_signal_209, new_AGEMA_signal_208, sbe_n2}), .c ({new_AGEMA_signal_217, new_AGEMA_signal_216, sbe_n9}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U5 ( .a ({new_AGEMA_signal_233, new_AGEMA_signal_232, sbe_n3}), .b ({new_AGEMA_signal_205, new_AGEMA_signal_204, sbe_n11}), .c ({new_AGEMA_signal_247, new_AGEMA_signal_246, sbe_B_3_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U4 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({new_AGEMA_signal_221, new_AGEMA_signal_220, sbe_n7}), .c ({new_AGEMA_signal_233, new_AGEMA_signal_232, sbe_n3}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U3 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({new_AGEMA_signal_209, new_AGEMA_signal_208, sbe_n2}), .c ({new_AGEMA_signal_221, new_AGEMA_signal_220, sbe_n7}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U2 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s2[7], X_s1[7], X_s0[7]}), .c ({new_AGEMA_signal_205, new_AGEMA_signal_204, sbe_n11}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_U1 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({new_AGEMA_signal_209, new_AGEMA_signal_208, sbe_n2}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m7_U2 ( .a ({new_AGEMA_signal_257, new_AGEMA_signal_256, sbe_sel_in_m7_n8}), .b ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_205, new_AGEMA_signal_204, sbe_n11}), .a ({new_AGEMA_signal_239, new_AGEMA_signal_238, sbe_n23}), .c ({new_AGEMA_signal_257, new_AGEMA_signal_256, sbe_sel_in_m7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m6_U2 ( .a ({new_AGEMA_signal_259, new_AGEMA_signal_258, sbe_sel_in_m6_n8}), .b ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_241, new_AGEMA_signal_240, sbe_Y_6_}), .a ({new_AGEMA_signal_245, new_AGEMA_signal_244, sbe_B_6_}), .c ({new_AGEMA_signal_259, new_AGEMA_signal_258, sbe_sel_in_m6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m5_U2 ( .a ({new_AGEMA_signal_261, new_AGEMA_signal_260, sbe_sel_in_m5_n8}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_197, new_AGEMA_signal_196, sbe_Y_5_}), .a ({new_AGEMA_signal_237, new_AGEMA_signal_236, sbe_n12}), .c ({new_AGEMA_signal_261, new_AGEMA_signal_260, sbe_sel_in_m5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m4_U2 ( .a ({new_AGEMA_signal_263, new_AGEMA_signal_262, sbe_sel_in_m4_n8}), .b ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_243, new_AGEMA_signal_242, sbe_Y_4_}), .a ({new_AGEMA_signal_223, new_AGEMA_signal_222, sbe_n22}), .c ({new_AGEMA_signal_263, new_AGEMA_signal_262, sbe_sel_in_m4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m3_U2 ( .a ({new_AGEMA_signal_265, new_AGEMA_signal_264, sbe_sel_in_m3_n8}), .b ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_211, new_AGEMA_signal_210, sbe_n21}), .a ({new_AGEMA_signal_247, new_AGEMA_signal_246, sbe_B_3_}), .c ({new_AGEMA_signal_265, new_AGEMA_signal_264, sbe_sel_in_m3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m2_U2 ( .a ({new_AGEMA_signal_235, new_AGEMA_signal_234, sbe_sel_in_m2_n8}), .b ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_215, new_AGEMA_signal_214, sbe_Y_2_}), .a ({new_AGEMA_signal_209, new_AGEMA_signal_208, sbe_n2}), .c ({new_AGEMA_signal_235, new_AGEMA_signal_234, sbe_sel_in_m2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m1_U2 ( .a ({new_AGEMA_signal_251, new_AGEMA_signal_250, sbe_sel_in_m1_n8}), .b ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_229, new_AGEMA_signal_228, sbe_Y_1_}), .a ({new_AGEMA_signal_231, new_AGEMA_signal_230, sbe_n25}), .c ({new_AGEMA_signal_251, new_AGEMA_signal_250, sbe_sel_in_m1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m0_U2 ( .a ({new_AGEMA_signal_279, new_AGEMA_signal_278, sbe_sel_in_m0_n8}), .b ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_in_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_255, new_AGEMA_signal_254, sbe_Y_0_}), .a ({new_AGEMA_signal_253, new_AGEMA_signal_252, sbe_n24}), .c ({new_AGEMA_signal_279, new_AGEMA_signal_278, sbe_sel_in_m0_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U10 ( .a ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}), .b ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}), .c ({new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_inv_bl}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U9 ( .a ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}), .b ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}), .c ({new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_inv_bh}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U8 ( .a ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}), .c ({new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_inv_bb}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U7 ( .a ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}), .b ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}), .c ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U6 ( .a ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}), .b ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}), .c ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U5 ( .a ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}), .c ({new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_inv_al}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U4 ( .a ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}), .b ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}), .c ({new_AGEMA_signal_295, new_AGEMA_signal_294, sbe_inv_ah}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U3 ( .a ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}), .c ({new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_inv_aa}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U2 ( .a ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}), .b ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}), .c ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U1 ( .a ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}), .c ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}) ) ;
    ClockGatingController #(9) ClockGatingInst ( .clk ( clk ), .rst ( rst ), .GatedClk ( clk_gated ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U34 ( .a ({new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_inv_n21}), .b ({new_AGEMA_signal_327, new_AGEMA_signal_326, sbe_inv_n20}), .c ({new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_inv_c[3]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U33 ( .a ({new_AGEMA_signal_315, new_AGEMA_signal_314, sbe_inv_n19}), .b ({new_AGEMA_signal_283, new_AGEMA_signal_282, sbe_inv_n18}), .c ({new_AGEMA_signal_327, new_AGEMA_signal_326, sbe_inv_n20}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U32 ( .a ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}), .b ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}), .clk ( clk ), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_283, new_AGEMA_signal_282, sbe_inv_n18}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U31 ( .a ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}), .clk ( clk ), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({new_AGEMA_signal_315, new_AGEMA_signal_314, sbe_inv_n19}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U30 ( .a ({new_AGEMA_signal_333, new_AGEMA_signal_332, sbe_inv_n17}), .b ({new_AGEMA_signal_303, new_AGEMA_signal_302, sbe_inv_n16}), .c ({new_AGEMA_signal_337, new_AGEMA_signal_336, sbe_inv_n21}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U29 ( .a ({new_AGEMA_signal_329, new_AGEMA_signal_328, sbe_inv_n15}), .b ({new_AGEMA_signal_317, new_AGEMA_signal_316, sbe_inv_n14}), .c ({new_AGEMA_signal_339, new_AGEMA_signal_338, sbe_inv_c[2]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U28 ( .a ({new_AGEMA_signal_301, new_AGEMA_signal_300, sbe_inv_n13}), .b ({new_AGEMA_signal_285, new_AGEMA_signal_284, sbe_inv_n12}), .c ({new_AGEMA_signal_317, new_AGEMA_signal_316, sbe_inv_n14}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U27 ( .a ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}), .b ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}), .clk ( clk ), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_285, new_AGEMA_signal_284, sbe_inv_n12}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U26 ( .a ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}), .clk ( clk ), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({new_AGEMA_signal_301, new_AGEMA_signal_300, sbe_inv_n13}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U25 ( .a ({new_AGEMA_signal_323, new_AGEMA_signal_322, sbe_inv_n11}), .b ({new_AGEMA_signal_303, new_AGEMA_signal_302, sbe_inv_n16}), .c ({new_AGEMA_signal_329, new_AGEMA_signal_328, sbe_inv_n15}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U24 ( .a ({new_AGEMA_signal_295, new_AGEMA_signal_294, sbe_inv_ah}), .b ({new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_inv_bh}), .clk ( clk ), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({new_AGEMA_signal_303, new_AGEMA_signal_302, sbe_inv_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U23 ( .a ({new_AGEMA_signal_341, new_AGEMA_signal_340, sbe_inv_n10}), .b ({new_AGEMA_signal_331, new_AGEMA_signal_330, sbe_inv_n9}), .c ({new_AGEMA_signal_347, new_AGEMA_signal_346, sbe_inv_c[1]}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U22 ( .a ({new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_inv_n8}), .b ({new_AGEMA_signal_287, new_AGEMA_signal_286, sbe_inv_n7}), .c ({new_AGEMA_signal_331, new_AGEMA_signal_330, sbe_inv_n9}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U21 ( .a ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}), .clk ( clk ), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({new_AGEMA_signal_287, new_AGEMA_signal_286, sbe_inv_n7}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U20 ( .a ({new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_inv_al}), .b ({new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_inv_bl}), .clk ( clk ), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({new_AGEMA_signal_319, new_AGEMA_signal_318, sbe_inv_n8}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U19 ( .a ({new_AGEMA_signal_333, new_AGEMA_signal_332, sbe_inv_n17}), .b ({new_AGEMA_signal_323, new_AGEMA_signal_322, sbe_inv_n11}), .c ({new_AGEMA_signal_341, new_AGEMA_signal_340, sbe_inv_n10}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U18 ( .a ({new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_inv_aa}), .b ({new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_inv_bb}), .clk ( clk ), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({new_AGEMA_signal_333, new_AGEMA_signal_332, sbe_inv_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U17 ( .a ({new_AGEMA_signal_323, new_AGEMA_signal_322, sbe_inv_n11}), .b ({new_AGEMA_signal_343, new_AGEMA_signal_342, sbe_inv_n6}), .c ({new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_c[0]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U16 ( .a ({new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_inv_n5}), .b ({new_AGEMA_signal_335, new_AGEMA_signal_334, sbe_inv_n4}), .c ({new_AGEMA_signal_343, new_AGEMA_signal_342, sbe_inv_n6}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U15 ( .a ({new_AGEMA_signal_305, new_AGEMA_signal_304, sbe_inv_n3}), .b ({new_AGEMA_signal_321, new_AGEMA_signal_320, sbe_inv_n2}), .c ({new_AGEMA_signal_335, new_AGEMA_signal_334, sbe_inv_n4}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U14 ( .a ({new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_inv_al}), .b ({new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_inv_bl}), .clk ( clk ), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({new_AGEMA_signal_321, new_AGEMA_signal_320, sbe_inv_n2}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U13 ( .a ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}), .b ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({new_AGEMA_signal_305, new_AGEMA_signal_304, sbe_inv_n3}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U12 ( .a ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}), .b ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}), .clk ( clk ), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_307, new_AGEMA_signal_306, sbe_inv_n5}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U11 ( .a ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}), .b ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}), .clk ( clk ), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({new_AGEMA_signal_323, new_AGEMA_signal_322, sbe_inv_n11}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U2 ( .a ({new_AGEMA_signal_339, new_AGEMA_signal_338, sbe_inv_c[2]}), .b ({new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_inv_c[3]}), .c ({new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_dinv_sa}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U1 ( .a ({new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_c[0]}), .b ({new_AGEMA_signal_347, new_AGEMA_signal_346, sbe_inv_c[1]}), .c ({new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_inv_dinv_sb}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U9 ( .a ({new_AGEMA_signal_363, new_AGEMA_signal_362, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_inv_dinv_d_1_}), .c ({new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_dinv_sd}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U8 ( .a ({new_AGEMA_signal_351, new_AGEMA_signal_350, sbe_inv_dinv_n4}), .b ({new_AGEMA_signal_359, new_AGEMA_signal_358, sbe_inv_dinv_n3}), .c ({new_AGEMA_signal_363, new_AGEMA_signal_362, sbe_inv_dinv_d_0_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U7 ( .a ({new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_inv_dinv_sb}), .b ({new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_dinv_sa}), .clk ( clk ), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({new_AGEMA_signal_359, new_AGEMA_signal_358, sbe_inv_dinv_n3}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U6 ( .a ({new_AGEMA_signal_347, new_AGEMA_signal_346, sbe_inv_c[1]}), .b ({new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_inv_c[3]}), .clk ( clk ), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({new_AGEMA_signal_351, new_AGEMA_signal_350, sbe_inv_dinv_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U5 ( .a ({new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_inv_dinv_n2}), .b ({new_AGEMA_signal_353, new_AGEMA_signal_352, sbe_inv_dinv_n1}), .c ({new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_inv_dinv_d_1_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U4 ( .a ({new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_c[0]}), .b ({new_AGEMA_signal_339, new_AGEMA_signal_338, sbe_inv_c[2]}), .clk ( clk ), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({new_AGEMA_signal_353, new_AGEMA_signal_352, sbe_inv_dinv_n1}) ) ;
    nor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_U3 ( .a ({new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_inv_dinv_sb}), .b ({new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_dinv_sa}), .clk ( clk ), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({new_AGEMA_signal_361, new_AGEMA_signal_360, sbe_inv_dinv_n2}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U39 ( .a ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}), .b ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}), .c ({new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_dl}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U38 ( .a ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}), .b ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}), .c ({new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_dh}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U37 ( .a ({new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_395, new_AGEMA_signal_394, sbe_inv_sd_1_}), .c ({new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_dd}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U36 ( .a ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}), .b ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}), .c ({new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_sd_0_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_U35 ( .a ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}), .b ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}), .c ({new_AGEMA_signal_395, new_AGEMA_signal_394, sbe_inv_sd_1_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_pmul_U5 ( .a ({new_AGEMA_signal_377, new_AGEMA_signal_376, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_369, new_AGEMA_signal_368, sbe_inv_dinv_pmul_n8}), .c ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_pmul_U4 ( .a ({new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_inv_dinv_d_1_}), .b ({new_AGEMA_signal_347, new_AGEMA_signal_346, sbe_inv_c[1]}), .clk ( clk ), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({new_AGEMA_signal_369, new_AGEMA_signal_368, sbe_inv_dinv_pmul_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_pmul_U3 ( .a ({new_AGEMA_signal_377, new_AGEMA_signal_376, sbe_inv_dinv_pmul_n9}), .b ({new_AGEMA_signal_371, new_AGEMA_signal_370, sbe_inv_dinv_pmul_n7}), .c ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_pmul_U2 ( .a ({new_AGEMA_signal_363, new_AGEMA_signal_362, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_349, new_AGEMA_signal_348, sbe_inv_c[0]}), .clk ( clk ), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({new_AGEMA_signal_371, new_AGEMA_signal_370, sbe_inv_dinv_pmul_n7}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_pmul_U1 ( .a ({new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_dinv_sd}), .b ({new_AGEMA_signal_357, new_AGEMA_signal_356, sbe_inv_dinv_sb}), .clk ( clk ), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({new_AGEMA_signal_377, new_AGEMA_signal_376, sbe_inv_dinv_pmul_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_qmul_U5 ( .a ({new_AGEMA_signal_379, new_AGEMA_signal_378, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_dinv_qmul_n8}), .c ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_qmul_U4 ( .a ({new_AGEMA_signal_365, new_AGEMA_signal_364, sbe_inv_dinv_d_1_}), .b ({new_AGEMA_signal_345, new_AGEMA_signal_344, sbe_inv_c[3]}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({new_AGEMA_signal_373, new_AGEMA_signal_372, sbe_inv_dinv_qmul_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_qmul_U3 ( .a ({new_AGEMA_signal_379, new_AGEMA_signal_378, sbe_inv_dinv_qmul_n9}), .b ({new_AGEMA_signal_375, new_AGEMA_signal_374, sbe_inv_dinv_qmul_n7}), .c ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_qmul_U2 ( .a ({new_AGEMA_signal_363, new_AGEMA_signal_362, sbe_inv_dinv_d_0_}), .b ({new_AGEMA_signal_339, new_AGEMA_signal_338, sbe_inv_c[2]}), .clk ( clk ), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_375, new_AGEMA_signal_374, sbe_inv_dinv_qmul_n7}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_dinv_qmul_U1 ( .a ({new_AGEMA_signal_367, new_AGEMA_signal_366, sbe_inv_dinv_sd}), .b ({new_AGEMA_signal_355, new_AGEMA_signal_354, sbe_inv_dinv_sa}), .clk ( clk ), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({new_AGEMA_signal_379, new_AGEMA_signal_378, sbe_inv_dinv_qmul_n9}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    not_masked #(.security_order(2), .pipeline(0)) sbe_U40 ( .a ({new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_C_2_}), .b ({new_AGEMA_signal_467, new_AGEMA_signal_466, sbe_n1}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U34 ( .a ({new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_C_7_}), .b ({new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_n17}), .c ({new_AGEMA_signal_503, new_AGEMA_signal_502, sbe_n16}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U33 ( .a ({new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_C_4_}), .b ({new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_n18}), .c ({new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_n17}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U32 ( .a ({new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_C_5_}), .b ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .c ({new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_n18}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U31 ( .a ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .b ({new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_C_4_}), .c ({new_AGEMA_signal_483, new_AGEMA_signal_482, sbe_n15}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U30 ( .a ({new_AGEMA_signal_455, new_AGEMA_signal_454, sbe_C_6_}), .b ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .c ({new_AGEMA_signal_485, new_AGEMA_signal_484, sbe_n14}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U21 ( .a ({new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_n6}), .b ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .c ({new_AGEMA_signal_521, new_AGEMA_signal_520, sbe_X[6]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U20 ( .a ({new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_C_2_}), .b ({new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_n6}), .c ({new_AGEMA_signal_523, new_AGEMA_signal_522, sbe_X[5]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U19 ( .a ({new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_D_5_}), .b ({new_AGEMA_signal_495, new_AGEMA_signal_494, sbe_n20}), .c ({new_AGEMA_signal_505, new_AGEMA_signal_504, sbe_n6}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U18 ( .a ({new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_n5}), .b ({new_AGEMA_signal_491, new_AGEMA_signal_490, sbe_D_0_}), .c ({new_AGEMA_signal_507, new_AGEMA_signal_506, sbe_X[3]}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U17 ( .a ({new_AGEMA_signal_495, new_AGEMA_signal_494, sbe_n20}), .b ({new_AGEMA_signal_471, new_AGEMA_signal_470, sbe_n4}), .c ({new_AGEMA_signal_509, new_AGEMA_signal_508, sbe_D_3_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U16 ( .a ({new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_C_5_}), .b ({new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_D_6_}), .c ({new_AGEMA_signal_495, new_AGEMA_signal_494, sbe_n20}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U15 ( .a ({new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_C_7_}), .b ({new_AGEMA_signal_477, new_AGEMA_signal_476, sbe_C_3_}), .c ({new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_D_6_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U14 ( .a ({new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_D_5_}), .b ({new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_n5}), .c ({new_AGEMA_signal_511, new_AGEMA_signal_510, sbe_D_2_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U13 ( .a ({new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_C_2_}), .b ({new_AGEMA_signal_489, new_AGEMA_signal_488, sbe_n19}), .c ({new_AGEMA_signal_497, new_AGEMA_signal_496, sbe_n5}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U12 ( .a ({new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_C_5_}), .b ({new_AGEMA_signal_477, new_AGEMA_signal_476, sbe_C_3_}), .c ({new_AGEMA_signal_489, new_AGEMA_signal_488, sbe_n19}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U11 ( .a ({new_AGEMA_signal_455, new_AGEMA_signal_454, sbe_C_6_}), .b ({new_AGEMA_signal_463, new_AGEMA_signal_462, sbe_C_0_}), .c ({new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_D_5_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U10 ( .a ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}), .b ({new_AGEMA_signal_471, new_AGEMA_signal_470, sbe_n4}), .c ({new_AGEMA_signal_491, new_AGEMA_signal_490, sbe_D_0_}) ) ;
    xnor_HPC2 #(.security_order(2), .pipeline(0)) sbe_U9 ( .a ({new_AGEMA_signal_455, new_AGEMA_signal_454, sbe_C_6_}), .b ({new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_C_4_}), .c ({new_AGEMA_signal_471, new_AGEMA_signal_470, sbe_n4}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_U4 ( .a ({new_AGEMA_signal_459, new_AGEMA_signal_458, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_431, new_AGEMA_signal_430, sbe_inv_pmul_ph[1]}), .c ({new_AGEMA_signal_473, new_AGEMA_signal_472, sbe_C_7_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_U3 ( .a ({new_AGEMA_signal_441, new_AGEMA_signal_440, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_433, new_AGEMA_signal_432, sbe_inv_pmul_ph[0]}), .c ({new_AGEMA_signal_455, new_AGEMA_signal_454, sbe_C_6_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_U2 ( .a ({new_AGEMA_signal_459, new_AGEMA_signal_458, sbe_inv_pmul_p_1_}), .b ({new_AGEMA_signal_435, new_AGEMA_signal_434, sbe_inv_pmul_pl[1]}), .c ({new_AGEMA_signal_475, new_AGEMA_signal_474, sbe_C_5_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_U1 ( .a ({new_AGEMA_signal_441, new_AGEMA_signal_440, sbe_inv_pmul_p_0_}), .b ({new_AGEMA_signal_437, new_AGEMA_signal_436, sbe_inv_pmul_pl[0]}), .c ({new_AGEMA_signal_457, new_AGEMA_signal_456, sbe_C_4_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_himul_U5 ( .a ({new_AGEMA_signal_415, new_AGEMA_signal_414, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_397, new_AGEMA_signal_396, sbe_inv_pmul_himul_n8}), .c ({new_AGEMA_signal_431, new_AGEMA_signal_430, sbe_inv_pmul_ph[1]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_himul_U4 ( .a ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}), .b ({new_AGEMA_signal_277, new_AGEMA_signal_276, sbe_Z[3]}), .clk ( clk ), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({new_AGEMA_signal_397, new_AGEMA_signal_396, sbe_inv_pmul_himul_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_himul_U3 ( .a ({new_AGEMA_signal_415, new_AGEMA_signal_414, sbe_inv_pmul_himul_n9}), .b ({new_AGEMA_signal_399, new_AGEMA_signal_398, sbe_inv_pmul_himul_n7}), .c ({new_AGEMA_signal_433, new_AGEMA_signal_432, sbe_inv_pmul_ph[0]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_himul_U2 ( .a ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}), .b ({new_AGEMA_signal_249, new_AGEMA_signal_248, sbe_Z[2]}), .clk ( clk ), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({new_AGEMA_signal_399, new_AGEMA_signal_398, sbe_inv_pmul_himul_n7}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_himul_U1 ( .a ({new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_dh}), .b ({new_AGEMA_signal_289, new_AGEMA_signal_288, sbe_inv_bh}), .clk ( clk ), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({new_AGEMA_signal_415, new_AGEMA_signal_414, sbe_inv_pmul_himul_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_lomul_U5 ( .a ({new_AGEMA_signal_417, new_AGEMA_signal_416, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_401, new_AGEMA_signal_400, sbe_inv_pmul_lomul_n8}), .c ({new_AGEMA_signal_435, new_AGEMA_signal_434, sbe_inv_pmul_pl[1]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_lomul_U4 ( .a ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}), .b ({new_AGEMA_signal_267, new_AGEMA_signal_266, sbe_Z[1]}), .clk ( clk ), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({new_AGEMA_signal_401, new_AGEMA_signal_400, sbe_inv_pmul_lomul_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_lomul_U3 ( .a ({new_AGEMA_signal_417, new_AGEMA_signal_416, sbe_inv_pmul_lomul_n9}), .b ({new_AGEMA_signal_403, new_AGEMA_signal_402, sbe_inv_pmul_lomul_n7}), .c ({new_AGEMA_signal_437, new_AGEMA_signal_436, sbe_inv_pmul_pl[0]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_lomul_U2 ( .a ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}), .b ({new_AGEMA_signal_281, new_AGEMA_signal_280, sbe_Z[0]}), .clk ( clk ), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({new_AGEMA_signal_403, new_AGEMA_signal_402, sbe_inv_pmul_lomul_n7}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_lomul_U1 ( .a ({new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_dl}), .b ({new_AGEMA_signal_309, new_AGEMA_signal_308, sbe_inv_bl}), .clk ( clk ), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({new_AGEMA_signal_417, new_AGEMA_signal_416, sbe_inv_pmul_lomul_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_summul_U5 ( .a ({new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_439, new_AGEMA_signal_438, sbe_inv_pmul_summul_n8}), .c ({new_AGEMA_signal_459, new_AGEMA_signal_458, sbe_inv_pmul_p_1_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_summul_U4 ( .a ({new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_dd}), .b ({new_AGEMA_signal_325, new_AGEMA_signal_324, sbe_inv_bb}), .clk ( clk ), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({new_AGEMA_signal_439, new_AGEMA_signal_438, sbe_inv_pmul_summul_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_summul_U3 ( .a ({new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_pmul_summul_n9}), .b ({new_AGEMA_signal_419, new_AGEMA_signal_418, sbe_inv_pmul_summul_n7}), .c ({new_AGEMA_signal_441, new_AGEMA_signal_440, sbe_inv_pmul_p_0_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_summul_U2 ( .a ({new_AGEMA_signal_395, new_AGEMA_signal_394, sbe_inv_sd_1_}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_290, sbe_inv_sb_1_}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({new_AGEMA_signal_419, new_AGEMA_signal_418, sbe_inv_pmul_summul_n7}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_pmul_summul_U1 ( .a ({new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_311, new_AGEMA_signal_310, sbe_inv_sb_0_}), .clk ( clk ), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_421, new_AGEMA_signal_420, sbe_inv_pmul_summul_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_U4 ( .a ({new_AGEMA_signal_465, new_AGEMA_signal_464, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_443, new_AGEMA_signal_442, sbe_inv_qmul_ph[1]}), .c ({new_AGEMA_signal_477, new_AGEMA_signal_476, sbe_C_3_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_U3 ( .a ({new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_445, new_AGEMA_signal_444, sbe_inv_qmul_ph[0]}), .c ({new_AGEMA_signal_461, new_AGEMA_signal_460, sbe_C_2_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_U2 ( .a ({new_AGEMA_signal_465, new_AGEMA_signal_464, sbe_inv_qmul_p_1_}), .b ({new_AGEMA_signal_447, new_AGEMA_signal_446, sbe_inv_qmul_pl[1]}), .c ({new_AGEMA_signal_479, new_AGEMA_signal_478, sbe_C_1_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_U1 ( .a ({new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_qmul_p_0_}), .b ({new_AGEMA_signal_449, new_AGEMA_signal_448, sbe_inv_qmul_pl[0]}), .c ({new_AGEMA_signal_463, new_AGEMA_signal_462, sbe_C_0_}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_himul_U5 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_405, new_AGEMA_signal_404, sbe_inv_qmul_himul_n8}), .c ({new_AGEMA_signal_443, new_AGEMA_signal_442, sbe_inv_qmul_ph[1]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_himul_U4 ( .a ({new_AGEMA_signal_381, new_AGEMA_signal_380, sbe_inv_d_3_}), .b ({new_AGEMA_signal_269, new_AGEMA_signal_268, sbe_Z[7]}), .clk ( clk ), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({new_AGEMA_signal_405, new_AGEMA_signal_404, sbe_inv_qmul_himul_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_himul_U3 ( .a ({new_AGEMA_signal_423, new_AGEMA_signal_422, sbe_inv_qmul_himul_n9}), .b ({new_AGEMA_signal_407, new_AGEMA_signal_406, sbe_inv_qmul_himul_n7}), .c ({new_AGEMA_signal_445, new_AGEMA_signal_444, sbe_inv_qmul_ph[0]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_himul_U2 ( .a ({new_AGEMA_signal_383, new_AGEMA_signal_382, sbe_inv_d_2_}), .b ({new_AGEMA_signal_271, new_AGEMA_signal_270, sbe_Z[6]}), .clk ( clk ), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({new_AGEMA_signal_407, new_AGEMA_signal_406, sbe_inv_qmul_himul_n7}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_himul_U1 ( .a ({new_AGEMA_signal_391, new_AGEMA_signal_390, sbe_inv_dh}), .b ({new_AGEMA_signal_295, new_AGEMA_signal_294, sbe_inv_ah}), .clk ( clk ), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({new_AGEMA_signal_423, new_AGEMA_signal_422, sbe_inv_qmul_himul_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_lomul_U5 ( .a ({new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_409, new_AGEMA_signal_408, sbe_inv_qmul_lomul_n8}), .c ({new_AGEMA_signal_447, new_AGEMA_signal_446, sbe_inv_qmul_pl[1]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_lomul_U4 ( .a ({new_AGEMA_signal_385, new_AGEMA_signal_384, sbe_inv_d_1_}), .b ({new_AGEMA_signal_273, new_AGEMA_signal_272, sbe_Z[5]}), .clk ( clk ), .r ({Fresh[104], Fresh[103], Fresh[102]}), .c ({new_AGEMA_signal_409, new_AGEMA_signal_408, sbe_inv_qmul_lomul_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_lomul_U3 ( .a ({new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_qmul_lomul_n9}), .b ({new_AGEMA_signal_411, new_AGEMA_signal_410, sbe_inv_qmul_lomul_n7}), .c ({new_AGEMA_signal_449, new_AGEMA_signal_448, sbe_inv_qmul_pl[0]}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_lomul_U2 ( .a ({new_AGEMA_signal_387, new_AGEMA_signal_386, sbe_inv_d_0_}), .b ({new_AGEMA_signal_275, new_AGEMA_signal_274, sbe_Z[4]}), .clk ( clk ), .r ({Fresh[107], Fresh[106], Fresh[105]}), .c ({new_AGEMA_signal_411, new_AGEMA_signal_410, sbe_inv_qmul_lomul_n7}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_lomul_U1 ( .a ({new_AGEMA_signal_389, new_AGEMA_signal_388, sbe_inv_dl}), .b ({new_AGEMA_signal_293, new_AGEMA_signal_292, sbe_inv_al}), .clk ( clk ), .r ({Fresh[110], Fresh[109], Fresh[108]}), .c ({new_AGEMA_signal_425, new_AGEMA_signal_424, sbe_inv_qmul_lomul_n9}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_summul_U5 ( .a ({new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_451, new_AGEMA_signal_450, sbe_inv_qmul_summul_n8}), .c ({new_AGEMA_signal_465, new_AGEMA_signal_464, sbe_inv_qmul_p_1_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_summul_U4 ( .a ({new_AGEMA_signal_413, new_AGEMA_signal_412, sbe_inv_dd}), .b ({new_AGEMA_signal_313, new_AGEMA_signal_312, sbe_inv_aa}), .clk ( clk ), .r ({Fresh[113], Fresh[112], Fresh[111]}), .c ({new_AGEMA_signal_451, new_AGEMA_signal_450, sbe_inv_qmul_summul_n8}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_summul_U3 ( .a ({new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_qmul_summul_n9}), .b ({new_AGEMA_signal_427, new_AGEMA_signal_426, sbe_inv_qmul_summul_n7}), .c ({new_AGEMA_signal_453, new_AGEMA_signal_452, sbe_inv_qmul_p_0_}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_summul_U2 ( .a ({new_AGEMA_signal_395, new_AGEMA_signal_394, sbe_inv_sd_1_}), .b ({new_AGEMA_signal_299, new_AGEMA_signal_298, sbe_inv_sa_1_}), .clk ( clk ), .r ({Fresh[116], Fresh[115], Fresh[114]}), .c ({new_AGEMA_signal_427, new_AGEMA_signal_426, sbe_inv_qmul_summul_n7}) ) ;
    nand_HPC2 #(.security_order(2), .pipeline(0)) sbe_inv_qmul_summul_U1 ( .a ({new_AGEMA_signal_393, new_AGEMA_signal_392, sbe_inv_sd_0_}), .b ({new_AGEMA_signal_297, new_AGEMA_signal_296, sbe_inv_sa_0_}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117]}), .c ({new_AGEMA_signal_429, new_AGEMA_signal_428, sbe_inv_qmul_summul_n9}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m7_U2 ( .a ({new_AGEMA_signal_499, new_AGEMA_signal_498, sbe_sel_out_m7_n8}), .b ({new_AGEMA_signal_513, new_AGEMA_signal_512, O[7]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m7_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_483, new_AGEMA_signal_482, sbe_n15}), .a ({new_AGEMA_signal_489, new_AGEMA_signal_488, sbe_n19}), .c ({new_AGEMA_signal_499, new_AGEMA_signal_498, sbe_sel_out_m7_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m6_U2 ( .a ({new_AGEMA_signal_533, new_AGEMA_signal_532, sbe_sel_out_m6_n8}), .b ({new_AGEMA_signal_541, new_AGEMA_signal_540, O[6]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m6_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_521, new_AGEMA_signal_520, sbe_X[6]}), .a ({new_AGEMA_signal_487, new_AGEMA_signal_486, sbe_D_6_}), .c ({new_AGEMA_signal_533, new_AGEMA_signal_532, sbe_sel_out_m6_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m5_U2 ( .a ({new_AGEMA_signal_535, new_AGEMA_signal_534, sbe_sel_out_m5_n8}), .b ({new_AGEMA_signal_543, new_AGEMA_signal_542, O[5]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m5_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_523, new_AGEMA_signal_522, sbe_X[5]}), .a ({new_AGEMA_signal_469, new_AGEMA_signal_468, sbe_D_5_}), .c ({new_AGEMA_signal_535, new_AGEMA_signal_534, sbe_sel_out_m5_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m4_U2 ( .a ({new_AGEMA_signal_515, new_AGEMA_signal_514, sbe_sel_out_m4_n8}), .b ({new_AGEMA_signal_525, new_AGEMA_signal_524, O[4]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m4_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_485, new_AGEMA_signal_484, sbe_n14}), .a ({new_AGEMA_signal_495, new_AGEMA_signal_494, sbe_n20}), .c ({new_AGEMA_signal_515, new_AGEMA_signal_514, sbe_sel_out_m4_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m3_U2 ( .a ({new_AGEMA_signal_527, new_AGEMA_signal_526, sbe_sel_out_m3_n8}), .b ({new_AGEMA_signal_537, new_AGEMA_signal_536, O[3]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m3_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_507, new_AGEMA_signal_506, sbe_X[3]}), .a ({new_AGEMA_signal_509, new_AGEMA_signal_508, sbe_D_3_}), .c ({new_AGEMA_signal_527, new_AGEMA_signal_526, sbe_sel_out_m3_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m2_U2 ( .a ({new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_sel_out_m2_n8}), .b ({new_AGEMA_signal_539, new_AGEMA_signal_538, O[2]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m2_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_503, new_AGEMA_signal_502, sbe_n16}), .a ({new_AGEMA_signal_511, new_AGEMA_signal_510, sbe_D_2_}), .c ({new_AGEMA_signal_529, new_AGEMA_signal_528, sbe_sel_out_m2_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m1_U2 ( .a ({new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_sel_out_m1_n8}), .b ({new_AGEMA_signal_531, new_AGEMA_signal_530, O[1]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m1_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_481, new_AGEMA_signal_480, sbe_n18}), .a ({new_AGEMA_signal_493, new_AGEMA_signal_492, sbe_n17}), .c ({new_AGEMA_signal_517, new_AGEMA_signal_516, sbe_sel_out_m1_n8}) ) ;
    not_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m0_U2 ( .a ({new_AGEMA_signal_501, new_AGEMA_signal_500, sbe_sel_out_m0_n8}), .b ({new_AGEMA_signal_519, new_AGEMA_signal_518, O[0]}) ) ;
    mux2_masked #(.security_order(2), .pipeline(0)) sbe_sel_out_m0_U1 ( .s ( 1'b1 ), .b ({new_AGEMA_signal_467, new_AGEMA_signal_466, sbe_n1}), .a ({new_AGEMA_signal_491, new_AGEMA_signal_490, sbe_D_0_}), .c ({new_AGEMA_signal_501, new_AGEMA_signal_500, sbe_sel_out_m0_n8}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(0)) Y_reg_7_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_513, new_AGEMA_signal_512, O[7]}), .Q ({Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Y_reg_6_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_541, new_AGEMA_signal_540, O[6]}), .Q ({Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Y_reg_5_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_543, new_AGEMA_signal_542, O[5]}), .Q ({Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Y_reg_4_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_525, new_AGEMA_signal_524, O[4]}), .Q ({Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Y_reg_3_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_537, new_AGEMA_signal_536, O[3]}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Y_reg_2_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_539, new_AGEMA_signal_538, O[2]}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Y_reg_1_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_531, new_AGEMA_signal_530, O[1]}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(0)) Y_reg_0_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_519, new_AGEMA_signal_518, O[0]}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
