/* modified netlist. Source: module sbox in file ../sbox_lookup/sbox.v */
/* 10 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 11 register stage(s) in total */

module sbox_HPC2_Pipeline_d4 (SI_s0, clk, SI_s1, SI_s2, SI_s3, SI_s4, Fresh, SO_s0, SO_s1, SO_s2, SO_s3, SO_s4);
    input [3:0] SI_s0 ;
    input clk ;
    input [3:0] SI_s1 ;
    input [3:0] SI_s2 ;
    input [3:0] SI_s3 ;
    input [3:0] SI_s4 ;
    input [129:0] Fresh ;
    output [3:0] SO_s0 ;
    output [3:0] SO_s1 ;
    output [3:0] SO_s2 ;
    output [3:0] SO_s3 ;
    output [3:0] SO_s4 ;
    wire N9 ;
    wire N12 ;
    wire N19 ;
    wire N27 ;
    wire n40 ;
    wire n41 ;
    wire n42 ;
    wire n43 ;
    wire n44 ;
    wire n45 ;
    wire n46 ;
    wire n47 ;
    wire n48 ;
    wire n49 ;
    wire n50 ;
    wire n51 ;
    wire n52 ;
    wire n53 ;
    wire n54 ;
    wire new_AGEMA_signal_38 ;
    wire new_AGEMA_signal_39 ;
    wire new_AGEMA_signal_40 ;
    wire new_AGEMA_signal_41 ;
    wire new_AGEMA_signal_50 ;
    wire new_AGEMA_signal_51 ;
    wire new_AGEMA_signal_52 ;
    wire new_AGEMA_signal_53 ;
    wire new_AGEMA_signal_58 ;
    wire new_AGEMA_signal_59 ;
    wire new_AGEMA_signal_60 ;
    wire new_AGEMA_signal_61 ;
    wire new_AGEMA_signal_62 ;
    wire new_AGEMA_signal_63 ;
    wire new_AGEMA_signal_64 ;
    wire new_AGEMA_signal_65 ;
    wire new_AGEMA_signal_66 ;
    wire new_AGEMA_signal_67 ;
    wire new_AGEMA_signal_68 ;
    wire new_AGEMA_signal_69 ;
    wire new_AGEMA_signal_70 ;
    wire new_AGEMA_signal_71 ;
    wire new_AGEMA_signal_72 ;
    wire new_AGEMA_signal_73 ;
    wire new_AGEMA_signal_74 ;
    wire new_AGEMA_signal_75 ;
    wire new_AGEMA_signal_76 ;
    wire new_AGEMA_signal_77 ;
    wire new_AGEMA_signal_78 ;
    wire new_AGEMA_signal_79 ;
    wire new_AGEMA_signal_80 ;
    wire new_AGEMA_signal_81 ;
    wire new_AGEMA_signal_82 ;
    wire new_AGEMA_signal_83 ;
    wire new_AGEMA_signal_84 ;
    wire new_AGEMA_signal_85 ;
    wire new_AGEMA_signal_86 ;
    wire new_AGEMA_signal_87 ;
    wire new_AGEMA_signal_88 ;
    wire new_AGEMA_signal_89 ;
    wire new_AGEMA_signal_90 ;
    wire new_AGEMA_signal_91 ;
    wire new_AGEMA_signal_92 ;
    wire new_AGEMA_signal_93 ;
    wire new_AGEMA_signal_94 ;
    wire new_AGEMA_signal_95 ;
    wire new_AGEMA_signal_96 ;
    wire new_AGEMA_signal_97 ;
    wire new_AGEMA_signal_98 ;
    wire new_AGEMA_signal_99 ;
    wire new_AGEMA_signal_100 ;
    wire new_AGEMA_signal_101 ;
    wire new_AGEMA_signal_102 ;
    wire new_AGEMA_signal_103 ;
    wire new_AGEMA_signal_104 ;
    wire new_AGEMA_signal_105 ;
    wire new_AGEMA_signal_106 ;
    wire new_AGEMA_signal_107 ;
    wire new_AGEMA_signal_108 ;
    wire new_AGEMA_signal_109 ;
    wire new_AGEMA_signal_110 ;
    wire new_AGEMA_signal_111 ;
    wire new_AGEMA_signal_112 ;
    wire new_AGEMA_signal_113 ;
    wire new_AGEMA_signal_114 ;
    wire new_AGEMA_signal_115 ;
    wire new_AGEMA_signal_116 ;
    wire new_AGEMA_signal_117 ;
    wire new_AGEMA_signal_118 ;
    wire new_AGEMA_signal_119 ;
    wire new_AGEMA_signal_120 ;
    wire new_AGEMA_signal_121 ;
    wire new_AGEMA_signal_122 ;
    wire new_AGEMA_signal_123 ;
    wire new_AGEMA_signal_124 ;
    wire new_AGEMA_signal_125 ;
    wire new_AGEMA_signal_272 ;
    wire new_AGEMA_signal_273 ;
    wire new_AGEMA_signal_274 ;
    wire new_AGEMA_signal_275 ;
    wire new_AGEMA_signal_276 ;
    wire new_AGEMA_signal_277 ;
    wire new_AGEMA_signal_278 ;
    wire new_AGEMA_signal_279 ;
    wire new_AGEMA_signal_280 ;
    wire new_AGEMA_signal_281 ;
    wire new_AGEMA_signal_282 ;
    wire new_AGEMA_signal_283 ;
    wire new_AGEMA_signal_284 ;
    wire new_AGEMA_signal_285 ;
    wire new_AGEMA_signal_286 ;
    wire new_AGEMA_signal_287 ;
    wire new_AGEMA_signal_288 ;
    wire new_AGEMA_signal_289 ;
    wire new_AGEMA_signal_290 ;
    wire new_AGEMA_signal_291 ;
    wire new_AGEMA_signal_292 ;
    wire new_AGEMA_signal_293 ;
    wire new_AGEMA_signal_294 ;
    wire new_AGEMA_signal_295 ;
    wire new_AGEMA_signal_296 ;
    wire new_AGEMA_signal_297 ;
    wire new_AGEMA_signal_298 ;
    wire new_AGEMA_signal_299 ;
    wire new_AGEMA_signal_300 ;
    wire new_AGEMA_signal_301 ;
    wire new_AGEMA_signal_302 ;
    wire new_AGEMA_signal_303 ;
    wire new_AGEMA_signal_304 ;
    wire new_AGEMA_signal_305 ;
    wire new_AGEMA_signal_306 ;
    wire new_AGEMA_signal_307 ;
    wire new_AGEMA_signal_308 ;
    wire new_AGEMA_signal_309 ;
    wire new_AGEMA_signal_310 ;
    wire new_AGEMA_signal_311 ;
    wire new_AGEMA_signal_312 ;
    wire new_AGEMA_signal_313 ;
    wire new_AGEMA_signal_314 ;
    wire new_AGEMA_signal_315 ;
    wire new_AGEMA_signal_316 ;
    wire new_AGEMA_signal_317 ;
    wire new_AGEMA_signal_318 ;
    wire new_AGEMA_signal_319 ;
    wire new_AGEMA_signal_320 ;
    wire new_AGEMA_signal_321 ;
    wire new_AGEMA_signal_322 ;
    wire new_AGEMA_signal_323 ;
    wire new_AGEMA_signal_324 ;
    wire new_AGEMA_signal_325 ;
    wire new_AGEMA_signal_326 ;
    wire new_AGEMA_signal_327 ;
    wire new_AGEMA_signal_328 ;
    wire new_AGEMA_signal_329 ;
    wire new_AGEMA_signal_330 ;
    wire new_AGEMA_signal_331 ;
    wire new_AGEMA_signal_332 ;
    wire new_AGEMA_signal_333 ;
    wire new_AGEMA_signal_334 ;
    wire new_AGEMA_signal_335 ;
    wire new_AGEMA_signal_336 ;
    wire new_AGEMA_signal_337 ;
    wire new_AGEMA_signal_338 ;
    wire new_AGEMA_signal_339 ;
    wire new_AGEMA_signal_340 ;
    wire new_AGEMA_signal_341 ;
    wire new_AGEMA_signal_342 ;
    wire new_AGEMA_signal_343 ;
    wire new_AGEMA_signal_344 ;
    wire new_AGEMA_signal_345 ;
    wire new_AGEMA_signal_346 ;
    wire new_AGEMA_signal_347 ;
    wire new_AGEMA_signal_348 ;
    wire new_AGEMA_signal_349 ;
    wire new_AGEMA_signal_350 ;
    wire new_AGEMA_signal_351 ;
    wire new_AGEMA_signal_352 ;
    wire new_AGEMA_signal_353 ;
    wire new_AGEMA_signal_354 ;
    wire new_AGEMA_signal_355 ;
    wire new_AGEMA_signal_356 ;
    wire new_AGEMA_signal_357 ;
    wire new_AGEMA_signal_358 ;
    wire new_AGEMA_signal_359 ;
    wire new_AGEMA_signal_360 ;
    wire new_AGEMA_signal_361 ;
    wire new_AGEMA_signal_362 ;
    wire new_AGEMA_signal_363 ;
    wire new_AGEMA_signal_364 ;
    wire new_AGEMA_signal_365 ;
    wire new_AGEMA_signal_366 ;
    wire new_AGEMA_signal_367 ;
    wire new_AGEMA_signal_368 ;
    wire new_AGEMA_signal_369 ;
    wire new_AGEMA_signal_370 ;
    wire new_AGEMA_signal_371 ;
    wire new_AGEMA_signal_372 ;
    wire new_AGEMA_signal_373 ;
    wire new_AGEMA_signal_374 ;
    wire new_AGEMA_signal_375 ;
    wire new_AGEMA_signal_376 ;
    wire new_AGEMA_signal_377 ;
    wire new_AGEMA_signal_378 ;
    wire new_AGEMA_signal_379 ;
    wire new_AGEMA_signal_380 ;
    wire new_AGEMA_signal_381 ;
    wire new_AGEMA_signal_382 ;
    wire new_AGEMA_signal_383 ;
    wire new_AGEMA_signal_384 ;
    wire new_AGEMA_signal_385 ;
    wire new_AGEMA_signal_386 ;
    wire new_AGEMA_signal_387 ;
    wire new_AGEMA_signal_388 ;
    wire new_AGEMA_signal_389 ;
    wire new_AGEMA_signal_390 ;
    wire new_AGEMA_signal_391 ;
    wire new_AGEMA_signal_392 ;
    wire new_AGEMA_signal_393 ;
    wire new_AGEMA_signal_394 ;
    wire new_AGEMA_signal_395 ;
    wire new_AGEMA_signal_396 ;
    wire new_AGEMA_signal_397 ;
    wire new_AGEMA_signal_398 ;
    wire new_AGEMA_signal_399 ;
    wire new_AGEMA_signal_400 ;
    wire new_AGEMA_signal_401 ;
    wire new_AGEMA_signal_402 ;
    wire new_AGEMA_signal_403 ;
    wire new_AGEMA_signal_404 ;
    wire new_AGEMA_signal_405 ;
    wire new_AGEMA_signal_406 ;
    wire new_AGEMA_signal_407 ;
    wire new_AGEMA_signal_408 ;
    wire new_AGEMA_signal_409 ;
    wire new_AGEMA_signal_410 ;
    wire new_AGEMA_signal_411 ;
    wire new_AGEMA_signal_412 ;
    wire new_AGEMA_signal_413 ;
    wire new_AGEMA_signal_414 ;
    wire new_AGEMA_signal_415 ;
    wire new_AGEMA_signal_416 ;
    wire new_AGEMA_signal_417 ;
    wire new_AGEMA_signal_418 ;
    wire new_AGEMA_signal_419 ;
    wire new_AGEMA_signal_420 ;
    wire new_AGEMA_signal_421 ;
    wire new_AGEMA_signal_422 ;
    wire new_AGEMA_signal_423 ;
    wire new_AGEMA_signal_424 ;
    wire new_AGEMA_signal_425 ;
    wire new_AGEMA_signal_426 ;
    wire new_AGEMA_signal_427 ;
    wire new_AGEMA_signal_428 ;
    wire new_AGEMA_signal_429 ;
    wire new_AGEMA_signal_430 ;
    wire new_AGEMA_signal_431 ;
    wire new_AGEMA_signal_432 ;
    wire new_AGEMA_signal_433 ;
    wire new_AGEMA_signal_434 ;
    wire new_AGEMA_signal_435 ;
    wire new_AGEMA_signal_436 ;
    wire new_AGEMA_signal_437 ;
    wire new_AGEMA_signal_438 ;
    wire new_AGEMA_signal_439 ;
    wire new_AGEMA_signal_440 ;
    wire new_AGEMA_signal_441 ;
    wire new_AGEMA_signal_442 ;
    wire new_AGEMA_signal_443 ;
    wire new_AGEMA_signal_444 ;
    wire new_AGEMA_signal_445 ;
    wire new_AGEMA_signal_446 ;
    wire new_AGEMA_signal_447 ;
    wire new_AGEMA_signal_448 ;
    wire new_AGEMA_signal_449 ;
    wire new_AGEMA_signal_450 ;
    wire new_AGEMA_signal_451 ;
    wire new_AGEMA_signal_452 ;
    wire new_AGEMA_signal_453 ;
    wire new_AGEMA_signal_454 ;
    wire new_AGEMA_signal_455 ;
    wire new_AGEMA_signal_456 ;
    wire new_AGEMA_signal_457 ;
    wire new_AGEMA_signal_458 ;
    wire new_AGEMA_signal_459 ;
    wire new_AGEMA_signal_460 ;
    wire new_AGEMA_signal_461 ;
    wire new_AGEMA_signal_462 ;
    wire new_AGEMA_signal_463 ;
    wire new_AGEMA_signal_464 ;
    wire new_AGEMA_signal_465 ;
    wire new_AGEMA_signal_466 ;
    wire new_AGEMA_signal_467 ;
    wire new_AGEMA_signal_468 ;
    wire new_AGEMA_signal_469 ;
    wire new_AGEMA_signal_470 ;
    wire new_AGEMA_signal_471 ;
    wire new_AGEMA_signal_472 ;
    wire new_AGEMA_signal_473 ;
    wire new_AGEMA_signal_474 ;
    wire new_AGEMA_signal_475 ;
    wire new_AGEMA_signal_476 ;
    wire new_AGEMA_signal_477 ;
    wire new_AGEMA_signal_478 ;
    wire new_AGEMA_signal_479 ;
    wire new_AGEMA_signal_480 ;
    wire new_AGEMA_signal_481 ;

    /* cells in depth 0 */
    not_masked #(.security_order(4), .pipeline(1)) U50 ( .a ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_41, new_AGEMA_signal_40, new_AGEMA_signal_39, new_AGEMA_signal_38, n53}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U53 ( .a ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_61, new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n52}) ) ;
    not_masked #(.security_order(4), .pipeline(1)) U59 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, new_AGEMA_signal_66, n51}) ) ;

    /* cells in depth 1 */
    buf_clk new_AGEMA_reg_buffer_23 ( .C ( clk ), .D ( SI_s0[3] ), .Q ( new_AGEMA_signal_272 ) ) ;
    buf_clk new_AGEMA_reg_buffer_25 ( .C ( clk ), .D ( SI_s1[3] ), .Q ( new_AGEMA_signal_274 ) ) ;
    buf_clk new_AGEMA_reg_buffer_27 ( .C ( clk ), .D ( SI_s2[3] ), .Q ( new_AGEMA_signal_276 ) ) ;
    buf_clk new_AGEMA_reg_buffer_29 ( .C ( clk ), .D ( SI_s3[3] ), .Q ( new_AGEMA_signal_278 ) ) ;
    buf_clk new_AGEMA_reg_buffer_31 ( .C ( clk ), .D ( SI_s4[3] ), .Q ( new_AGEMA_signal_280 ) ) ;
    buf_clk new_AGEMA_reg_buffer_33 ( .C ( clk ), .D ( n53 ), .Q ( new_AGEMA_signal_282 ) ) ;
    buf_clk new_AGEMA_reg_buffer_35 ( .C ( clk ), .D ( new_AGEMA_signal_38 ), .Q ( new_AGEMA_signal_284 ) ) ;
    buf_clk new_AGEMA_reg_buffer_37 ( .C ( clk ), .D ( new_AGEMA_signal_39 ), .Q ( new_AGEMA_signal_286 ) ) ;
    buf_clk new_AGEMA_reg_buffer_39 ( .C ( clk ), .D ( new_AGEMA_signal_40 ), .Q ( new_AGEMA_signal_288 ) ) ;
    buf_clk new_AGEMA_reg_buffer_41 ( .C ( clk ), .D ( new_AGEMA_signal_41 ), .Q ( new_AGEMA_signal_290 ) ) ;
    buf_clk new_AGEMA_reg_buffer_43 ( .C ( clk ), .D ( SI_s0[1] ), .Q ( new_AGEMA_signal_292 ) ) ;
    buf_clk new_AGEMA_reg_buffer_45 ( .C ( clk ), .D ( SI_s1[1] ), .Q ( new_AGEMA_signal_294 ) ) ;
    buf_clk new_AGEMA_reg_buffer_47 ( .C ( clk ), .D ( SI_s2[1] ), .Q ( new_AGEMA_signal_296 ) ) ;
    buf_clk new_AGEMA_reg_buffer_49 ( .C ( clk ), .D ( SI_s3[1] ), .Q ( new_AGEMA_signal_298 ) ) ;
    buf_clk new_AGEMA_reg_buffer_51 ( .C ( clk ), .D ( SI_s4[1] ), .Q ( new_AGEMA_signal_300 ) ) ;
    buf_clk new_AGEMA_reg_buffer_53 ( .C ( clk ), .D ( SI_s0[2] ), .Q ( new_AGEMA_signal_302 ) ) ;
    buf_clk new_AGEMA_reg_buffer_55 ( .C ( clk ), .D ( SI_s1[2] ), .Q ( new_AGEMA_signal_304 ) ) ;
    buf_clk new_AGEMA_reg_buffer_57 ( .C ( clk ), .D ( SI_s2[2] ), .Q ( new_AGEMA_signal_306 ) ) ;
    buf_clk new_AGEMA_reg_buffer_59 ( .C ( clk ), .D ( SI_s3[2] ), .Q ( new_AGEMA_signal_308 ) ) ;
    buf_clk new_AGEMA_reg_buffer_61 ( .C ( clk ), .D ( SI_s4[2] ), .Q ( new_AGEMA_signal_310 ) ) ;

    /* cells in depth 2 */
    nor_HPC2 #(.security_order(4), .pipeline(1)) U51 ( .a ({SI_s4[1], SI_s3[1], SI_s2[1], SI_s1[1], SI_s0[1]}), .b ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ({Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_53, new_AGEMA_signal_52, new_AGEMA_signal_51, new_AGEMA_signal_50, n40}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) U52 ( .a ({new_AGEMA_signal_53, new_AGEMA_signal_52, new_AGEMA_signal_51, new_AGEMA_signal_50, n40}), .b ({new_AGEMA_signal_281, new_AGEMA_signal_279, new_AGEMA_signal_277, new_AGEMA_signal_275, new_AGEMA_signal_273}), .c ({new_AGEMA_signal_77, new_AGEMA_signal_76, new_AGEMA_signal_75, new_AGEMA_signal_74, N12}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) U54 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_61, new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n52}), .clk ( clk ), .r ({Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10]}), .c ({new_AGEMA_signal_81, new_AGEMA_signal_80, new_AGEMA_signal_79, new_AGEMA_signal_78, n41}) ) ;
    xnor_HPC2 #(.security_order(4), .pipeline(1)) U55 ( .a ({new_AGEMA_signal_291, new_AGEMA_signal_289, new_AGEMA_signal_287, new_AGEMA_signal_285, new_AGEMA_signal_283}), .b ({new_AGEMA_signal_81, new_AGEMA_signal_80, new_AGEMA_signal_79, new_AGEMA_signal_78, n41}), .c ({new_AGEMA_signal_105, new_AGEMA_signal_104, new_AGEMA_signal_103, new_AGEMA_signal_102, n42}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) U57 ( .a ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .b ({SI_s4[3], SI_s3[3], SI_s2[3], SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ({Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20]}), .c ({new_AGEMA_signal_65, new_AGEMA_signal_64, new_AGEMA_signal_63, new_AGEMA_signal_62, n43}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) U60 ( .a ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, new_AGEMA_signal_66, n51}), .b ({new_AGEMA_signal_41, new_AGEMA_signal_40, new_AGEMA_signal_39, new_AGEMA_signal_38, n53}), .clk ( clk ), .r ({Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30]}), .c ({new_AGEMA_signal_89, new_AGEMA_signal_88, new_AGEMA_signal_87, new_AGEMA_signal_86, n45}) ) ;
    nor_HPC2 #(.security_order(4), .pipeline(1)) U61 ( .a ({SI_s4[2], SI_s3[2], SI_s2[2], SI_s1[2], SI_s0[2]}), .b ({SI_s4[0], SI_s3[0], SI_s2[0], SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ({Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40]}), .c ({new_AGEMA_signal_73, new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, n48}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) U67 ( .a ({new_AGEMA_signal_61, new_AGEMA_signal_60, new_AGEMA_signal_59, new_AGEMA_signal_58, n52}), .b ({new_AGEMA_signal_69, new_AGEMA_signal_68, new_AGEMA_signal_67, new_AGEMA_signal_66, n51}), .clk ( clk ), .r ({Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50]}), .c ({new_AGEMA_signal_101, new_AGEMA_signal_100, new_AGEMA_signal_99, new_AGEMA_signal_98, n54}) ) ;
    xor_HPC2 #(.security_order(4), .pipeline(1)) U68 ( .a ({new_AGEMA_signal_101, new_AGEMA_signal_100, new_AGEMA_signal_99, new_AGEMA_signal_98, n54}), .b ({new_AGEMA_signal_291, new_AGEMA_signal_289, new_AGEMA_signal_287, new_AGEMA_signal_285, new_AGEMA_signal_283}), .c ({new_AGEMA_signal_113, new_AGEMA_signal_112, new_AGEMA_signal_111, new_AGEMA_signal_110, N9}) ) ;
    buf_clk new_AGEMA_reg_buffer_24 ( .C ( clk ), .D ( new_AGEMA_signal_272 ), .Q ( new_AGEMA_signal_273 ) ) ;
    buf_clk new_AGEMA_reg_buffer_26 ( .C ( clk ), .D ( new_AGEMA_signal_274 ), .Q ( new_AGEMA_signal_275 ) ) ;
    buf_clk new_AGEMA_reg_buffer_28 ( .C ( clk ), .D ( new_AGEMA_signal_276 ), .Q ( new_AGEMA_signal_277 ) ) ;
    buf_clk new_AGEMA_reg_buffer_30 ( .C ( clk ), .D ( new_AGEMA_signal_278 ), .Q ( new_AGEMA_signal_279 ) ) ;
    buf_clk new_AGEMA_reg_buffer_32 ( .C ( clk ), .D ( new_AGEMA_signal_280 ), .Q ( new_AGEMA_signal_281 ) ) ;
    buf_clk new_AGEMA_reg_buffer_34 ( .C ( clk ), .D ( new_AGEMA_signal_282 ), .Q ( new_AGEMA_signal_283 ) ) ;
    buf_clk new_AGEMA_reg_buffer_36 ( .C ( clk ), .D ( new_AGEMA_signal_284 ), .Q ( new_AGEMA_signal_285 ) ) ;
    buf_clk new_AGEMA_reg_buffer_38 ( .C ( clk ), .D ( new_AGEMA_signal_286 ), .Q ( new_AGEMA_signal_287 ) ) ;
    buf_clk new_AGEMA_reg_buffer_40 ( .C ( clk ), .D ( new_AGEMA_signal_288 ), .Q ( new_AGEMA_signal_289 ) ) ;
    buf_clk new_AGEMA_reg_buffer_42 ( .C ( clk ), .D ( new_AGEMA_signal_290 ), .Q ( new_AGEMA_signal_291 ) ) ;
    buf_clk new_AGEMA_reg_buffer_44 ( .C ( clk ), .D ( new_AGEMA_signal_292 ), .Q ( new_AGEMA_signal_293 ) ) ;
    buf_clk new_AGEMA_reg_buffer_46 ( .C ( clk ), .D ( new_AGEMA_signal_294 ), .Q ( new_AGEMA_signal_295 ) ) ;
    buf_clk new_AGEMA_reg_buffer_48 ( .C ( clk ), .D ( new_AGEMA_signal_296 ), .Q ( new_AGEMA_signal_297 ) ) ;
    buf_clk new_AGEMA_reg_buffer_50 ( .C ( clk ), .D ( new_AGEMA_signal_298 ), .Q ( new_AGEMA_signal_299 ) ) ;
    buf_clk new_AGEMA_reg_buffer_52 ( .C ( clk ), .D ( new_AGEMA_signal_300 ), .Q ( new_AGEMA_signal_301 ) ) ;
    buf_clk new_AGEMA_reg_buffer_54 ( .C ( clk ), .D ( new_AGEMA_signal_302 ), .Q ( new_AGEMA_signal_303 ) ) ;
    buf_clk new_AGEMA_reg_buffer_56 ( .C ( clk ), .D ( new_AGEMA_signal_304 ), .Q ( new_AGEMA_signal_305 ) ) ;
    buf_clk new_AGEMA_reg_buffer_58 ( .C ( clk ), .D ( new_AGEMA_signal_306 ), .Q ( new_AGEMA_signal_307 ) ) ;
    buf_clk new_AGEMA_reg_buffer_60 ( .C ( clk ), .D ( new_AGEMA_signal_308 ), .Q ( new_AGEMA_signal_309 ) ) ;
    buf_clk new_AGEMA_reg_buffer_62 ( .C ( clk ), .D ( new_AGEMA_signal_310 ), .Q ( new_AGEMA_signal_311 ) ) ;

    /* cells in depth 3 */
    buf_clk new_AGEMA_reg_buffer_63 ( .C ( clk ), .D ( n45 ), .Q ( new_AGEMA_signal_312 ) ) ;
    buf_clk new_AGEMA_reg_buffer_65 ( .C ( clk ), .D ( new_AGEMA_signal_86 ), .Q ( new_AGEMA_signal_314 ) ) ;
    buf_clk new_AGEMA_reg_buffer_67 ( .C ( clk ), .D ( new_AGEMA_signal_87 ), .Q ( new_AGEMA_signal_316 ) ) ;
    buf_clk new_AGEMA_reg_buffer_69 ( .C ( clk ), .D ( new_AGEMA_signal_88 ), .Q ( new_AGEMA_signal_318 ) ) ;
    buf_clk new_AGEMA_reg_buffer_71 ( .C ( clk ), .D ( new_AGEMA_signal_89 ), .Q ( new_AGEMA_signal_320 ) ) ;
    buf_clk new_AGEMA_reg_buffer_73 ( .C ( clk ), .D ( new_AGEMA_signal_293 ), .Q ( new_AGEMA_signal_322 ) ) ;
    buf_clk new_AGEMA_reg_buffer_77 ( .C ( clk ), .D ( new_AGEMA_signal_295 ), .Q ( new_AGEMA_signal_326 ) ) ;
    buf_clk new_AGEMA_reg_buffer_81 ( .C ( clk ), .D ( new_AGEMA_signal_297 ), .Q ( new_AGEMA_signal_330 ) ) ;
    buf_clk new_AGEMA_reg_buffer_85 ( .C ( clk ), .D ( new_AGEMA_signal_299 ), .Q ( new_AGEMA_signal_334 ) ) ;
    buf_clk new_AGEMA_reg_buffer_89 ( .C ( clk ), .D ( new_AGEMA_signal_301 ), .Q ( new_AGEMA_signal_338 ) ) ;
    buf_clk new_AGEMA_reg_buffer_123 ( .C ( clk ), .D ( N9 ), .Q ( new_AGEMA_signal_372 ) ) ;
    buf_clk new_AGEMA_reg_buffer_131 ( .C ( clk ), .D ( new_AGEMA_signal_110 ), .Q ( new_AGEMA_signal_380 ) ) ;
    buf_clk new_AGEMA_reg_buffer_139 ( .C ( clk ), .D ( new_AGEMA_signal_111 ), .Q ( new_AGEMA_signal_388 ) ) ;
    buf_clk new_AGEMA_reg_buffer_147 ( .C ( clk ), .D ( new_AGEMA_signal_112 ), .Q ( new_AGEMA_signal_396 ) ) ;
    buf_clk new_AGEMA_reg_buffer_155 ( .C ( clk ), .D ( new_AGEMA_signal_113 ), .Q ( new_AGEMA_signal_404 ) ) ;
    buf_clk new_AGEMA_reg_buffer_163 ( .C ( clk ), .D ( N12 ), .Q ( new_AGEMA_signal_412 ) ) ;
    buf_clk new_AGEMA_reg_buffer_171 ( .C ( clk ), .D ( new_AGEMA_signal_74 ), .Q ( new_AGEMA_signal_420 ) ) ;
    buf_clk new_AGEMA_reg_buffer_179 ( .C ( clk ), .D ( new_AGEMA_signal_75 ), .Q ( new_AGEMA_signal_428 ) ) ;
    buf_clk new_AGEMA_reg_buffer_187 ( .C ( clk ), .D ( new_AGEMA_signal_76 ), .Q ( new_AGEMA_signal_436 ) ) ;
    buf_clk new_AGEMA_reg_buffer_195 ( .C ( clk ), .D ( new_AGEMA_signal_77 ), .Q ( new_AGEMA_signal_444 ) ) ;

    /* cells in depth 4 */
    mux2_HPC2 #(.security_order(4), .pipeline(1)) U56 ( .s ({new_AGEMA_signal_301, new_AGEMA_signal_299, new_AGEMA_signal_297, new_AGEMA_signal_295, new_AGEMA_signal_293}), .b ({new_AGEMA_signal_105, new_AGEMA_signal_104, new_AGEMA_signal_103, new_AGEMA_signal_102, n42}), .a ({new_AGEMA_signal_311, new_AGEMA_signal_309, new_AGEMA_signal_307, new_AGEMA_signal_305, new_AGEMA_signal_303}), .clk ( clk ), .r ({Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60]}), .c ({new_AGEMA_signal_117, new_AGEMA_signal_116, new_AGEMA_signal_115, new_AGEMA_signal_114, N19}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) U58 ( .a ({new_AGEMA_signal_65, new_AGEMA_signal_64, new_AGEMA_signal_63, new_AGEMA_signal_62, n43}), .b ({new_AGEMA_signal_311, new_AGEMA_signal_309, new_AGEMA_signal_307, new_AGEMA_signal_305, new_AGEMA_signal_303}), .clk ( clk ), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70]}), .c ({new_AGEMA_signal_85, new_AGEMA_signal_84, new_AGEMA_signal_83, new_AGEMA_signal_82, n47}) ) ;
    or_HPC2 #(.security_order(4), .pipeline(1)) U62 ( .a ({new_AGEMA_signal_281, new_AGEMA_signal_279, new_AGEMA_signal_277, new_AGEMA_signal_275, new_AGEMA_signal_273}), .b ({new_AGEMA_signal_73, new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, n48}), .clk ( clk ), .r ({Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .c ({new_AGEMA_signal_93, new_AGEMA_signal_92, new_AGEMA_signal_91, new_AGEMA_signal_90, n44}) ) ;
    nand_HPC2 #(.security_order(4), .pipeline(1)) U65 ( .a ({new_AGEMA_signal_281, new_AGEMA_signal_279, new_AGEMA_signal_277, new_AGEMA_signal_275, new_AGEMA_signal_273}), .b ({new_AGEMA_signal_73, new_AGEMA_signal_72, new_AGEMA_signal_71, new_AGEMA_signal_70, n48}), .clk ( clk ), .r ({Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90]}), .c ({new_AGEMA_signal_97, new_AGEMA_signal_96, new_AGEMA_signal_95, new_AGEMA_signal_94, n49}) ) ;
    buf_clk new_AGEMA_reg_buffer_64 ( .C ( clk ), .D ( new_AGEMA_signal_312 ), .Q ( new_AGEMA_signal_313 ) ) ;
    buf_clk new_AGEMA_reg_buffer_66 ( .C ( clk ), .D ( new_AGEMA_signal_314 ), .Q ( new_AGEMA_signal_315 ) ) ;
    buf_clk new_AGEMA_reg_buffer_68 ( .C ( clk ), .D ( new_AGEMA_signal_316 ), .Q ( new_AGEMA_signal_317 ) ) ;
    buf_clk new_AGEMA_reg_buffer_70 ( .C ( clk ), .D ( new_AGEMA_signal_318 ), .Q ( new_AGEMA_signal_319 ) ) ;
    buf_clk new_AGEMA_reg_buffer_72 ( .C ( clk ), .D ( new_AGEMA_signal_320 ), .Q ( new_AGEMA_signal_321 ) ) ;
    buf_clk new_AGEMA_reg_buffer_74 ( .C ( clk ), .D ( new_AGEMA_signal_322 ), .Q ( new_AGEMA_signal_323 ) ) ;
    buf_clk new_AGEMA_reg_buffer_78 ( .C ( clk ), .D ( new_AGEMA_signal_326 ), .Q ( new_AGEMA_signal_327 ) ) ;
    buf_clk new_AGEMA_reg_buffer_82 ( .C ( clk ), .D ( new_AGEMA_signal_330 ), .Q ( new_AGEMA_signal_331 ) ) ;
    buf_clk new_AGEMA_reg_buffer_86 ( .C ( clk ), .D ( new_AGEMA_signal_334 ), .Q ( new_AGEMA_signal_335 ) ) ;
    buf_clk new_AGEMA_reg_buffer_90 ( .C ( clk ), .D ( new_AGEMA_signal_338 ), .Q ( new_AGEMA_signal_339 ) ) ;
    buf_clk new_AGEMA_reg_buffer_124 ( .C ( clk ), .D ( new_AGEMA_signal_372 ), .Q ( new_AGEMA_signal_373 ) ) ;
    buf_clk new_AGEMA_reg_buffer_132 ( .C ( clk ), .D ( new_AGEMA_signal_380 ), .Q ( new_AGEMA_signal_381 ) ) ;
    buf_clk new_AGEMA_reg_buffer_140 ( .C ( clk ), .D ( new_AGEMA_signal_388 ), .Q ( new_AGEMA_signal_389 ) ) ;
    buf_clk new_AGEMA_reg_buffer_148 ( .C ( clk ), .D ( new_AGEMA_signal_396 ), .Q ( new_AGEMA_signal_397 ) ) ;
    buf_clk new_AGEMA_reg_buffer_156 ( .C ( clk ), .D ( new_AGEMA_signal_404 ), .Q ( new_AGEMA_signal_405 ) ) ;
    buf_clk new_AGEMA_reg_buffer_164 ( .C ( clk ), .D ( new_AGEMA_signal_412 ), .Q ( new_AGEMA_signal_413 ) ) ;
    buf_clk new_AGEMA_reg_buffer_172 ( .C ( clk ), .D ( new_AGEMA_signal_420 ), .Q ( new_AGEMA_signal_421 ) ) ;
    buf_clk new_AGEMA_reg_buffer_180 ( .C ( clk ), .D ( new_AGEMA_signal_428 ), .Q ( new_AGEMA_signal_429 ) ) ;
    buf_clk new_AGEMA_reg_buffer_188 ( .C ( clk ), .D ( new_AGEMA_signal_436 ), .Q ( new_AGEMA_signal_437 ) ) ;
    buf_clk new_AGEMA_reg_buffer_196 ( .C ( clk ), .D ( new_AGEMA_signal_444 ), .Q ( new_AGEMA_signal_445 ) ) ;

    /* cells in depth 5 */
    buf_clk new_AGEMA_reg_buffer_75 ( .C ( clk ), .D ( new_AGEMA_signal_323 ), .Q ( new_AGEMA_signal_324 ) ) ;
    buf_clk new_AGEMA_reg_buffer_79 ( .C ( clk ), .D ( new_AGEMA_signal_327 ), .Q ( new_AGEMA_signal_328 ) ) ;
    buf_clk new_AGEMA_reg_buffer_83 ( .C ( clk ), .D ( new_AGEMA_signal_331 ), .Q ( new_AGEMA_signal_332 ) ) ;
    buf_clk new_AGEMA_reg_buffer_87 ( .C ( clk ), .D ( new_AGEMA_signal_335 ), .Q ( new_AGEMA_signal_336 ) ) ;
    buf_clk new_AGEMA_reg_buffer_91 ( .C ( clk ), .D ( new_AGEMA_signal_339 ), .Q ( new_AGEMA_signal_340 ) ) ;
    buf_clk new_AGEMA_reg_buffer_93 ( .C ( clk ), .D ( n47 ), .Q ( new_AGEMA_signal_342 ) ) ;
    buf_clk new_AGEMA_reg_buffer_95 ( .C ( clk ), .D ( new_AGEMA_signal_82 ), .Q ( new_AGEMA_signal_344 ) ) ;
    buf_clk new_AGEMA_reg_buffer_97 ( .C ( clk ), .D ( new_AGEMA_signal_83 ), .Q ( new_AGEMA_signal_346 ) ) ;
    buf_clk new_AGEMA_reg_buffer_99 ( .C ( clk ), .D ( new_AGEMA_signal_84 ), .Q ( new_AGEMA_signal_348 ) ) ;
    buf_clk new_AGEMA_reg_buffer_101 ( .C ( clk ), .D ( new_AGEMA_signal_85 ), .Q ( new_AGEMA_signal_350 ) ) ;
    buf_clk new_AGEMA_reg_buffer_103 ( .C ( clk ), .D ( n49 ), .Q ( new_AGEMA_signal_352 ) ) ;
    buf_clk new_AGEMA_reg_buffer_107 ( .C ( clk ), .D ( new_AGEMA_signal_94 ), .Q ( new_AGEMA_signal_356 ) ) ;
    buf_clk new_AGEMA_reg_buffer_111 ( .C ( clk ), .D ( new_AGEMA_signal_95 ), .Q ( new_AGEMA_signal_360 ) ) ;
    buf_clk new_AGEMA_reg_buffer_115 ( .C ( clk ), .D ( new_AGEMA_signal_96 ), .Q ( new_AGEMA_signal_364 ) ) ;
    buf_clk new_AGEMA_reg_buffer_119 ( .C ( clk ), .D ( new_AGEMA_signal_97 ), .Q ( new_AGEMA_signal_368 ) ) ;
    buf_clk new_AGEMA_reg_buffer_125 ( .C ( clk ), .D ( new_AGEMA_signal_373 ), .Q ( new_AGEMA_signal_374 ) ) ;
    buf_clk new_AGEMA_reg_buffer_133 ( .C ( clk ), .D ( new_AGEMA_signal_381 ), .Q ( new_AGEMA_signal_382 ) ) ;
    buf_clk new_AGEMA_reg_buffer_141 ( .C ( clk ), .D ( new_AGEMA_signal_389 ), .Q ( new_AGEMA_signal_390 ) ) ;
    buf_clk new_AGEMA_reg_buffer_149 ( .C ( clk ), .D ( new_AGEMA_signal_397 ), .Q ( new_AGEMA_signal_398 ) ) ;
    buf_clk new_AGEMA_reg_buffer_157 ( .C ( clk ), .D ( new_AGEMA_signal_405 ), .Q ( new_AGEMA_signal_406 ) ) ;
    buf_clk new_AGEMA_reg_buffer_165 ( .C ( clk ), .D ( new_AGEMA_signal_413 ), .Q ( new_AGEMA_signal_414 ) ) ;
    buf_clk new_AGEMA_reg_buffer_173 ( .C ( clk ), .D ( new_AGEMA_signal_421 ), .Q ( new_AGEMA_signal_422 ) ) ;
    buf_clk new_AGEMA_reg_buffer_181 ( .C ( clk ), .D ( new_AGEMA_signal_429 ), .Q ( new_AGEMA_signal_430 ) ) ;
    buf_clk new_AGEMA_reg_buffer_189 ( .C ( clk ), .D ( new_AGEMA_signal_437 ), .Q ( new_AGEMA_signal_438 ) ) ;
    buf_clk new_AGEMA_reg_buffer_197 ( .C ( clk ), .D ( new_AGEMA_signal_445 ), .Q ( new_AGEMA_signal_446 ) ) ;
    buf_clk new_AGEMA_reg_buffer_203 ( .C ( clk ), .D ( N19 ), .Q ( new_AGEMA_signal_452 ) ) ;
    buf_clk new_AGEMA_reg_buffer_209 ( .C ( clk ), .D ( new_AGEMA_signal_114 ), .Q ( new_AGEMA_signal_458 ) ) ;
    buf_clk new_AGEMA_reg_buffer_215 ( .C ( clk ), .D ( new_AGEMA_signal_115 ), .Q ( new_AGEMA_signal_464 ) ) ;
    buf_clk new_AGEMA_reg_buffer_221 ( .C ( clk ), .D ( new_AGEMA_signal_116 ), .Q ( new_AGEMA_signal_470 ) ) ;
    buf_clk new_AGEMA_reg_buffer_227 ( .C ( clk ), .D ( new_AGEMA_signal_117 ), .Q ( new_AGEMA_signal_476 ) ) ;

    /* cells in depth 6 */
    nor_HPC2 #(.security_order(4), .pipeline(1)) U63 ( .a ({new_AGEMA_signal_321, new_AGEMA_signal_319, new_AGEMA_signal_317, new_AGEMA_signal_315, new_AGEMA_signal_313}), .b ({new_AGEMA_signal_93, new_AGEMA_signal_92, new_AGEMA_signal_91, new_AGEMA_signal_90, n44}), .clk ( clk ), .r ({Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100]}), .c ({new_AGEMA_signal_109, new_AGEMA_signal_108, new_AGEMA_signal_107, new_AGEMA_signal_106, n46}) ) ;
    buf_clk new_AGEMA_reg_buffer_76 ( .C ( clk ), .D ( new_AGEMA_signal_324 ), .Q ( new_AGEMA_signal_325 ) ) ;
    buf_clk new_AGEMA_reg_buffer_80 ( .C ( clk ), .D ( new_AGEMA_signal_328 ), .Q ( new_AGEMA_signal_329 ) ) ;
    buf_clk new_AGEMA_reg_buffer_84 ( .C ( clk ), .D ( new_AGEMA_signal_332 ), .Q ( new_AGEMA_signal_333 ) ) ;
    buf_clk new_AGEMA_reg_buffer_88 ( .C ( clk ), .D ( new_AGEMA_signal_336 ), .Q ( new_AGEMA_signal_337 ) ) ;
    buf_clk new_AGEMA_reg_buffer_92 ( .C ( clk ), .D ( new_AGEMA_signal_340 ), .Q ( new_AGEMA_signal_341 ) ) ;
    buf_clk new_AGEMA_reg_buffer_94 ( .C ( clk ), .D ( new_AGEMA_signal_342 ), .Q ( new_AGEMA_signal_343 ) ) ;
    buf_clk new_AGEMA_reg_buffer_96 ( .C ( clk ), .D ( new_AGEMA_signal_344 ), .Q ( new_AGEMA_signal_345 ) ) ;
    buf_clk new_AGEMA_reg_buffer_98 ( .C ( clk ), .D ( new_AGEMA_signal_346 ), .Q ( new_AGEMA_signal_347 ) ) ;
    buf_clk new_AGEMA_reg_buffer_100 ( .C ( clk ), .D ( new_AGEMA_signal_348 ), .Q ( new_AGEMA_signal_349 ) ) ;
    buf_clk new_AGEMA_reg_buffer_102 ( .C ( clk ), .D ( new_AGEMA_signal_350 ), .Q ( new_AGEMA_signal_351 ) ) ;
    buf_clk new_AGEMA_reg_buffer_104 ( .C ( clk ), .D ( new_AGEMA_signal_352 ), .Q ( new_AGEMA_signal_353 ) ) ;
    buf_clk new_AGEMA_reg_buffer_108 ( .C ( clk ), .D ( new_AGEMA_signal_356 ), .Q ( new_AGEMA_signal_357 ) ) ;
    buf_clk new_AGEMA_reg_buffer_112 ( .C ( clk ), .D ( new_AGEMA_signal_360 ), .Q ( new_AGEMA_signal_361 ) ) ;
    buf_clk new_AGEMA_reg_buffer_116 ( .C ( clk ), .D ( new_AGEMA_signal_364 ), .Q ( new_AGEMA_signal_365 ) ) ;
    buf_clk new_AGEMA_reg_buffer_120 ( .C ( clk ), .D ( new_AGEMA_signal_368 ), .Q ( new_AGEMA_signal_369 ) ) ;
    buf_clk new_AGEMA_reg_buffer_126 ( .C ( clk ), .D ( new_AGEMA_signal_374 ), .Q ( new_AGEMA_signal_375 ) ) ;
    buf_clk new_AGEMA_reg_buffer_134 ( .C ( clk ), .D ( new_AGEMA_signal_382 ), .Q ( new_AGEMA_signal_383 ) ) ;
    buf_clk new_AGEMA_reg_buffer_142 ( .C ( clk ), .D ( new_AGEMA_signal_390 ), .Q ( new_AGEMA_signal_391 ) ) ;
    buf_clk new_AGEMA_reg_buffer_150 ( .C ( clk ), .D ( new_AGEMA_signal_398 ), .Q ( new_AGEMA_signal_399 ) ) ;
    buf_clk new_AGEMA_reg_buffer_158 ( .C ( clk ), .D ( new_AGEMA_signal_406 ), .Q ( new_AGEMA_signal_407 ) ) ;
    buf_clk new_AGEMA_reg_buffer_166 ( .C ( clk ), .D ( new_AGEMA_signal_414 ), .Q ( new_AGEMA_signal_415 ) ) ;
    buf_clk new_AGEMA_reg_buffer_174 ( .C ( clk ), .D ( new_AGEMA_signal_422 ), .Q ( new_AGEMA_signal_423 ) ) ;
    buf_clk new_AGEMA_reg_buffer_182 ( .C ( clk ), .D ( new_AGEMA_signal_430 ), .Q ( new_AGEMA_signal_431 ) ) ;
    buf_clk new_AGEMA_reg_buffer_190 ( .C ( clk ), .D ( new_AGEMA_signal_438 ), .Q ( new_AGEMA_signal_439 ) ) ;
    buf_clk new_AGEMA_reg_buffer_198 ( .C ( clk ), .D ( new_AGEMA_signal_446 ), .Q ( new_AGEMA_signal_447 ) ) ;
    buf_clk new_AGEMA_reg_buffer_204 ( .C ( clk ), .D ( new_AGEMA_signal_452 ), .Q ( new_AGEMA_signal_453 ) ) ;
    buf_clk new_AGEMA_reg_buffer_210 ( .C ( clk ), .D ( new_AGEMA_signal_458 ), .Q ( new_AGEMA_signal_459 ) ) ;
    buf_clk new_AGEMA_reg_buffer_216 ( .C ( clk ), .D ( new_AGEMA_signal_464 ), .Q ( new_AGEMA_signal_465 ) ) ;
    buf_clk new_AGEMA_reg_buffer_222 ( .C ( clk ), .D ( new_AGEMA_signal_470 ), .Q ( new_AGEMA_signal_471 ) ) ;
    buf_clk new_AGEMA_reg_buffer_228 ( .C ( clk ), .D ( new_AGEMA_signal_476 ), .Q ( new_AGEMA_signal_477 ) ) ;

    /* cells in depth 7 */
    buf_clk new_AGEMA_reg_buffer_105 ( .C ( clk ), .D ( new_AGEMA_signal_353 ), .Q ( new_AGEMA_signal_354 ) ) ;
    buf_clk new_AGEMA_reg_buffer_109 ( .C ( clk ), .D ( new_AGEMA_signal_357 ), .Q ( new_AGEMA_signal_358 ) ) ;
    buf_clk new_AGEMA_reg_buffer_113 ( .C ( clk ), .D ( new_AGEMA_signal_361 ), .Q ( new_AGEMA_signal_362 ) ) ;
    buf_clk new_AGEMA_reg_buffer_117 ( .C ( clk ), .D ( new_AGEMA_signal_365 ), .Q ( new_AGEMA_signal_366 ) ) ;
    buf_clk new_AGEMA_reg_buffer_121 ( .C ( clk ), .D ( new_AGEMA_signal_369 ), .Q ( new_AGEMA_signal_370 ) ) ;
    buf_clk new_AGEMA_reg_buffer_127 ( .C ( clk ), .D ( new_AGEMA_signal_375 ), .Q ( new_AGEMA_signal_376 ) ) ;
    buf_clk new_AGEMA_reg_buffer_135 ( .C ( clk ), .D ( new_AGEMA_signal_383 ), .Q ( new_AGEMA_signal_384 ) ) ;
    buf_clk new_AGEMA_reg_buffer_143 ( .C ( clk ), .D ( new_AGEMA_signal_391 ), .Q ( new_AGEMA_signal_392 ) ) ;
    buf_clk new_AGEMA_reg_buffer_151 ( .C ( clk ), .D ( new_AGEMA_signal_399 ), .Q ( new_AGEMA_signal_400 ) ) ;
    buf_clk new_AGEMA_reg_buffer_159 ( .C ( clk ), .D ( new_AGEMA_signal_407 ), .Q ( new_AGEMA_signal_408 ) ) ;
    buf_clk new_AGEMA_reg_buffer_167 ( .C ( clk ), .D ( new_AGEMA_signal_415 ), .Q ( new_AGEMA_signal_416 ) ) ;
    buf_clk new_AGEMA_reg_buffer_175 ( .C ( clk ), .D ( new_AGEMA_signal_423 ), .Q ( new_AGEMA_signal_424 ) ) ;
    buf_clk new_AGEMA_reg_buffer_183 ( .C ( clk ), .D ( new_AGEMA_signal_431 ), .Q ( new_AGEMA_signal_432 ) ) ;
    buf_clk new_AGEMA_reg_buffer_191 ( .C ( clk ), .D ( new_AGEMA_signal_439 ), .Q ( new_AGEMA_signal_440 ) ) ;
    buf_clk new_AGEMA_reg_buffer_199 ( .C ( clk ), .D ( new_AGEMA_signal_447 ), .Q ( new_AGEMA_signal_448 ) ) ;
    buf_clk new_AGEMA_reg_buffer_205 ( .C ( clk ), .D ( new_AGEMA_signal_453 ), .Q ( new_AGEMA_signal_454 ) ) ;
    buf_clk new_AGEMA_reg_buffer_211 ( .C ( clk ), .D ( new_AGEMA_signal_459 ), .Q ( new_AGEMA_signal_460 ) ) ;
    buf_clk new_AGEMA_reg_buffer_217 ( .C ( clk ), .D ( new_AGEMA_signal_465 ), .Q ( new_AGEMA_signal_466 ) ) ;
    buf_clk new_AGEMA_reg_buffer_223 ( .C ( clk ), .D ( new_AGEMA_signal_471 ), .Q ( new_AGEMA_signal_472 ) ) ;
    buf_clk new_AGEMA_reg_buffer_229 ( .C ( clk ), .D ( new_AGEMA_signal_477 ), .Q ( new_AGEMA_signal_478 ) ) ;

    /* cells in depth 8 */
    mux2_HPC2 #(.security_order(4), .pipeline(1)) U64 ( .s ({new_AGEMA_signal_341, new_AGEMA_signal_337, new_AGEMA_signal_333, new_AGEMA_signal_329, new_AGEMA_signal_325}), .b ({new_AGEMA_signal_351, new_AGEMA_signal_349, new_AGEMA_signal_347, new_AGEMA_signal_345, new_AGEMA_signal_343}), .a ({new_AGEMA_signal_109, new_AGEMA_signal_108, new_AGEMA_signal_107, new_AGEMA_signal_106, n46}), .clk ( clk ), .r ({Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110]}), .c ({new_AGEMA_signal_121, new_AGEMA_signal_120, new_AGEMA_signal_119, new_AGEMA_signal_118, n50}) ) ;
    buf_clk new_AGEMA_reg_buffer_106 ( .C ( clk ), .D ( new_AGEMA_signal_354 ), .Q ( new_AGEMA_signal_355 ) ) ;
    buf_clk new_AGEMA_reg_buffer_110 ( .C ( clk ), .D ( new_AGEMA_signal_358 ), .Q ( new_AGEMA_signal_359 ) ) ;
    buf_clk new_AGEMA_reg_buffer_114 ( .C ( clk ), .D ( new_AGEMA_signal_362 ), .Q ( new_AGEMA_signal_363 ) ) ;
    buf_clk new_AGEMA_reg_buffer_118 ( .C ( clk ), .D ( new_AGEMA_signal_366 ), .Q ( new_AGEMA_signal_367 ) ) ;
    buf_clk new_AGEMA_reg_buffer_122 ( .C ( clk ), .D ( new_AGEMA_signal_370 ), .Q ( new_AGEMA_signal_371 ) ) ;
    buf_clk new_AGEMA_reg_buffer_128 ( .C ( clk ), .D ( new_AGEMA_signal_376 ), .Q ( new_AGEMA_signal_377 ) ) ;
    buf_clk new_AGEMA_reg_buffer_136 ( .C ( clk ), .D ( new_AGEMA_signal_384 ), .Q ( new_AGEMA_signal_385 ) ) ;
    buf_clk new_AGEMA_reg_buffer_144 ( .C ( clk ), .D ( new_AGEMA_signal_392 ), .Q ( new_AGEMA_signal_393 ) ) ;
    buf_clk new_AGEMA_reg_buffer_152 ( .C ( clk ), .D ( new_AGEMA_signal_400 ), .Q ( new_AGEMA_signal_401 ) ) ;
    buf_clk new_AGEMA_reg_buffer_160 ( .C ( clk ), .D ( new_AGEMA_signal_408 ), .Q ( new_AGEMA_signal_409 ) ) ;
    buf_clk new_AGEMA_reg_buffer_168 ( .C ( clk ), .D ( new_AGEMA_signal_416 ), .Q ( new_AGEMA_signal_417 ) ) ;
    buf_clk new_AGEMA_reg_buffer_176 ( .C ( clk ), .D ( new_AGEMA_signal_424 ), .Q ( new_AGEMA_signal_425 ) ) ;
    buf_clk new_AGEMA_reg_buffer_184 ( .C ( clk ), .D ( new_AGEMA_signal_432 ), .Q ( new_AGEMA_signal_433 ) ) ;
    buf_clk new_AGEMA_reg_buffer_192 ( .C ( clk ), .D ( new_AGEMA_signal_440 ), .Q ( new_AGEMA_signal_441 ) ) ;
    buf_clk new_AGEMA_reg_buffer_200 ( .C ( clk ), .D ( new_AGEMA_signal_448 ), .Q ( new_AGEMA_signal_449 ) ) ;
    buf_clk new_AGEMA_reg_buffer_206 ( .C ( clk ), .D ( new_AGEMA_signal_454 ), .Q ( new_AGEMA_signal_455 ) ) ;
    buf_clk new_AGEMA_reg_buffer_212 ( .C ( clk ), .D ( new_AGEMA_signal_460 ), .Q ( new_AGEMA_signal_461 ) ) ;
    buf_clk new_AGEMA_reg_buffer_218 ( .C ( clk ), .D ( new_AGEMA_signal_466 ), .Q ( new_AGEMA_signal_467 ) ) ;
    buf_clk new_AGEMA_reg_buffer_224 ( .C ( clk ), .D ( new_AGEMA_signal_472 ), .Q ( new_AGEMA_signal_473 ) ) ;
    buf_clk new_AGEMA_reg_buffer_230 ( .C ( clk ), .D ( new_AGEMA_signal_478 ), .Q ( new_AGEMA_signal_479 ) ) ;

    /* cells in depth 9 */
    buf_clk new_AGEMA_reg_buffer_129 ( .C ( clk ), .D ( new_AGEMA_signal_377 ), .Q ( new_AGEMA_signal_378 ) ) ;
    buf_clk new_AGEMA_reg_buffer_137 ( .C ( clk ), .D ( new_AGEMA_signal_385 ), .Q ( new_AGEMA_signal_386 ) ) ;
    buf_clk new_AGEMA_reg_buffer_145 ( .C ( clk ), .D ( new_AGEMA_signal_393 ), .Q ( new_AGEMA_signal_394 ) ) ;
    buf_clk new_AGEMA_reg_buffer_153 ( .C ( clk ), .D ( new_AGEMA_signal_401 ), .Q ( new_AGEMA_signal_402 ) ) ;
    buf_clk new_AGEMA_reg_buffer_161 ( .C ( clk ), .D ( new_AGEMA_signal_409 ), .Q ( new_AGEMA_signal_410 ) ) ;
    buf_clk new_AGEMA_reg_buffer_169 ( .C ( clk ), .D ( new_AGEMA_signal_417 ), .Q ( new_AGEMA_signal_418 ) ) ;
    buf_clk new_AGEMA_reg_buffer_177 ( .C ( clk ), .D ( new_AGEMA_signal_425 ), .Q ( new_AGEMA_signal_426 ) ) ;
    buf_clk new_AGEMA_reg_buffer_185 ( .C ( clk ), .D ( new_AGEMA_signal_433 ), .Q ( new_AGEMA_signal_434 ) ) ;
    buf_clk new_AGEMA_reg_buffer_193 ( .C ( clk ), .D ( new_AGEMA_signal_441 ), .Q ( new_AGEMA_signal_442 ) ) ;
    buf_clk new_AGEMA_reg_buffer_201 ( .C ( clk ), .D ( new_AGEMA_signal_449 ), .Q ( new_AGEMA_signal_450 ) ) ;
    buf_clk new_AGEMA_reg_buffer_207 ( .C ( clk ), .D ( new_AGEMA_signal_455 ), .Q ( new_AGEMA_signal_456 ) ) ;
    buf_clk new_AGEMA_reg_buffer_213 ( .C ( clk ), .D ( new_AGEMA_signal_461 ), .Q ( new_AGEMA_signal_462 ) ) ;
    buf_clk new_AGEMA_reg_buffer_219 ( .C ( clk ), .D ( new_AGEMA_signal_467 ), .Q ( new_AGEMA_signal_468 ) ) ;
    buf_clk new_AGEMA_reg_buffer_225 ( .C ( clk ), .D ( new_AGEMA_signal_473 ), .Q ( new_AGEMA_signal_474 ) ) ;
    buf_clk new_AGEMA_reg_buffer_231 ( .C ( clk ), .D ( new_AGEMA_signal_479 ), .Q ( new_AGEMA_signal_480 ) ) ;

    /* cells in depth 10 */
    nand_HPC2 #(.security_order(4), .pipeline(1)) U66 ( .a ({new_AGEMA_signal_121, new_AGEMA_signal_120, new_AGEMA_signal_119, new_AGEMA_signal_118, n50}), .b ({new_AGEMA_signal_371, new_AGEMA_signal_367, new_AGEMA_signal_363, new_AGEMA_signal_359, new_AGEMA_signal_355}), .clk ( clk ), .r ({Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120]}), .c ({new_AGEMA_signal_125, new_AGEMA_signal_124, new_AGEMA_signal_123, new_AGEMA_signal_122, N27}) ) ;
    buf_clk new_AGEMA_reg_buffer_130 ( .C ( clk ), .D ( new_AGEMA_signal_378 ), .Q ( new_AGEMA_signal_379 ) ) ;
    buf_clk new_AGEMA_reg_buffer_138 ( .C ( clk ), .D ( new_AGEMA_signal_386 ), .Q ( new_AGEMA_signal_387 ) ) ;
    buf_clk new_AGEMA_reg_buffer_146 ( .C ( clk ), .D ( new_AGEMA_signal_394 ), .Q ( new_AGEMA_signal_395 ) ) ;
    buf_clk new_AGEMA_reg_buffer_154 ( .C ( clk ), .D ( new_AGEMA_signal_402 ), .Q ( new_AGEMA_signal_403 ) ) ;
    buf_clk new_AGEMA_reg_buffer_162 ( .C ( clk ), .D ( new_AGEMA_signal_410 ), .Q ( new_AGEMA_signal_411 ) ) ;
    buf_clk new_AGEMA_reg_buffer_170 ( .C ( clk ), .D ( new_AGEMA_signal_418 ), .Q ( new_AGEMA_signal_419 ) ) ;
    buf_clk new_AGEMA_reg_buffer_178 ( .C ( clk ), .D ( new_AGEMA_signal_426 ), .Q ( new_AGEMA_signal_427 ) ) ;
    buf_clk new_AGEMA_reg_buffer_186 ( .C ( clk ), .D ( new_AGEMA_signal_434 ), .Q ( new_AGEMA_signal_435 ) ) ;
    buf_clk new_AGEMA_reg_buffer_194 ( .C ( clk ), .D ( new_AGEMA_signal_442 ), .Q ( new_AGEMA_signal_443 ) ) ;
    buf_clk new_AGEMA_reg_buffer_202 ( .C ( clk ), .D ( new_AGEMA_signal_450 ), .Q ( new_AGEMA_signal_451 ) ) ;
    buf_clk new_AGEMA_reg_buffer_208 ( .C ( clk ), .D ( new_AGEMA_signal_456 ), .Q ( new_AGEMA_signal_457 ) ) ;
    buf_clk new_AGEMA_reg_buffer_214 ( .C ( clk ), .D ( new_AGEMA_signal_462 ), .Q ( new_AGEMA_signal_463 ) ) ;
    buf_clk new_AGEMA_reg_buffer_220 ( .C ( clk ), .D ( new_AGEMA_signal_468 ), .Q ( new_AGEMA_signal_469 ) ) ;
    buf_clk new_AGEMA_reg_buffer_226 ( .C ( clk ), .D ( new_AGEMA_signal_474 ), .Q ( new_AGEMA_signal_475 ) ) ;
    buf_clk new_AGEMA_reg_buffer_232 ( .C ( clk ), .D ( new_AGEMA_signal_480 ), .Q ( new_AGEMA_signal_481 ) ) ;

    /* register cells */
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_3_ ( .clk ( clk ), .D ({new_AGEMA_signal_411, new_AGEMA_signal_403, new_AGEMA_signal_395, new_AGEMA_signal_387, new_AGEMA_signal_379}), .Q ({SO_s4[3], SO_s3[3], SO_s2[3], SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_2_ ( .clk ( clk ), .D ({new_AGEMA_signal_451, new_AGEMA_signal_443, new_AGEMA_signal_435, new_AGEMA_signal_427, new_AGEMA_signal_419}), .Q ({SO_s4[2], SO_s3[2], SO_s2[2], SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_1_ ( .clk ( clk ), .D ({new_AGEMA_signal_481, new_AGEMA_signal_475, new_AGEMA_signal_469, new_AGEMA_signal_463, new_AGEMA_signal_457}), .Q ({SO_s4[1], SO_s3[1], SO_s2[1], SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(4), .pipeline(1)) SO_reg_0_ ( .clk ( clk ), .D ({new_AGEMA_signal_125, new_AGEMA_signal_124, new_AGEMA_signal_123, new_AGEMA_signal_122, N27}), .Q ({SO_s4[0], SO_s3[0], SO_s2[0], SO_s1[0], SO_s0[0]}) ) ;
endmodule
