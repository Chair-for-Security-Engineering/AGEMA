////////////////////////////////////////////////////////////////////////////
// COMPANY : Ruhr University Bochum
// AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Low-Latency Hardware Private Circuits] https://eprint.iacr.org/2022/507
// /////////////////////////////////////////////////////////////////
//
// Copyright c 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// INCLUDING NEGLIGENCE OR OTHERWISE ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//
/* modified netlist. Source: module PRESENT in file /AGEMA/Designs/PRESENT_nibble-serial/AGEMA/PRESENT.v */
/* 2 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 3 register stage(s) in total */

module PRESENT_HPC3_Pipeline_d1 (data_in_s0, key_s0, clk, reset, data_in_s1, key_s1, Fresh, data_out_s0, done, data_out_s1);
    input [63:0] data_in_s0 ;
    input [79:0] key_s0 ;
    input clk ;
    input reset ;
    input [63:0] data_in_s1 ;
    input [79:0] key_s1 ;
    input [7:0] Fresh ;
    output [63:0] data_out_s0 ;
    output done ;
    output [63:0] data_out_s1 ;
    wire selSbox ;
    wire ctrlData_0_ ;
    wire intDone ;
    wire fsm_n15 ;
    wire fsm_n14 ;
    wire fsm_n13 ;
    wire fsm_n12 ;
    wire fsm_n11 ;
    wire fsm_n10 ;
    wire fsm_n9 ;
    wire fsm_n8 ;
    wire fsm_n7 ;
    wire fsm_n6 ;
    wire fsm_n4 ;
    wire fsm_n2 ;
    wire fsm_n5 ;
    wire fsm_n20 ;
    wire fsm_ps_state_0_ ;
    wire fsm_ps_state_1_ ;
    wire fsm_n21 ;
    wire fsm_n3 ;
    wire fsm_rst_countSerial ;
    wire fsm_en_countRound ;
    wire fsm_cnt_rnd_n33 ;
    wire fsm_cnt_rnd_n32 ;
    wire fsm_cnt_rnd_n31 ;
    wire fsm_cnt_rnd_n30 ;
    wire fsm_cnt_rnd_n29 ;
    wire fsm_cnt_rnd_n28 ;
    wire fsm_cnt_rnd_n27 ;
    wire fsm_cnt_rnd_n26 ;
    wire fsm_cnt_rnd_n23 ;
    wire fsm_cnt_rnd_n22 ;
    wire fsm_cnt_rnd_n21 ;
    wire fsm_cnt_rnd_n20 ;
    wire fsm_cnt_rnd_n19 ;
    wire fsm_cnt_rnd_n17 ;
    wire fsm_cnt_rnd_n15 ;
    wire fsm_cnt_rnd_n13 ;
    wire fsm_cnt_rnd_n12 ;
    wire fsm_cnt_rnd_n11 ;
    wire fsm_cnt_rnd_n10 ;
    wire fsm_cnt_rnd_n9 ;
    wire fsm_cnt_rnd_n8 ;
    wire fsm_cnt_rnd_n7 ;
    wire fsm_cnt_rnd_n6 ;
    wire fsm_cnt_rnd_n5 ;
    wire fsm_cnt_rnd_n3 ;
    wire fsm_cnt_rnd_n24 ;
    wire fsm_cnt_rnd_n41 ;
    wire fsm_cnt_rnd_n25 ;
    wire fsm_cnt_rnd_n1 ;
    wire fsm_cnt_rnd_n18 ;
    wire fsm_cnt_rnd_n16 ;
    wire fsm_cnt_rnd_n14 ;
    wire fsm_cnt_ser_n10 ;
    wire fsm_cnt_ser_n9 ;
    wire fsm_cnt_ser_n8 ;
    wire fsm_cnt_ser_n7 ;
    wire fsm_cnt_ser_n6 ;
    wire fsm_cnt_ser_n5 ;
    wire fsm_cnt_ser_n4 ;
    wire fsm_cnt_ser_n2 ;
    wire fsm_cnt_ser_n20 ;
    wire fsm_cnt_ser_n28 ;
    wire fsm_cnt_ser_n26 ;
    wire fsm_cnt_ser_n3 ;
    wire fsm_cnt_ser_n1 ;
    wire stateFF_state_n7 ;
    wire stateFF_state_n6 ;
    wire stateFF_state_n5 ;
    wire keyFF_keystate_n8 ;
    wire keyFF_keystate_n7 ;
    wire keyFF_keystate_n6 ;
    wire sboxInst_n3 ;
    wire sboxInst_n2 ;
    wire sboxInst_n1 ;
    wire sboxInst_L8 ;
    wire sboxInst_L7 ;
    wire sboxInst_T3 ;
    wire sboxInst_T1 ;
    wire sboxInst_Q7 ;
    wire sboxInst_Q6 ;
    wire sboxInst_L5 ;
    wire sboxInst_T2 ;
    wire sboxInst_L4 ;
    wire sboxInst_Q3 ;
    wire sboxInst_L3 ;
    wire sboxInst_Q2 ;
    wire sboxInst_T0 ;
    wire sboxInst_L2 ;
    wire sboxInst_L1 ;
    wire sboxInst_L0 ;
    wire [4:0] counter ;
    wire [3:0] serialIn ;
    wire [3:0] sboxOut ;
    wire [3:0] roundkey ;
    wire [3:1] keyRegKS ;
    wire [3:0] sboxIn ;
    wire [3:0] stateXORroundkey ;
    wire [3:0] fsm_countSerial ;
    wire [63:0] stateFF_inputPar ;
    wire [3:0] stateFF_state_gff_1_s_next_state ;
    wire [3:0] stateFF_state_gff_2_s_next_state ;
    wire [3:0] stateFF_state_gff_3_s_next_state ;
    wire [3:0] stateFF_state_gff_4_s_next_state ;
    wire [3:0] stateFF_state_gff_5_s_next_state ;
    wire [3:0] stateFF_state_gff_6_s_next_state ;
    wire [3:0] stateFF_state_gff_7_s_next_state ;
    wire [3:0] stateFF_state_gff_8_s_next_state ;
    wire [3:0] stateFF_state_gff_9_s_next_state ;
    wire [3:0] stateFF_state_gff_10_s_next_state ;
    wire [3:0] stateFF_state_gff_11_s_next_state ;
    wire [3:0] stateFF_state_gff_12_s_next_state ;
    wire [3:0] stateFF_state_gff_13_s_next_state ;
    wire [3:0] stateFF_state_gff_14_s_next_state ;
    wire [3:0] stateFF_state_gff_15_s_next_state ;
    wire [3:0] stateFF_state_gff_16_s_next_state ;
    wire [4:0] keyFF_counterAdd ;
    wire [75:3] keyFF_outputPar ;
    wire [79:0] keyFF_inputPar ;
    wire [3:0] keyFF_keystate_gff_1_s_next_state ;
    wire [3:0] keyFF_keystate_gff_2_s_next_state ;
    wire [3:0] keyFF_keystate_gff_3_s_next_state ;
    wire [3:0] keyFF_keystate_gff_4_s_next_state ;
    wire [3:0] keyFF_keystate_gff_5_s_next_state ;
    wire [3:0] keyFF_keystate_gff_6_s_next_state ;
    wire [3:0] keyFF_keystate_gff_7_s_next_state ;
    wire [3:0] keyFF_keystate_gff_8_s_next_state ;
    wire [3:0] keyFF_keystate_gff_9_s_next_state ;
    wire [3:0] keyFF_keystate_gff_10_s_next_state ;
    wire [3:0] keyFF_keystate_gff_11_s_next_state ;
    wire [3:0] keyFF_keystate_gff_12_s_next_state ;
    wire [3:0] keyFF_keystate_gff_13_s_next_state ;
    wire [3:0] keyFF_keystate_gff_14_s_next_state ;
    wire [3:0] keyFF_keystate_gff_15_s_next_state ;
    wire [3:0] keyFF_keystate_gff_16_s_next_state ;
    wire [3:0] keyFF_keystate_gff_17_s_next_state ;
    wire [3:0] keyFF_keystate_gff_18_s_next_state ;
    wire [3:0] keyFF_keystate_gff_19_s_next_state ;
    wire [3:0] keyFF_keystate_gff_20_s_next_state ;
    wire new_AGEMA_signal_856 ;
    wire new_AGEMA_signal_858 ;
    wire new_AGEMA_signal_859 ;
    wire new_AGEMA_signal_861 ;
    wire new_AGEMA_signal_862 ;
    wire new_AGEMA_signal_864 ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_867 ;
    wire new_AGEMA_signal_870 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_876 ;
    wire new_AGEMA_signal_879 ;
    wire new_AGEMA_signal_882 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_888 ;
    wire new_AGEMA_signal_891 ;
    wire new_AGEMA_signal_894 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_900 ;
    wire new_AGEMA_signal_903 ;
    wire new_AGEMA_signal_906 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_912 ;
    wire new_AGEMA_signal_914 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_920 ;
    wire new_AGEMA_signal_923 ;
    wire new_AGEMA_signal_926 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_932 ;
    wire new_AGEMA_signal_935 ;
    wire new_AGEMA_signal_938 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_944 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_950 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_956 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire new_AGEMA_signal_1869 ;
    wire new_AGEMA_signal_1870 ;
    wire new_AGEMA_signal_1871 ;
    wire new_AGEMA_signal_1872 ;
    wire new_AGEMA_signal_1873 ;
    wire new_AGEMA_signal_1874 ;
    wire new_AGEMA_signal_1875 ;
    wire new_AGEMA_signal_1876 ;
    wire new_AGEMA_signal_1877 ;
    wire new_AGEMA_signal_1878 ;
    wire new_AGEMA_signal_1879 ;
    wire new_AGEMA_signal_1880 ;
    wire new_AGEMA_signal_1881 ;
    wire new_AGEMA_signal_1882 ;
    wire new_AGEMA_signal_1883 ;
    wire new_AGEMA_signal_1884 ;
    wire new_AGEMA_signal_1885 ;
    wire new_AGEMA_signal_1886 ;
    wire new_AGEMA_signal_1887 ;
    wire new_AGEMA_signal_1888 ;
    wire new_AGEMA_signal_1889 ;
    wire new_AGEMA_signal_1890 ;
    wire new_AGEMA_signal_1891 ;
    wire new_AGEMA_signal_1892 ;
    wire new_AGEMA_signal_1893 ;
    wire new_AGEMA_signal_1894 ;
    wire new_AGEMA_signal_1895 ;
    wire new_AGEMA_signal_1896 ;
    wire new_AGEMA_signal_1897 ;
    wire new_AGEMA_signal_1898 ;
    wire new_AGEMA_signal_1899 ;
    wire new_AGEMA_signal_1900 ;
    wire new_AGEMA_signal_1901 ;
    wire new_AGEMA_signal_1902 ;
    wire new_AGEMA_signal_1903 ;
    wire new_AGEMA_signal_1904 ;
    wire new_AGEMA_signal_1905 ;
    wire new_AGEMA_signal_1906 ;
    wire new_AGEMA_signal_1907 ;
    wire new_AGEMA_signal_1908 ;
    wire new_AGEMA_signal_1909 ;
    wire new_AGEMA_signal_1910 ;
    wire new_AGEMA_signal_1911 ;
    wire new_AGEMA_signal_1912 ;
    wire new_AGEMA_signal_1913 ;
    wire new_AGEMA_signal_1914 ;
    wire new_AGEMA_signal_1915 ;
    wire new_AGEMA_signal_1916 ;
    wire new_AGEMA_signal_1917 ;
    wire new_AGEMA_signal_1918 ;
    wire new_AGEMA_signal_1919 ;
    wire new_AGEMA_signal_1920 ;
    wire new_AGEMA_signal_1921 ;
    wire new_AGEMA_signal_1922 ;
    wire new_AGEMA_signal_1923 ;
    wire new_AGEMA_signal_1924 ;
    wire new_AGEMA_signal_1925 ;
    wire new_AGEMA_signal_1926 ;
    wire new_AGEMA_signal_1927 ;
    wire new_AGEMA_signal_1928 ;
    wire new_AGEMA_signal_1929 ;
    wire new_AGEMA_signal_1930 ;
    wire new_AGEMA_signal_1931 ;
    wire new_AGEMA_signal_1932 ;
    wire new_AGEMA_signal_1933 ;
    wire new_AGEMA_signal_1934 ;
    wire new_AGEMA_signal_1935 ;
    wire new_AGEMA_signal_1936 ;
    wire new_AGEMA_signal_1937 ;
    wire new_AGEMA_signal_1938 ;
    wire new_AGEMA_signal_1939 ;
    wire new_AGEMA_signal_1940 ;
    wire new_AGEMA_signal_1941 ;
    wire new_AGEMA_signal_1942 ;
    wire new_AGEMA_signal_1943 ;
    wire new_AGEMA_signal_1944 ;
    wire new_AGEMA_signal_1945 ;
    wire new_AGEMA_signal_1946 ;
    wire new_AGEMA_signal_1947 ;
    wire new_AGEMA_signal_1948 ;
    wire new_AGEMA_signal_1949 ;
    wire new_AGEMA_signal_1950 ;
    wire new_AGEMA_signal_1951 ;
    wire new_AGEMA_signal_1952 ;
    wire new_AGEMA_signal_1953 ;
    wire new_AGEMA_signal_1954 ;
    wire new_AGEMA_signal_1955 ;
    wire new_AGEMA_signal_1956 ;
    wire new_AGEMA_signal_1957 ;
    wire new_AGEMA_signal_1958 ;
    wire new_AGEMA_signal_1959 ;
    wire new_AGEMA_signal_1960 ;
    wire new_AGEMA_signal_1961 ;
    wire new_AGEMA_signal_1962 ;
    wire new_AGEMA_signal_1963 ;
    wire new_AGEMA_signal_1964 ;
    wire new_AGEMA_signal_1965 ;
    wire new_AGEMA_signal_1966 ;
    wire new_AGEMA_signal_1967 ;
    wire new_AGEMA_signal_1968 ;
    wire new_AGEMA_signal_1969 ;
    wire new_AGEMA_signal_1970 ;
    wire new_AGEMA_signal_1971 ;
    wire new_AGEMA_signal_1972 ;
    wire new_AGEMA_signal_1973 ;
    wire new_AGEMA_signal_1974 ;
    wire new_AGEMA_signal_1975 ;
    wire new_AGEMA_signal_1976 ;
    wire new_AGEMA_signal_1977 ;
    wire new_AGEMA_signal_1978 ;
    wire new_AGEMA_signal_1979 ;
    wire new_AGEMA_signal_1980 ;
    wire new_AGEMA_signal_1981 ;
    wire new_AGEMA_signal_1982 ;
    wire new_AGEMA_signal_1983 ;
    wire new_AGEMA_signal_1984 ;
    wire new_AGEMA_signal_1985 ;
    wire new_AGEMA_signal_1986 ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1992 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1998 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2004 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2010 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2016 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2022 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2028 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2066 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2068 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2072 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2074 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2078 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2080 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2084 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2086 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2090 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2092 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2096 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2098 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2102 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2104 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2108 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2110 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2120 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2122 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2126 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2130 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2134 ;
    wire new_AGEMA_signal_2135 ;

    /* cells in depth 0 */
    xor_HPC3 #(.security_order(1), .pipeline(1)) U9 ( .a ({new_AGEMA_signal_856, roundkey[0]}), .b ({data_out_s1[60], data_out_s0[60]}), .c ({new_AGEMA_signal_858, stateXORroundkey[0]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U10 ( .a ({new_AGEMA_signal_859, roundkey[1]}), .b ({data_out_s1[61], data_out_s0[61]}), .c ({new_AGEMA_signal_861, stateXORroundkey[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U11 ( .a ({new_AGEMA_signal_862, roundkey[2]}), .b ({data_out_s1[62], data_out_s0[62]}), .c ({new_AGEMA_signal_864, stateXORroundkey[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) U12 ( .a ({new_AGEMA_signal_865, roundkey[3]}), .b ({data_out_s1[63], data_out_s0[63]}), .c ({new_AGEMA_signal_867, stateXORroundkey[3]}) ) ;
    NOR2_X1 fsm_U20 ( .A1 (reset), .A2 (fsm_n15), .ZN (fsm_n21) ) ;
    NOR2_X1 fsm_U19 ( .A1 (fsm_n14), .A2 (done), .ZN (fsm_n15) ) ;
    NOR2_X1 fsm_U18 ( .A1 (reset), .A2 (fsm_n13), .ZN (fsm_n20) ) ;
    NOR2_X1 fsm_U17 ( .A1 (fsm_ps_state_1_), .A2 (fsm_n12), .ZN (fsm_n13) ) ;
    NOR2_X1 fsm_U16 ( .A1 (fsm_n11), .A2 (fsm_n10), .ZN (fsm_n12) ) ;
    NAND2_X1 fsm_U15 ( .A1 (counter[3]), .A2 (counter[1]), .ZN (fsm_n10) ) ;
    OR2_X1 fsm_U14 ( .A1 (fsm_n9), .A2 (fsm_n8), .ZN (fsm_n11) ) ;
    NAND2_X1 fsm_U13 ( .A1 (counter[0]), .A2 (counter[4]), .ZN (fsm_n8) ) ;
    NAND2_X1 fsm_U12 ( .A1 (counter[2]), .A2 (fsm_ps_state_0_), .ZN (fsm_n9) ) ;
    NOR2_X1 fsm_U11 ( .A1 (fsm_n3), .A2 (fsm_n5), .ZN (done) ) ;
    AND2_X1 fsm_U10 ( .A1 (fsm_n14), .A2 (fsm_n5), .ZN (fsm_en_countRound) ) ;
    AND2_X1 fsm_U9 ( .A1 (fsm_countSerial[2]), .A2 (fsm_n7), .ZN (fsm_n14) ) ;
    NOR2_X1 fsm_U8 ( .A1 (fsm_n6), .A2 (fsm_n4), .ZN (fsm_n7) ) ;
    NAND2_X1 fsm_U7 ( .A1 (fsm_countSerial[1]), .A2 (fsm_countSerial[0]), .ZN (fsm_n4) ) ;
    NAND2_X1 fsm_U6 ( .A1 (fsm_n3), .A2 (fsm_countSerial[3]), .ZN (fsm_n6) ) ;
    NOR2_X1 fsm_U5 ( .A1 (fsm_ps_state_0_), .A2 (fsm_n5), .ZN (intDone) ) ;
    NOR2_X1 fsm_U4 ( .A1 (fsm_ps_state_1_), .A2 (fsm_n3), .ZN (selSbox) ) ;
    NOR2_X1 fsm_U3 ( .A1 (reset), .A2 (selSbox), .ZN (fsm_rst_countSerial) ) ;
    INV_X1 fsm_U2 ( .A (reset), .ZN (fsm_n2) ) ;
    INV_X1 fsm_U1 ( .A (fsm_rst_countSerial), .ZN (ctrlData_0_) ) ;
    NAND2_X1 fsm_cnt_rnd_U28 ( .A1 (fsm_cnt_rnd_n33), .A2 (fsm_cnt_rnd_n32), .ZN (fsm_cnt_rnd_n41) ) ;
    NAND2_X1 fsm_cnt_rnd_U27 ( .A1 (fsm_cnt_rnd_n31), .A2 (counter[1]), .ZN (fsm_cnt_rnd_n32) ) ;
    NAND2_X1 fsm_cnt_rnd_U26 ( .A1 (fsm_cnt_rnd_n30), .A2 (fsm_cnt_rnd_n24), .ZN (fsm_cnt_rnd_n33) ) ;
    NAND2_X1 fsm_cnt_rnd_U25 ( .A1 (fsm_cnt_rnd_n29), .A2 (counter[0]), .ZN (fsm_cnt_rnd_n30) ) ;
    NAND2_X1 fsm_cnt_rnd_U24 ( .A1 (fsm_cnt_rnd_n28), .A2 (fsm_cnt_rnd_n27), .ZN (fsm_cnt_rnd_n18) ) ;
    NAND2_X1 fsm_cnt_rnd_U23 ( .A1 (fsm_cnt_rnd_n26), .A2 (counter[0]), .ZN (fsm_cnt_rnd_n27) ) ;
    MUX2_X1 fsm_cnt_rnd_U22 ( .S (fsm_cnt_rnd_n5), .A (fsm_cnt_rnd_n23), .B (fsm_cnt_rnd_n22), .Z (fsm_cnt_rnd_n16) ) ;
    NAND2_X1 fsm_cnt_rnd_U21 ( .A1 (fsm_cnt_rnd_n31), .A2 (fsm_cnt_rnd_n21), .ZN (fsm_cnt_rnd_n23) ) ;
    NAND2_X1 fsm_cnt_rnd_U20 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n24), .ZN (fsm_cnt_rnd_n21) ) ;
    NOR2_X1 fsm_cnt_rnd_U19 ( .A1 (fsm_cnt_rnd_n20), .A2 (fsm_cnt_rnd_n26), .ZN (fsm_cnt_rnd_n31) ) ;
    NOR2_X1 fsm_cnt_rnd_U18 ( .A1 (fsm_en_countRound), .A2 (fsm_cnt_rnd_n6), .ZN (fsm_cnt_rnd_n26) ) ;
    INV_X1 fsm_cnt_rnd_U17 ( .A (fsm_cnt_rnd_n28), .ZN (fsm_cnt_rnd_n20) ) ;
    NAND2_X1 fsm_cnt_rnd_U16 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n3), .ZN (fsm_cnt_rnd_n28) ) ;
    MUX2_X1 fsm_cnt_rnd_U15 ( .S (counter[4]), .A (fsm_cnt_rnd_n19), .B (fsm_cnt_rnd_n17), .Z (fsm_cnt_rnd_n14) ) ;
    NAND2_X1 fsm_cnt_rnd_U14 ( .A1 (fsm_cnt_rnd_n15), .A2 (fsm_cnt_rnd_n13), .ZN (fsm_cnt_rnd_n17) ) ;
    NAND2_X1 fsm_cnt_rnd_U13 ( .A1 (fsm_cnt_rnd_n29), .A2 (fsm_cnt_rnd_n25), .ZN (fsm_cnt_rnd_n15) ) ;
    INV_X1 fsm_cnt_rnd_U12 ( .A (fsm_cnt_rnd_n12), .ZN (fsm_cnt_rnd_n29) ) ;
    NOR2_X1 fsm_cnt_rnd_U11 ( .A1 (fsm_cnt_rnd_n25), .A2 (fsm_cnt_rnd_n11), .ZN (fsm_cnt_rnd_n19) ) ;
    INV_X1 fsm_cnt_rnd_U10 ( .A (fsm_cnt_rnd_n10), .ZN (fsm_cnt_rnd_n1) ) ;
    MUX2_X1 fsm_cnt_rnd_U9 ( .S (fsm_cnt_rnd_n25), .A (fsm_cnt_rnd_n13), .B (fsm_cnt_rnd_n11), .Z (fsm_cnt_rnd_n10) ) ;
    NAND2_X1 fsm_cnt_rnd_U8 ( .A1 (counter[2]), .A2 (fsm_cnt_rnd_n22), .ZN (fsm_cnt_rnd_n11) ) ;
    NOR2_X1 fsm_cnt_rnd_U7 ( .A1 (fsm_cnt_rnd_n12), .A2 (fsm_cnt_rnd_n9), .ZN (fsm_cnt_rnd_n22) ) ;
    NAND2_X1 fsm_cnt_rnd_U6 ( .A1 (fsm_en_countRound), .A2 (fsm_n2), .ZN (fsm_cnt_rnd_n12) ) ;
    NAND2_X1 fsm_cnt_rnd_U5 ( .A1 (fsm_n2), .A2 (fsm_cnt_rnd_n8), .ZN (fsm_cnt_rnd_n13) ) ;
    NAND2_X1 fsm_cnt_rnd_U4 ( .A1 (fsm_en_countRound), .A2 (fsm_cnt_rnd_n7), .ZN (fsm_cnt_rnd_n8) ) ;
    NOR2_X1 fsm_cnt_rnd_U3 ( .A1 (fsm_cnt_rnd_n5), .A2 (fsm_cnt_rnd_n9), .ZN (fsm_cnt_rnd_n7) ) ;
    OR2_X1 fsm_cnt_rnd_U2 ( .A1 (fsm_cnt_rnd_n24), .A2 (fsm_cnt_rnd_n3), .ZN (fsm_cnt_rnd_n9) ) ;
    INV_X1 fsm_cnt_rnd_U1 ( .A (fsm_n2), .ZN (fsm_cnt_rnd_n6) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_2__U1 ( .A (counter[2]), .ZN (fsm_cnt_rnd_n5) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_0__U1 ( .A (counter[0]), .ZN (fsm_cnt_rnd_n3) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_3__U1 ( .A (counter[3]), .ZN (fsm_cnt_rnd_n25) ) ;
    INV_X1 fsm_cnt_rnd_count_reg_reg_1__U1 ( .A (fsm_cnt_rnd_n24), .ZN (counter[1]) ) ;
    NOR2_X1 fsm_cnt_ser_U12 ( .A1 (fsm_cnt_ser_n10), .A2 (fsm_cnt_ser_n9), .ZN (fsm_cnt_ser_n3) ) ;
    XNOR2_X1 fsm_cnt_ser_U11 ( .A (fsm_n3), .B (fsm_countSerial[0]), .ZN (fsm_cnt_ser_n10) ) ;
    NOR2_X1 fsm_cnt_ser_U10 ( .A1 (fsm_cnt_ser_n9), .A2 (fsm_cnt_ser_n8), .ZN (fsm_cnt_ser_n28) ) ;
    XOR2_X1 fsm_cnt_ser_U9 ( .A (fsm_countSerial[1]), .B (fsm_cnt_ser_n7), .Z (fsm_cnt_ser_n8) ) ;
    NOR2_X1 fsm_cnt_ser_U8 ( .A1 (fsm_cnt_ser_n9), .A2 (fsm_cnt_ser_n6), .ZN (fsm_cnt_ser_n26) ) ;
    XOR2_X1 fsm_cnt_ser_U7 ( .A (fsm_countSerial[3]), .B (fsm_cnt_ser_n5), .Z (fsm_cnt_ser_n6) ) ;
    NAND2_X1 fsm_cnt_ser_U6 ( .A1 (fsm_cnt_ser_n4), .A2 (fsm_countSerial[2]), .ZN (fsm_cnt_ser_n5) ) ;
    NOR2_X1 fsm_cnt_ser_U5 ( .A1 (fsm_cnt_ser_n2), .A2 (fsm_cnt_ser_n9), .ZN (fsm_cnt_ser_n1) ) ;
    INV_X1 fsm_cnt_ser_U4 ( .A (fsm_rst_countSerial), .ZN (fsm_cnt_ser_n9) ) ;
    XNOR2_X1 fsm_cnt_ser_U3 ( .A (fsm_cnt_ser_n4), .B (fsm_countSerial[2]), .ZN (fsm_cnt_ser_n2) ) ;
    NOR2_X1 fsm_cnt_ser_U2 ( .A1 (fsm_cnt_ser_n20), .A2 (fsm_cnt_ser_n7), .ZN (fsm_cnt_ser_n4) ) ;
    NAND2_X1 fsm_cnt_ser_U1 ( .A1 (fsm_n3), .A2 (fsm_countSerial[0]), .ZN (fsm_cnt_ser_n7) ) ;
    INV_X1 fsm_cnt_ser_count_reg_reg_1__U1 ( .A (fsm_countSerial[1]), .ZN (fsm_cnt_ser_n20) ) ;
    INV_X1 fsm_ps_state_reg_0__U1 ( .A (fsm_ps_state_0_), .ZN (fsm_n3) ) ;
    INV_X1 fsm_ps_state_reg_1__U1 ( .A (fsm_ps_state_1_), .ZN (fsm_n5) ) ;
    INV_X1 stateFF_state_U3 ( .A (stateFF_state_n7), .ZN (stateFF_state_n6) ) ;
    INV_X1 stateFF_state_U2 ( .A (stateFF_state_n7), .ZN (stateFF_state_n5) ) ;
    INV_X1 stateFF_state_U1 ( .A (ctrlData_0_), .ZN (stateFF_state_n7) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_2_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({data_out_s1[0], data_out_s0[0]}), .a ({new_AGEMA_signal_882, stateFF_inputPar[4]}), .c ({new_AGEMA_signal_1299, stateFF_state_gff_2_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_2_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({data_out_s1[1], data_out_s0[1]}), .a ({new_AGEMA_signal_885, stateFF_inputPar[5]}), .c ({new_AGEMA_signal_1300, stateFF_state_gff_2_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_2_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({data_out_s1[2], data_out_s0[2]}), .a ({new_AGEMA_signal_888, stateFF_inputPar[6]}), .c ({new_AGEMA_signal_1301, stateFF_state_gff_2_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_2_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({data_out_s1[3], data_out_s0[3]}), .a ({new_AGEMA_signal_891, stateFF_inputPar[7]}), .c ({new_AGEMA_signal_1302, stateFF_state_gff_2_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_3_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[4], data_out_s0[4]}), .a ({new_AGEMA_signal_894, stateFF_inputPar[8]}), .c ({new_AGEMA_signal_1318, stateFF_state_gff_3_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_3_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[5], data_out_s0[5]}), .a ({new_AGEMA_signal_897, stateFF_inputPar[9]}), .c ({new_AGEMA_signal_1319, stateFF_state_gff_3_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_3_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[6], data_out_s0[6]}), .a ({new_AGEMA_signal_900, stateFF_inputPar[10]}), .c ({new_AGEMA_signal_1320, stateFF_state_gff_3_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_3_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[7], data_out_s0[7]}), .a ({new_AGEMA_signal_903, stateFF_inputPar[11]}), .c ({new_AGEMA_signal_1321, stateFF_state_gff_3_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_4_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[8], data_out_s0[8]}), .a ({new_AGEMA_signal_906, stateFF_inputPar[12]}), .c ({new_AGEMA_signal_1322, stateFF_state_gff_4_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_4_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[9], data_out_s0[9]}), .a ({new_AGEMA_signal_909, stateFF_inputPar[13]}), .c ({new_AGEMA_signal_1323, stateFF_state_gff_4_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_4_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[10], data_out_s0[10]}), .a ({new_AGEMA_signal_912, stateFF_inputPar[14]}), .c ({new_AGEMA_signal_1324, stateFF_state_gff_4_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_4_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[11], data_out_s0[11]}), .a ({new_AGEMA_signal_914, stateFF_inputPar[15]}), .c ({new_AGEMA_signal_1325, stateFF_state_gff_4_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_5_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[12], data_out_s0[12]}), .a ({new_AGEMA_signal_917, stateFF_inputPar[16]}), .c ({new_AGEMA_signal_1326, stateFF_state_gff_5_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_5_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[13], data_out_s0[13]}), .a ({new_AGEMA_signal_920, stateFF_inputPar[17]}), .c ({new_AGEMA_signal_1327, stateFF_state_gff_5_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_5_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[14], data_out_s0[14]}), .a ({new_AGEMA_signal_923, stateFF_inputPar[18]}), .c ({new_AGEMA_signal_1328, stateFF_state_gff_5_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_5_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[15], data_out_s0[15]}), .a ({new_AGEMA_signal_926, stateFF_inputPar[19]}), .c ({new_AGEMA_signal_1329, stateFF_state_gff_5_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_6_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[16], data_out_s0[16]}), .a ({new_AGEMA_signal_929, stateFF_inputPar[20]}), .c ({new_AGEMA_signal_1330, stateFF_state_gff_6_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_6_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[17], data_out_s0[17]}), .a ({new_AGEMA_signal_932, stateFF_inputPar[21]}), .c ({new_AGEMA_signal_1331, stateFF_state_gff_6_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_6_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[18], data_out_s0[18]}), .a ({new_AGEMA_signal_935, stateFF_inputPar[22]}), .c ({new_AGEMA_signal_1332, stateFF_state_gff_6_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_6_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[19], data_out_s0[19]}), .a ({new_AGEMA_signal_938, stateFF_inputPar[23]}), .c ({new_AGEMA_signal_1333, stateFF_state_gff_6_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_7_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[20], data_out_s0[20]}), .a ({new_AGEMA_signal_941, stateFF_inputPar[24]}), .c ({new_AGEMA_signal_1334, stateFF_state_gff_7_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_7_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[21], data_out_s0[21]}), .a ({new_AGEMA_signal_944, stateFF_inputPar[25]}), .c ({new_AGEMA_signal_1335, stateFF_state_gff_7_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_7_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[22], data_out_s0[22]}), .a ({new_AGEMA_signal_947, stateFF_inputPar[26]}), .c ({new_AGEMA_signal_1336, stateFF_state_gff_7_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_7_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[23], data_out_s0[23]}), .a ({new_AGEMA_signal_950, stateFF_inputPar[27]}), .c ({new_AGEMA_signal_1337, stateFF_state_gff_7_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_8_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[24], data_out_s0[24]}), .a ({new_AGEMA_signal_953, stateFF_inputPar[28]}), .c ({new_AGEMA_signal_1338, stateFF_state_gff_8_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_8_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[25], data_out_s0[25]}), .a ({new_AGEMA_signal_956, stateFF_inputPar[29]}), .c ({new_AGEMA_signal_1339, stateFF_state_gff_8_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_8_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[26], data_out_s0[26]}), .a ({new_AGEMA_signal_959, stateFF_inputPar[30]}), .c ({new_AGEMA_signal_1340, stateFF_state_gff_8_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_8_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[27], data_out_s0[27]}), .a ({new_AGEMA_signal_961, stateFF_inputPar[31]}), .c ({new_AGEMA_signal_1341, stateFF_state_gff_8_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_9_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[28], data_out_s0[28]}), .a ({new_AGEMA_signal_964, stateFF_inputPar[32]}), .c ({new_AGEMA_signal_1342, stateFF_state_gff_9_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_9_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[29], data_out_s0[29]}), .a ({new_AGEMA_signal_967, stateFF_inputPar[33]}), .c ({new_AGEMA_signal_1343, stateFF_state_gff_9_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_9_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[30], data_out_s0[30]}), .a ({new_AGEMA_signal_970, stateFF_inputPar[34]}), .c ({new_AGEMA_signal_1344, stateFF_state_gff_9_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_9_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n6), .b ({data_out_s1[31], data_out_s0[31]}), .a ({new_AGEMA_signal_973, stateFF_inputPar[35]}), .c ({new_AGEMA_signal_1345, stateFF_state_gff_9_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_10_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[32], data_out_s0[32]}), .a ({new_AGEMA_signal_976, stateFF_inputPar[36]}), .c ({new_AGEMA_signal_1346, stateFF_state_gff_10_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_10_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[33], data_out_s0[33]}), .a ({new_AGEMA_signal_979, stateFF_inputPar[37]}), .c ({new_AGEMA_signal_1347, stateFF_state_gff_10_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_10_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[34], data_out_s0[34]}), .a ({new_AGEMA_signal_982, stateFF_inputPar[38]}), .c ({new_AGEMA_signal_1348, stateFF_state_gff_10_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_10_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[35], data_out_s0[35]}), .a ({new_AGEMA_signal_985, stateFF_inputPar[39]}), .c ({new_AGEMA_signal_1349, stateFF_state_gff_10_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_11_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[36], data_out_s0[36]}), .a ({new_AGEMA_signal_988, stateFF_inputPar[40]}), .c ({new_AGEMA_signal_1350, stateFF_state_gff_11_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_11_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[37], data_out_s0[37]}), .a ({new_AGEMA_signal_991, stateFF_inputPar[41]}), .c ({new_AGEMA_signal_1351, stateFF_state_gff_11_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_11_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[38], data_out_s0[38]}), .a ({new_AGEMA_signal_994, stateFF_inputPar[42]}), .c ({new_AGEMA_signal_1352, stateFF_state_gff_11_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_11_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[39], data_out_s0[39]}), .a ({new_AGEMA_signal_997, stateFF_inputPar[43]}), .c ({new_AGEMA_signal_1353, stateFF_state_gff_11_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_12_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[40], data_out_s0[40]}), .a ({new_AGEMA_signal_1000, stateFF_inputPar[44]}), .c ({new_AGEMA_signal_1354, stateFF_state_gff_12_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_12_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[41], data_out_s0[41]}), .a ({new_AGEMA_signal_1003, stateFF_inputPar[45]}), .c ({new_AGEMA_signal_1355, stateFF_state_gff_12_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_12_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[42], data_out_s0[42]}), .a ({new_AGEMA_signal_1006, stateFF_inputPar[46]}), .c ({new_AGEMA_signal_1356, stateFF_state_gff_12_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_12_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[43], data_out_s0[43]}), .a ({new_AGEMA_signal_1008, stateFF_inputPar[47]}), .c ({new_AGEMA_signal_1357, stateFF_state_gff_12_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_13_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[44], data_out_s0[44]}), .a ({new_AGEMA_signal_1011, stateFF_inputPar[48]}), .c ({new_AGEMA_signal_1358, stateFF_state_gff_13_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_13_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[45], data_out_s0[45]}), .a ({new_AGEMA_signal_1014, stateFF_inputPar[49]}), .c ({new_AGEMA_signal_1359, stateFF_state_gff_13_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_13_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[46], data_out_s0[46]}), .a ({new_AGEMA_signal_1017, stateFF_inputPar[50]}), .c ({new_AGEMA_signal_1360, stateFF_state_gff_13_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_13_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[47], data_out_s0[47]}), .a ({new_AGEMA_signal_1020, stateFF_inputPar[51]}), .c ({new_AGEMA_signal_1361, stateFF_state_gff_13_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_14_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[48], data_out_s0[48]}), .a ({new_AGEMA_signal_1023, stateFF_inputPar[52]}), .c ({new_AGEMA_signal_1362, stateFF_state_gff_14_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_14_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[49], data_out_s0[49]}), .a ({new_AGEMA_signal_1026, stateFF_inputPar[53]}), .c ({new_AGEMA_signal_1363, stateFF_state_gff_14_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_14_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[50], data_out_s0[50]}), .a ({new_AGEMA_signal_1029, stateFF_inputPar[54]}), .c ({new_AGEMA_signal_1364, stateFF_state_gff_14_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_14_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[51], data_out_s0[51]}), .a ({new_AGEMA_signal_1032, stateFF_inputPar[55]}), .c ({new_AGEMA_signal_1365, stateFF_state_gff_14_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_15_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[52], data_out_s0[52]}), .a ({new_AGEMA_signal_1035, stateFF_inputPar[56]}), .c ({new_AGEMA_signal_1366, stateFF_state_gff_15_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_15_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[53], data_out_s0[53]}), .a ({new_AGEMA_signal_1038, stateFF_inputPar[57]}), .c ({new_AGEMA_signal_1367, stateFF_state_gff_15_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_15_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[54], data_out_s0[54]}), .a ({new_AGEMA_signal_1041, stateFF_inputPar[58]}), .c ({new_AGEMA_signal_1368, stateFF_state_gff_15_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_15_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[55], data_out_s0[55]}), .a ({new_AGEMA_signal_1044, stateFF_inputPar[59]}), .c ({new_AGEMA_signal_1369, stateFF_state_gff_15_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_16_MUX_inst1_mux_inst_0_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[56], data_out_s0[56]}), .a ({new_AGEMA_signal_1047, stateFF_inputPar[60]}), .c ({new_AGEMA_signal_1370, stateFF_state_gff_16_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_16_MUX_inst1_mux_inst_1_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[57], data_out_s0[57]}), .a ({new_AGEMA_signal_1050, stateFF_inputPar[61]}), .c ({new_AGEMA_signal_1371, stateFF_state_gff_16_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_16_MUX_inst1_mux_inst_2_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[58], data_out_s0[58]}), .a ({new_AGEMA_signal_1053, stateFF_inputPar[62]}), .c ({new_AGEMA_signal_1372, stateFF_state_gff_16_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_16_MUX_inst1_mux_inst_3_U1 ( .s (stateFF_state_n5), .b ({data_out_s1[59], data_out_s0[59]}), .a ({new_AGEMA_signal_1055, stateFF_inputPar[63]}), .c ({new_AGEMA_signal_1373, stateFF_state_gff_16_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_0_U1 ( .s (reset), .b ({data_out_s1[0], data_out_s0[0]}), .a ({data_in_s1[0], data_in_s0[0]}), .c ({new_AGEMA_signal_870, stateFF_inputPar[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_1_U1 ( .s (reset), .b ({data_out_s1[4], data_out_s0[4]}), .a ({data_in_s1[1], data_in_s0[1]}), .c ({new_AGEMA_signal_873, stateFF_inputPar[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_2_U1 ( .s (reset), .b ({data_out_s1[8], data_out_s0[8]}), .a ({data_in_s1[2], data_in_s0[2]}), .c ({new_AGEMA_signal_876, stateFF_inputPar[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_3_U1 ( .s (reset), .b ({data_out_s1[12], data_out_s0[12]}), .a ({data_in_s1[3], data_in_s0[3]}), .c ({new_AGEMA_signal_879, stateFF_inputPar[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_4_U1 ( .s (reset), .b ({data_out_s1[16], data_out_s0[16]}), .a ({data_in_s1[4], data_in_s0[4]}), .c ({new_AGEMA_signal_882, stateFF_inputPar[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_5_U1 ( .s (reset), .b ({data_out_s1[20], data_out_s0[20]}), .a ({data_in_s1[5], data_in_s0[5]}), .c ({new_AGEMA_signal_885, stateFF_inputPar[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_6_U1 ( .s (reset), .b ({data_out_s1[24], data_out_s0[24]}), .a ({data_in_s1[6], data_in_s0[6]}), .c ({new_AGEMA_signal_888, stateFF_inputPar[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_7_U1 ( .s (reset), .b ({data_out_s1[28], data_out_s0[28]}), .a ({data_in_s1[7], data_in_s0[7]}), .c ({new_AGEMA_signal_891, stateFF_inputPar[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_8_U1 ( .s (reset), .b ({data_out_s1[32], data_out_s0[32]}), .a ({data_in_s1[8], data_in_s0[8]}), .c ({new_AGEMA_signal_894, stateFF_inputPar[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_9_U1 ( .s (reset), .b ({data_out_s1[36], data_out_s0[36]}), .a ({data_in_s1[9], data_in_s0[9]}), .c ({new_AGEMA_signal_897, stateFF_inputPar[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_10_U1 ( .s (reset), .b ({data_out_s1[40], data_out_s0[40]}), .a ({data_in_s1[10], data_in_s0[10]}), .c ({new_AGEMA_signal_900, stateFF_inputPar[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_11_U1 ( .s (reset), .b ({data_out_s1[44], data_out_s0[44]}), .a ({data_in_s1[11], data_in_s0[11]}), .c ({new_AGEMA_signal_903, stateFF_inputPar[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_12_U1 ( .s (reset), .b ({data_out_s1[48], data_out_s0[48]}), .a ({data_in_s1[12], data_in_s0[12]}), .c ({new_AGEMA_signal_906, stateFF_inputPar[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_13_U1 ( .s (reset), .b ({data_out_s1[52], data_out_s0[52]}), .a ({data_in_s1[13], data_in_s0[13]}), .c ({new_AGEMA_signal_909, stateFF_inputPar[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_14_U1 ( .s (reset), .b ({data_out_s1[56], data_out_s0[56]}), .a ({data_in_s1[14], data_in_s0[14]}), .c ({new_AGEMA_signal_912, stateFF_inputPar[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_15_U1 ( .s (reset), .b ({data_out_s1[60], data_out_s0[60]}), .a ({data_in_s1[15], data_in_s0[15]}), .c ({new_AGEMA_signal_914, stateFF_inputPar[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_16_U1 ( .s (reset), .b ({data_out_s1[1], data_out_s0[1]}), .a ({data_in_s1[16], data_in_s0[16]}), .c ({new_AGEMA_signal_917, stateFF_inputPar[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_17_U1 ( .s (reset), .b ({data_out_s1[5], data_out_s0[5]}), .a ({data_in_s1[17], data_in_s0[17]}), .c ({new_AGEMA_signal_920, stateFF_inputPar[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_18_U1 ( .s (reset), .b ({data_out_s1[9], data_out_s0[9]}), .a ({data_in_s1[18], data_in_s0[18]}), .c ({new_AGEMA_signal_923, stateFF_inputPar[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_19_U1 ( .s (reset), .b ({data_out_s1[13], data_out_s0[13]}), .a ({data_in_s1[19], data_in_s0[19]}), .c ({new_AGEMA_signal_926, stateFF_inputPar[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_20_U1 ( .s (reset), .b ({data_out_s1[17], data_out_s0[17]}), .a ({data_in_s1[20], data_in_s0[20]}), .c ({new_AGEMA_signal_929, stateFF_inputPar[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_21_U1 ( .s (reset), .b ({data_out_s1[21], data_out_s0[21]}), .a ({data_in_s1[21], data_in_s0[21]}), .c ({new_AGEMA_signal_932, stateFF_inputPar[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_22_U1 ( .s (reset), .b ({data_out_s1[25], data_out_s0[25]}), .a ({data_in_s1[22], data_in_s0[22]}), .c ({new_AGEMA_signal_935, stateFF_inputPar[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_23_U1 ( .s (reset), .b ({data_out_s1[29], data_out_s0[29]}), .a ({data_in_s1[23], data_in_s0[23]}), .c ({new_AGEMA_signal_938, stateFF_inputPar[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_24_U1 ( .s (reset), .b ({data_out_s1[33], data_out_s0[33]}), .a ({data_in_s1[24], data_in_s0[24]}), .c ({new_AGEMA_signal_941, stateFF_inputPar[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_25_U1 ( .s (reset), .b ({data_out_s1[37], data_out_s0[37]}), .a ({data_in_s1[25], data_in_s0[25]}), .c ({new_AGEMA_signal_944, stateFF_inputPar[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_26_U1 ( .s (reset), .b ({data_out_s1[41], data_out_s0[41]}), .a ({data_in_s1[26], data_in_s0[26]}), .c ({new_AGEMA_signal_947, stateFF_inputPar[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_27_U1 ( .s (reset), .b ({data_out_s1[45], data_out_s0[45]}), .a ({data_in_s1[27], data_in_s0[27]}), .c ({new_AGEMA_signal_950, stateFF_inputPar[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_28_U1 ( .s (reset), .b ({data_out_s1[49], data_out_s0[49]}), .a ({data_in_s1[28], data_in_s0[28]}), .c ({new_AGEMA_signal_953, stateFF_inputPar[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_29_U1 ( .s (reset), .b ({data_out_s1[53], data_out_s0[53]}), .a ({data_in_s1[29], data_in_s0[29]}), .c ({new_AGEMA_signal_956, stateFF_inputPar[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_30_U1 ( .s (reset), .b ({data_out_s1[57], data_out_s0[57]}), .a ({data_in_s1[30], data_in_s0[30]}), .c ({new_AGEMA_signal_959, stateFF_inputPar[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_31_U1 ( .s (reset), .b ({data_out_s1[61], data_out_s0[61]}), .a ({data_in_s1[31], data_in_s0[31]}), .c ({new_AGEMA_signal_961, stateFF_inputPar[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_32_U1 ( .s (reset), .b ({data_out_s1[2], data_out_s0[2]}), .a ({data_in_s1[32], data_in_s0[32]}), .c ({new_AGEMA_signal_964, stateFF_inputPar[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_33_U1 ( .s (reset), .b ({data_out_s1[6], data_out_s0[6]}), .a ({data_in_s1[33], data_in_s0[33]}), .c ({new_AGEMA_signal_967, stateFF_inputPar[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_34_U1 ( .s (reset), .b ({data_out_s1[10], data_out_s0[10]}), .a ({data_in_s1[34], data_in_s0[34]}), .c ({new_AGEMA_signal_970, stateFF_inputPar[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_35_U1 ( .s (reset), .b ({data_out_s1[14], data_out_s0[14]}), .a ({data_in_s1[35], data_in_s0[35]}), .c ({new_AGEMA_signal_973, stateFF_inputPar[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_36_U1 ( .s (reset), .b ({data_out_s1[18], data_out_s0[18]}), .a ({data_in_s1[36], data_in_s0[36]}), .c ({new_AGEMA_signal_976, stateFF_inputPar[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_37_U1 ( .s (reset), .b ({data_out_s1[22], data_out_s0[22]}), .a ({data_in_s1[37], data_in_s0[37]}), .c ({new_AGEMA_signal_979, stateFF_inputPar[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_38_U1 ( .s (reset), .b ({data_out_s1[26], data_out_s0[26]}), .a ({data_in_s1[38], data_in_s0[38]}), .c ({new_AGEMA_signal_982, stateFF_inputPar[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_39_U1 ( .s (reset), .b ({data_out_s1[30], data_out_s0[30]}), .a ({data_in_s1[39], data_in_s0[39]}), .c ({new_AGEMA_signal_985, stateFF_inputPar[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_40_U1 ( .s (reset), .b ({data_out_s1[34], data_out_s0[34]}), .a ({data_in_s1[40], data_in_s0[40]}), .c ({new_AGEMA_signal_988, stateFF_inputPar[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_41_U1 ( .s (reset), .b ({data_out_s1[38], data_out_s0[38]}), .a ({data_in_s1[41], data_in_s0[41]}), .c ({new_AGEMA_signal_991, stateFF_inputPar[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_42_U1 ( .s (reset), .b ({data_out_s1[42], data_out_s0[42]}), .a ({data_in_s1[42], data_in_s0[42]}), .c ({new_AGEMA_signal_994, stateFF_inputPar[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_43_U1 ( .s (reset), .b ({data_out_s1[46], data_out_s0[46]}), .a ({data_in_s1[43], data_in_s0[43]}), .c ({new_AGEMA_signal_997, stateFF_inputPar[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_44_U1 ( .s (reset), .b ({data_out_s1[50], data_out_s0[50]}), .a ({data_in_s1[44], data_in_s0[44]}), .c ({new_AGEMA_signal_1000, stateFF_inputPar[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_45_U1 ( .s (reset), .b ({data_out_s1[54], data_out_s0[54]}), .a ({data_in_s1[45], data_in_s0[45]}), .c ({new_AGEMA_signal_1003, stateFF_inputPar[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_46_U1 ( .s (reset), .b ({data_out_s1[58], data_out_s0[58]}), .a ({data_in_s1[46], data_in_s0[46]}), .c ({new_AGEMA_signal_1006, stateFF_inputPar[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_47_U1 ( .s (reset), .b ({data_out_s1[62], data_out_s0[62]}), .a ({data_in_s1[47], data_in_s0[47]}), .c ({new_AGEMA_signal_1008, stateFF_inputPar[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_48_U1 ( .s (reset), .b ({data_out_s1[3], data_out_s0[3]}), .a ({data_in_s1[48], data_in_s0[48]}), .c ({new_AGEMA_signal_1011, stateFF_inputPar[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_49_U1 ( .s (reset), .b ({data_out_s1[7], data_out_s0[7]}), .a ({data_in_s1[49], data_in_s0[49]}), .c ({new_AGEMA_signal_1014, stateFF_inputPar[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_50_U1 ( .s (reset), .b ({data_out_s1[11], data_out_s0[11]}), .a ({data_in_s1[50], data_in_s0[50]}), .c ({new_AGEMA_signal_1017, stateFF_inputPar[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_51_U1 ( .s (reset), .b ({data_out_s1[15], data_out_s0[15]}), .a ({data_in_s1[51], data_in_s0[51]}), .c ({new_AGEMA_signal_1020, stateFF_inputPar[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_52_U1 ( .s (reset), .b ({data_out_s1[19], data_out_s0[19]}), .a ({data_in_s1[52], data_in_s0[52]}), .c ({new_AGEMA_signal_1023, stateFF_inputPar[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_53_U1 ( .s (reset), .b ({data_out_s1[23], data_out_s0[23]}), .a ({data_in_s1[53], data_in_s0[53]}), .c ({new_AGEMA_signal_1026, stateFF_inputPar[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_54_U1 ( .s (reset), .b ({data_out_s1[27], data_out_s0[27]}), .a ({data_in_s1[54], data_in_s0[54]}), .c ({new_AGEMA_signal_1029, stateFF_inputPar[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_55_U1 ( .s (reset), .b ({data_out_s1[31], data_out_s0[31]}), .a ({data_in_s1[55], data_in_s0[55]}), .c ({new_AGEMA_signal_1032, stateFF_inputPar[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_56_U1 ( .s (reset), .b ({data_out_s1[35], data_out_s0[35]}), .a ({data_in_s1[56], data_in_s0[56]}), .c ({new_AGEMA_signal_1035, stateFF_inputPar[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_57_U1 ( .s (reset), .b ({data_out_s1[39], data_out_s0[39]}), .a ({data_in_s1[57], data_in_s0[57]}), .c ({new_AGEMA_signal_1038, stateFF_inputPar[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_58_U1 ( .s (reset), .b ({data_out_s1[43], data_out_s0[43]}), .a ({data_in_s1[58], data_in_s0[58]}), .c ({new_AGEMA_signal_1041, stateFF_inputPar[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_59_U1 ( .s (reset), .b ({data_out_s1[47], data_out_s0[47]}), .a ({data_in_s1[59], data_in_s0[59]}), .c ({new_AGEMA_signal_1044, stateFF_inputPar[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_60_U1 ( .s (reset), .b ({data_out_s1[51], data_out_s0[51]}), .a ({data_in_s1[60], data_in_s0[60]}), .c ({new_AGEMA_signal_1047, stateFF_inputPar[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_61_U1 ( .s (reset), .b ({data_out_s1[55], data_out_s0[55]}), .a ({data_in_s1[61], data_in_s0[61]}), .c ({new_AGEMA_signal_1050, stateFF_inputPar[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_62_U1 ( .s (reset), .b ({data_out_s1[59], data_out_s0[59]}), .a ({data_in_s1[62], data_in_s0[62]}), .c ({new_AGEMA_signal_1053, stateFF_inputPar[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_MUX_inputPar_mux_inst_63_U1 ( .s (reset), .b ({data_out_s1[63], data_out_s0[63]}), .a ({data_in_s1[63], data_in_s0[63]}), .c ({new_AGEMA_signal_1055, stateFF_inputPar[63]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) keyFF_U5 ( .a ({1'b0, counter[4]}), .b ({new_AGEMA_signal_1056, keyFF_outputPar[22]}), .c ({new_AGEMA_signal_1057, keyFF_counterAdd[4]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) keyFF_U4 ( .a ({1'b0, counter[3]}), .b ({new_AGEMA_signal_1058, keyFF_outputPar[21]}), .c ({new_AGEMA_signal_1059, keyFF_counterAdd[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) keyFF_U3 ( .a ({1'b0, counter[2]}), .b ({new_AGEMA_signal_1060, keyFF_outputPar[20]}), .c ({new_AGEMA_signal_1061, keyFF_counterAdd[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) keyFF_U2 ( .a ({1'b0, counter[1]}), .b ({new_AGEMA_signal_1274, keyFF_outputPar[19]}), .c ({new_AGEMA_signal_1275, keyFF_counterAdd[1]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) keyFF_U1 ( .a ({1'b0, counter[0]}), .b ({new_AGEMA_signal_1062, keyFF_outputPar[18]}), .c ({new_AGEMA_signal_1063, keyFF_counterAdd[0]}) ) ;
    INV_X1 keyFF_keystate_U3 ( .A (keyFF_keystate_n8), .ZN (keyFF_keystate_n6) ) ;
    INV_X1 keyFF_keystate_U2 ( .A (keyFF_keystate_n8), .ZN (keyFF_keystate_n7) ) ;
    INV_X1 keyFF_keystate_U1 ( .A (ctrlData_0_), .ZN (keyFF_keystate_n8) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_856, roundkey[0]}), .a ({new_AGEMA_signal_1066, keyFF_inputPar[0]}), .c ({new_AGEMA_signal_1374, keyFF_keystate_gff_1_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_859, roundkey[1]}), .a ({new_AGEMA_signal_1069, keyFF_inputPar[1]}), .c ({new_AGEMA_signal_1375, keyFF_keystate_gff_1_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_862, roundkey[2]}), .a ({new_AGEMA_signal_1072, keyFF_inputPar[2]}), .c ({new_AGEMA_signal_1376, keyFF_keystate_gff_1_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_1_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_865, roundkey[3]}), .a ({new_AGEMA_signal_1075, keyFF_inputPar[3]}), .c ({new_AGEMA_signal_1377, keyFF_keystate_gff_1_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1287, keyRegKS[1]}), .a ({new_AGEMA_signal_1078, keyFF_inputPar[4]}), .c ({new_AGEMA_signal_1378, keyFF_keystate_gff_2_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1289, keyRegKS[2]}), .a ({new_AGEMA_signal_1081, keyFF_inputPar[5]}), .c ({new_AGEMA_signal_1379, keyFF_keystate_gff_2_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1291, keyRegKS[3]}), .a ({new_AGEMA_signal_1084, keyFF_inputPar[6]}), .c ({new_AGEMA_signal_1380, keyFF_keystate_gff_2_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_2_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1064, keyFF_outputPar[3]}), .a ({new_AGEMA_signal_1087, keyFF_inputPar[7]}), .c ({new_AGEMA_signal_1381, keyFF_keystate_gff_2_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1067, keyFF_outputPar[4]}), .a ({new_AGEMA_signal_1090, keyFF_inputPar[8]}), .c ({new_AGEMA_signal_1382, keyFF_keystate_gff_3_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1070, keyFF_outputPar[5]}), .a ({new_AGEMA_signal_1093, keyFF_inputPar[9]}), .c ({new_AGEMA_signal_1383, keyFF_keystate_gff_3_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1073, keyFF_outputPar[6]}), .a ({new_AGEMA_signal_1096, keyFF_inputPar[10]}), .c ({new_AGEMA_signal_1384, keyFF_keystate_gff_3_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_3_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1076, keyFF_outputPar[7]}), .a ({new_AGEMA_signal_1099, keyFF_inputPar[11]}), .c ({new_AGEMA_signal_1385, keyFF_keystate_gff_3_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1079, keyFF_outputPar[8]}), .a ({new_AGEMA_signal_1102, keyFF_inputPar[12]}), .c ({new_AGEMA_signal_1386, keyFF_keystate_gff_4_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1082, keyFF_outputPar[9]}), .a ({new_AGEMA_signal_1105, keyFF_inputPar[13]}), .c ({new_AGEMA_signal_1387, keyFF_keystate_gff_4_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1085, keyFF_outputPar[10]}), .a ({new_AGEMA_signal_1108, keyFF_inputPar[14]}), .c ({new_AGEMA_signal_1388, keyFF_keystate_gff_4_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_4_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1088, keyFF_outputPar[11]}), .a ({new_AGEMA_signal_1277, keyFF_inputPar[15]}), .c ({new_AGEMA_signal_1389, keyFF_keystate_gff_4_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1091, keyFF_outputPar[12]}), .a ({new_AGEMA_signal_1285, keyFF_inputPar[16]}), .c ({new_AGEMA_signal_1303, keyFF_keystate_gff_5_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1094, keyFF_outputPar[13]}), .a ({new_AGEMA_signal_1279, keyFF_inputPar[17]}), .c ({new_AGEMA_signal_1304, keyFF_keystate_gff_5_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1097, keyFF_outputPar[14]}), .a ({new_AGEMA_signal_1281, keyFF_inputPar[18]}), .c ({new_AGEMA_signal_1305, keyFF_keystate_gff_5_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_5_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1100, keyFF_outputPar[15]}), .a ({new_AGEMA_signal_1283, keyFF_inputPar[19]}), .c ({new_AGEMA_signal_1306, keyFF_keystate_gff_5_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_0_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1103, keyFF_outputPar[16]}), .a ({new_AGEMA_signal_1111, keyFF_inputPar[20]}), .c ({new_AGEMA_signal_1307, keyFF_keystate_gff_6_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_1_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1106, keyFF_outputPar[17]}), .a ({new_AGEMA_signal_1114, keyFF_inputPar[21]}), .c ({new_AGEMA_signal_1308, keyFF_keystate_gff_6_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_2_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1062, keyFF_outputPar[18]}), .a ({new_AGEMA_signal_1117, keyFF_inputPar[22]}), .c ({new_AGEMA_signal_1309, keyFF_keystate_gff_6_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_6_MUX_inst1_mux_inst_3_U1 ( .s (ctrlData_0_), .b ({new_AGEMA_signal_1274, keyFF_outputPar[19]}), .a ({new_AGEMA_signal_1120, keyFF_inputPar[23]}), .c ({new_AGEMA_signal_1310, keyFF_keystate_gff_6_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1060, keyFF_outputPar[20]}), .a ({new_AGEMA_signal_1123, keyFF_inputPar[24]}), .c ({new_AGEMA_signal_1390, keyFF_keystate_gff_7_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1058, keyFF_outputPar[21]}), .a ({new_AGEMA_signal_1126, keyFF_inputPar[25]}), .c ({new_AGEMA_signal_1391, keyFF_keystate_gff_7_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1056, keyFF_outputPar[22]}), .a ({new_AGEMA_signal_1129, keyFF_inputPar[26]}), .c ({new_AGEMA_signal_1392, keyFF_keystate_gff_7_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_7_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1109, keyFF_outputPar[23]}), .a ({new_AGEMA_signal_1132, keyFF_inputPar[27]}), .c ({new_AGEMA_signal_1393, keyFF_keystate_gff_7_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1112, keyFF_outputPar[24]}), .a ({new_AGEMA_signal_1135, keyFF_inputPar[28]}), .c ({new_AGEMA_signal_1394, keyFF_keystate_gff_8_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1115, keyFF_outputPar[25]}), .a ({new_AGEMA_signal_1138, keyFF_inputPar[29]}), .c ({new_AGEMA_signal_1395, keyFF_keystate_gff_8_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1118, keyFF_outputPar[26]}), .a ({new_AGEMA_signal_1141, keyFF_inputPar[30]}), .c ({new_AGEMA_signal_1396, keyFF_keystate_gff_8_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_8_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1121, keyFF_outputPar[27]}), .a ({new_AGEMA_signal_1144, keyFF_inputPar[31]}), .c ({new_AGEMA_signal_1397, keyFF_keystate_gff_8_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1124, keyFF_outputPar[28]}), .a ({new_AGEMA_signal_1147, keyFF_inputPar[32]}), .c ({new_AGEMA_signal_1398, keyFF_keystate_gff_9_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1127, keyFF_outputPar[29]}), .a ({new_AGEMA_signal_1150, keyFF_inputPar[33]}), .c ({new_AGEMA_signal_1399, keyFF_keystate_gff_9_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1130, keyFF_outputPar[30]}), .a ({new_AGEMA_signal_1153, keyFF_inputPar[34]}), .c ({new_AGEMA_signal_1400, keyFF_keystate_gff_9_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_9_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1133, keyFF_outputPar[31]}), .a ({new_AGEMA_signal_1156, keyFF_inputPar[35]}), .c ({new_AGEMA_signal_1401, keyFF_keystate_gff_9_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1136, keyFF_outputPar[32]}), .a ({new_AGEMA_signal_1159, keyFF_inputPar[36]}), .c ({new_AGEMA_signal_1402, keyFF_keystate_gff_10_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1139, keyFF_outputPar[33]}), .a ({new_AGEMA_signal_1162, keyFF_inputPar[37]}), .c ({new_AGEMA_signal_1403, keyFF_keystate_gff_10_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1142, keyFF_outputPar[34]}), .a ({new_AGEMA_signal_1165, keyFF_inputPar[38]}), .c ({new_AGEMA_signal_1404, keyFF_keystate_gff_10_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_10_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1145, keyFF_outputPar[35]}), .a ({new_AGEMA_signal_1168, keyFF_inputPar[39]}), .c ({new_AGEMA_signal_1405, keyFF_keystate_gff_10_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1148, keyFF_outputPar[36]}), .a ({new_AGEMA_signal_1171, keyFF_inputPar[40]}), .c ({new_AGEMA_signal_1406, keyFF_keystate_gff_11_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1151, keyFF_outputPar[37]}), .a ({new_AGEMA_signal_1174, keyFF_inputPar[41]}), .c ({new_AGEMA_signal_1407, keyFF_keystate_gff_11_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1154, keyFF_outputPar[38]}), .a ({new_AGEMA_signal_1177, keyFF_inputPar[42]}), .c ({new_AGEMA_signal_1408, keyFF_keystate_gff_11_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_11_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1157, keyFF_outputPar[39]}), .a ({new_AGEMA_signal_1180, keyFF_inputPar[43]}), .c ({new_AGEMA_signal_1409, keyFF_keystate_gff_11_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1160, keyFF_outputPar[40]}), .a ({new_AGEMA_signal_1183, keyFF_inputPar[44]}), .c ({new_AGEMA_signal_1410, keyFF_keystate_gff_12_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1163, keyFF_outputPar[41]}), .a ({new_AGEMA_signal_1186, keyFF_inputPar[45]}), .c ({new_AGEMA_signal_1411, keyFF_keystate_gff_12_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1166, keyFF_outputPar[42]}), .a ({new_AGEMA_signal_1189, keyFF_inputPar[46]}), .c ({new_AGEMA_signal_1412, keyFF_keystate_gff_12_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_12_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1169, keyFF_outputPar[43]}), .a ({new_AGEMA_signal_1192, keyFF_inputPar[47]}), .c ({new_AGEMA_signal_1413, keyFF_keystate_gff_12_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1172, keyFF_outputPar[44]}), .a ({new_AGEMA_signal_1195, keyFF_inputPar[48]}), .c ({new_AGEMA_signal_1414, keyFF_keystate_gff_13_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1175, keyFF_outputPar[45]}), .a ({new_AGEMA_signal_1198, keyFF_inputPar[49]}), .c ({new_AGEMA_signal_1415, keyFF_keystate_gff_13_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1178, keyFF_outputPar[46]}), .a ({new_AGEMA_signal_1201, keyFF_inputPar[50]}), .c ({new_AGEMA_signal_1416, keyFF_keystate_gff_13_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_13_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n7), .b ({new_AGEMA_signal_1181, keyFF_outputPar[47]}), .a ({new_AGEMA_signal_1204, keyFF_inputPar[51]}), .c ({new_AGEMA_signal_1417, keyFF_keystate_gff_13_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1184, keyFF_outputPar[48]}), .a ({new_AGEMA_signal_1207, keyFF_inputPar[52]}), .c ({new_AGEMA_signal_1418, keyFF_keystate_gff_14_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1187, keyFF_outputPar[49]}), .a ({new_AGEMA_signal_1210, keyFF_inputPar[53]}), .c ({new_AGEMA_signal_1419, keyFF_keystate_gff_14_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1190, keyFF_outputPar[50]}), .a ({new_AGEMA_signal_1213, keyFF_inputPar[54]}), .c ({new_AGEMA_signal_1420, keyFF_keystate_gff_14_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_14_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1193, keyFF_outputPar[51]}), .a ({new_AGEMA_signal_1216, keyFF_inputPar[55]}), .c ({new_AGEMA_signal_1421, keyFF_keystate_gff_14_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1196, keyFF_outputPar[52]}), .a ({new_AGEMA_signal_1219, keyFF_inputPar[56]}), .c ({new_AGEMA_signal_1422, keyFF_keystate_gff_15_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1199, keyFF_outputPar[53]}), .a ({new_AGEMA_signal_1222, keyFF_inputPar[57]}), .c ({new_AGEMA_signal_1423, keyFF_keystate_gff_15_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1202, keyFF_outputPar[54]}), .a ({new_AGEMA_signal_1225, keyFF_inputPar[58]}), .c ({new_AGEMA_signal_1424, keyFF_keystate_gff_15_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_15_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1205, keyFF_outputPar[55]}), .a ({new_AGEMA_signal_1228, keyFF_inputPar[59]}), .c ({new_AGEMA_signal_1425, keyFF_keystate_gff_15_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1208, keyFF_outputPar[56]}), .a ({new_AGEMA_signal_1231, keyFF_inputPar[60]}), .c ({new_AGEMA_signal_1426, keyFF_keystate_gff_16_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1211, keyFF_outputPar[57]}), .a ({new_AGEMA_signal_1234, keyFF_inputPar[61]}), .c ({new_AGEMA_signal_1427, keyFF_keystate_gff_16_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1214, keyFF_outputPar[58]}), .a ({new_AGEMA_signal_1237, keyFF_inputPar[62]}), .c ({new_AGEMA_signal_1428, keyFF_keystate_gff_16_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_16_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1217, keyFF_outputPar[59]}), .a ({new_AGEMA_signal_1240, keyFF_inputPar[63]}), .c ({new_AGEMA_signal_1429, keyFF_keystate_gff_16_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1220, keyFF_outputPar[60]}), .a ({new_AGEMA_signal_1243, keyFF_inputPar[64]}), .c ({new_AGEMA_signal_1430, keyFF_keystate_gff_17_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1223, keyFF_outputPar[61]}), .a ({new_AGEMA_signal_1246, keyFF_inputPar[65]}), .c ({new_AGEMA_signal_1431, keyFF_keystate_gff_17_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1226, keyFF_outputPar[62]}), .a ({new_AGEMA_signal_1249, keyFF_inputPar[66]}), .c ({new_AGEMA_signal_1432, keyFF_keystate_gff_17_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_17_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1229, keyFF_outputPar[63]}), .a ({new_AGEMA_signal_1252, keyFF_inputPar[67]}), .c ({new_AGEMA_signal_1433, keyFF_keystate_gff_17_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1232, keyFF_outputPar[64]}), .a ({new_AGEMA_signal_1255, keyFF_inputPar[68]}), .c ({new_AGEMA_signal_1434, keyFF_keystate_gff_18_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1235, keyFF_outputPar[65]}), .a ({new_AGEMA_signal_1258, keyFF_inputPar[69]}), .c ({new_AGEMA_signal_1435, keyFF_keystate_gff_18_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1238, keyFF_outputPar[66]}), .a ({new_AGEMA_signal_1261, keyFF_inputPar[70]}), .c ({new_AGEMA_signal_1436, keyFF_keystate_gff_18_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_18_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1241, keyFF_outputPar[67]}), .a ({new_AGEMA_signal_1264, keyFF_inputPar[71]}), .c ({new_AGEMA_signal_1437, keyFF_keystate_gff_18_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_0_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1244, keyFF_outputPar[68]}), .a ({new_AGEMA_signal_1267, keyFF_inputPar[72]}), .c ({new_AGEMA_signal_1438, keyFF_keystate_gff_19_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_1_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1247, keyFF_outputPar[69]}), .a ({new_AGEMA_signal_1269, keyFF_inputPar[73]}), .c ({new_AGEMA_signal_1439, keyFF_keystate_gff_19_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_2_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1250, keyFF_outputPar[70]}), .a ({new_AGEMA_signal_1271, keyFF_inputPar[74]}), .c ({new_AGEMA_signal_1440, keyFF_keystate_gff_19_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_19_MUX_inst1_mux_inst_3_U1 ( .s (keyFF_keystate_n6), .b ({new_AGEMA_signal_1253, keyFF_outputPar[71]}), .a ({new_AGEMA_signal_1273, keyFF_inputPar[75]}), .c ({new_AGEMA_signal_1441, keyFF_keystate_gff_19_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_0_U1 ( .s (reset), .b ({new_AGEMA_signal_1064, keyFF_outputPar[3]}), .a ({key_s1[0], key_s0[0]}), .c ({new_AGEMA_signal_1066, keyFF_inputPar[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_1_U1 ( .s (reset), .b ({new_AGEMA_signal_1067, keyFF_outputPar[4]}), .a ({key_s1[1], key_s0[1]}), .c ({new_AGEMA_signal_1069, keyFF_inputPar[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_2_U1 ( .s (reset), .b ({new_AGEMA_signal_1070, keyFF_outputPar[5]}), .a ({key_s1[2], key_s0[2]}), .c ({new_AGEMA_signal_1072, keyFF_inputPar[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_3_U1 ( .s (reset), .b ({new_AGEMA_signal_1073, keyFF_outputPar[6]}), .a ({key_s1[3], key_s0[3]}), .c ({new_AGEMA_signal_1075, keyFF_inputPar[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_4_U1 ( .s (reset), .b ({new_AGEMA_signal_1076, keyFF_outputPar[7]}), .a ({key_s1[4], key_s0[4]}), .c ({new_AGEMA_signal_1078, keyFF_inputPar[4]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_5_U1 ( .s (reset), .b ({new_AGEMA_signal_1079, keyFF_outputPar[8]}), .a ({key_s1[5], key_s0[5]}), .c ({new_AGEMA_signal_1081, keyFF_inputPar[5]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_6_U1 ( .s (reset), .b ({new_AGEMA_signal_1082, keyFF_outputPar[9]}), .a ({key_s1[6], key_s0[6]}), .c ({new_AGEMA_signal_1084, keyFF_inputPar[6]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_7_U1 ( .s (reset), .b ({new_AGEMA_signal_1085, keyFF_outputPar[10]}), .a ({key_s1[7], key_s0[7]}), .c ({new_AGEMA_signal_1087, keyFF_inputPar[7]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_8_U1 ( .s (reset), .b ({new_AGEMA_signal_1088, keyFF_outputPar[11]}), .a ({key_s1[8], key_s0[8]}), .c ({new_AGEMA_signal_1090, keyFF_inputPar[8]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_9_U1 ( .s (reset), .b ({new_AGEMA_signal_1091, keyFF_outputPar[12]}), .a ({key_s1[9], key_s0[9]}), .c ({new_AGEMA_signal_1093, keyFF_inputPar[9]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_10_U1 ( .s (reset), .b ({new_AGEMA_signal_1094, keyFF_outputPar[13]}), .a ({key_s1[10], key_s0[10]}), .c ({new_AGEMA_signal_1096, keyFF_inputPar[10]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_11_U1 ( .s (reset), .b ({new_AGEMA_signal_1097, keyFF_outputPar[14]}), .a ({key_s1[11], key_s0[11]}), .c ({new_AGEMA_signal_1099, keyFF_inputPar[11]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_12_U1 ( .s (reset), .b ({new_AGEMA_signal_1100, keyFF_outputPar[15]}), .a ({key_s1[12], key_s0[12]}), .c ({new_AGEMA_signal_1102, keyFF_inputPar[12]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_13_U1 ( .s (reset), .b ({new_AGEMA_signal_1103, keyFF_outputPar[16]}), .a ({key_s1[13], key_s0[13]}), .c ({new_AGEMA_signal_1105, keyFF_inputPar[13]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_14_U1 ( .s (reset), .b ({new_AGEMA_signal_1106, keyFF_outputPar[17]}), .a ({key_s1[14], key_s0[14]}), .c ({new_AGEMA_signal_1108, keyFF_inputPar[14]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_15_U1 ( .s (reset), .b ({new_AGEMA_signal_1063, keyFF_counterAdd[0]}), .a ({key_s1[15], key_s0[15]}), .c ({new_AGEMA_signal_1277, keyFF_inputPar[15]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_16_U1 ( .s (reset), .b ({new_AGEMA_signal_1275, keyFF_counterAdd[1]}), .a ({key_s1[16], key_s0[16]}), .c ({new_AGEMA_signal_1285, keyFF_inputPar[16]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_17_U1 ( .s (reset), .b ({new_AGEMA_signal_1061, keyFF_counterAdd[2]}), .a ({key_s1[17], key_s0[17]}), .c ({new_AGEMA_signal_1279, keyFF_inputPar[17]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_18_U1 ( .s (reset), .b ({new_AGEMA_signal_1059, keyFF_counterAdd[3]}), .a ({key_s1[18], key_s0[18]}), .c ({new_AGEMA_signal_1281, keyFF_inputPar[18]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_19_U1 ( .s (reset), .b ({new_AGEMA_signal_1057, keyFF_counterAdd[4]}), .a ({key_s1[19], key_s0[19]}), .c ({new_AGEMA_signal_1283, keyFF_inputPar[19]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_20_U1 ( .s (reset), .b ({new_AGEMA_signal_1109, keyFF_outputPar[23]}), .a ({key_s1[20], key_s0[20]}), .c ({new_AGEMA_signal_1111, keyFF_inputPar[20]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_21_U1 ( .s (reset), .b ({new_AGEMA_signal_1112, keyFF_outputPar[24]}), .a ({key_s1[21], key_s0[21]}), .c ({new_AGEMA_signal_1114, keyFF_inputPar[21]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_22_U1 ( .s (reset), .b ({new_AGEMA_signal_1115, keyFF_outputPar[25]}), .a ({key_s1[22], key_s0[22]}), .c ({new_AGEMA_signal_1117, keyFF_inputPar[22]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_23_U1 ( .s (reset), .b ({new_AGEMA_signal_1118, keyFF_outputPar[26]}), .a ({key_s1[23], key_s0[23]}), .c ({new_AGEMA_signal_1120, keyFF_inputPar[23]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_24_U1 ( .s (reset), .b ({new_AGEMA_signal_1121, keyFF_outputPar[27]}), .a ({key_s1[24], key_s0[24]}), .c ({new_AGEMA_signal_1123, keyFF_inputPar[24]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_25_U1 ( .s (reset), .b ({new_AGEMA_signal_1124, keyFF_outputPar[28]}), .a ({key_s1[25], key_s0[25]}), .c ({new_AGEMA_signal_1126, keyFF_inputPar[25]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_26_U1 ( .s (reset), .b ({new_AGEMA_signal_1127, keyFF_outputPar[29]}), .a ({key_s1[26], key_s0[26]}), .c ({new_AGEMA_signal_1129, keyFF_inputPar[26]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_27_U1 ( .s (reset), .b ({new_AGEMA_signal_1130, keyFF_outputPar[30]}), .a ({key_s1[27], key_s0[27]}), .c ({new_AGEMA_signal_1132, keyFF_inputPar[27]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_28_U1 ( .s (reset), .b ({new_AGEMA_signal_1133, keyFF_outputPar[31]}), .a ({key_s1[28], key_s0[28]}), .c ({new_AGEMA_signal_1135, keyFF_inputPar[28]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_29_U1 ( .s (reset), .b ({new_AGEMA_signal_1136, keyFF_outputPar[32]}), .a ({key_s1[29], key_s0[29]}), .c ({new_AGEMA_signal_1138, keyFF_inputPar[29]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_30_U1 ( .s (reset), .b ({new_AGEMA_signal_1139, keyFF_outputPar[33]}), .a ({key_s1[30], key_s0[30]}), .c ({new_AGEMA_signal_1141, keyFF_inputPar[30]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_31_U1 ( .s (reset), .b ({new_AGEMA_signal_1142, keyFF_outputPar[34]}), .a ({key_s1[31], key_s0[31]}), .c ({new_AGEMA_signal_1144, keyFF_inputPar[31]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_32_U1 ( .s (reset), .b ({new_AGEMA_signal_1145, keyFF_outputPar[35]}), .a ({key_s1[32], key_s0[32]}), .c ({new_AGEMA_signal_1147, keyFF_inputPar[32]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_33_U1 ( .s (reset), .b ({new_AGEMA_signal_1148, keyFF_outputPar[36]}), .a ({key_s1[33], key_s0[33]}), .c ({new_AGEMA_signal_1150, keyFF_inputPar[33]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_34_U1 ( .s (reset), .b ({new_AGEMA_signal_1151, keyFF_outputPar[37]}), .a ({key_s1[34], key_s0[34]}), .c ({new_AGEMA_signal_1153, keyFF_inputPar[34]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_35_U1 ( .s (reset), .b ({new_AGEMA_signal_1154, keyFF_outputPar[38]}), .a ({key_s1[35], key_s0[35]}), .c ({new_AGEMA_signal_1156, keyFF_inputPar[35]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_36_U1 ( .s (reset), .b ({new_AGEMA_signal_1157, keyFF_outputPar[39]}), .a ({key_s1[36], key_s0[36]}), .c ({new_AGEMA_signal_1159, keyFF_inputPar[36]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_37_U1 ( .s (reset), .b ({new_AGEMA_signal_1160, keyFF_outputPar[40]}), .a ({key_s1[37], key_s0[37]}), .c ({new_AGEMA_signal_1162, keyFF_inputPar[37]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_38_U1 ( .s (reset), .b ({new_AGEMA_signal_1163, keyFF_outputPar[41]}), .a ({key_s1[38], key_s0[38]}), .c ({new_AGEMA_signal_1165, keyFF_inputPar[38]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_39_U1 ( .s (reset), .b ({new_AGEMA_signal_1166, keyFF_outputPar[42]}), .a ({key_s1[39], key_s0[39]}), .c ({new_AGEMA_signal_1168, keyFF_inputPar[39]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_40_U1 ( .s (reset), .b ({new_AGEMA_signal_1169, keyFF_outputPar[43]}), .a ({key_s1[40], key_s0[40]}), .c ({new_AGEMA_signal_1171, keyFF_inputPar[40]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_41_U1 ( .s (reset), .b ({new_AGEMA_signal_1172, keyFF_outputPar[44]}), .a ({key_s1[41], key_s0[41]}), .c ({new_AGEMA_signal_1174, keyFF_inputPar[41]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_42_U1 ( .s (reset), .b ({new_AGEMA_signal_1175, keyFF_outputPar[45]}), .a ({key_s1[42], key_s0[42]}), .c ({new_AGEMA_signal_1177, keyFF_inputPar[42]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_43_U1 ( .s (reset), .b ({new_AGEMA_signal_1178, keyFF_outputPar[46]}), .a ({key_s1[43], key_s0[43]}), .c ({new_AGEMA_signal_1180, keyFF_inputPar[43]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_44_U1 ( .s (reset), .b ({new_AGEMA_signal_1181, keyFF_outputPar[47]}), .a ({key_s1[44], key_s0[44]}), .c ({new_AGEMA_signal_1183, keyFF_inputPar[44]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_45_U1 ( .s (reset), .b ({new_AGEMA_signal_1184, keyFF_outputPar[48]}), .a ({key_s1[45], key_s0[45]}), .c ({new_AGEMA_signal_1186, keyFF_inputPar[45]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_46_U1 ( .s (reset), .b ({new_AGEMA_signal_1187, keyFF_outputPar[49]}), .a ({key_s1[46], key_s0[46]}), .c ({new_AGEMA_signal_1189, keyFF_inputPar[46]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_47_U1 ( .s (reset), .b ({new_AGEMA_signal_1190, keyFF_outputPar[50]}), .a ({key_s1[47], key_s0[47]}), .c ({new_AGEMA_signal_1192, keyFF_inputPar[47]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_48_U1 ( .s (reset), .b ({new_AGEMA_signal_1193, keyFF_outputPar[51]}), .a ({key_s1[48], key_s0[48]}), .c ({new_AGEMA_signal_1195, keyFF_inputPar[48]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_49_U1 ( .s (reset), .b ({new_AGEMA_signal_1196, keyFF_outputPar[52]}), .a ({key_s1[49], key_s0[49]}), .c ({new_AGEMA_signal_1198, keyFF_inputPar[49]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_50_U1 ( .s (reset), .b ({new_AGEMA_signal_1199, keyFF_outputPar[53]}), .a ({key_s1[50], key_s0[50]}), .c ({new_AGEMA_signal_1201, keyFF_inputPar[50]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_51_U1 ( .s (reset), .b ({new_AGEMA_signal_1202, keyFF_outputPar[54]}), .a ({key_s1[51], key_s0[51]}), .c ({new_AGEMA_signal_1204, keyFF_inputPar[51]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_52_U1 ( .s (reset), .b ({new_AGEMA_signal_1205, keyFF_outputPar[55]}), .a ({key_s1[52], key_s0[52]}), .c ({new_AGEMA_signal_1207, keyFF_inputPar[52]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_53_U1 ( .s (reset), .b ({new_AGEMA_signal_1208, keyFF_outputPar[56]}), .a ({key_s1[53], key_s0[53]}), .c ({new_AGEMA_signal_1210, keyFF_inputPar[53]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_54_U1 ( .s (reset), .b ({new_AGEMA_signal_1211, keyFF_outputPar[57]}), .a ({key_s1[54], key_s0[54]}), .c ({new_AGEMA_signal_1213, keyFF_inputPar[54]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_55_U1 ( .s (reset), .b ({new_AGEMA_signal_1214, keyFF_outputPar[58]}), .a ({key_s1[55], key_s0[55]}), .c ({new_AGEMA_signal_1216, keyFF_inputPar[55]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_56_U1 ( .s (reset), .b ({new_AGEMA_signal_1217, keyFF_outputPar[59]}), .a ({key_s1[56], key_s0[56]}), .c ({new_AGEMA_signal_1219, keyFF_inputPar[56]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_57_U1 ( .s (reset), .b ({new_AGEMA_signal_1220, keyFF_outputPar[60]}), .a ({key_s1[57], key_s0[57]}), .c ({new_AGEMA_signal_1222, keyFF_inputPar[57]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_58_U1 ( .s (reset), .b ({new_AGEMA_signal_1223, keyFF_outputPar[61]}), .a ({key_s1[58], key_s0[58]}), .c ({new_AGEMA_signal_1225, keyFF_inputPar[58]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_59_U1 ( .s (reset), .b ({new_AGEMA_signal_1226, keyFF_outputPar[62]}), .a ({key_s1[59], key_s0[59]}), .c ({new_AGEMA_signal_1228, keyFF_inputPar[59]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_60_U1 ( .s (reset), .b ({new_AGEMA_signal_1229, keyFF_outputPar[63]}), .a ({key_s1[60], key_s0[60]}), .c ({new_AGEMA_signal_1231, keyFF_inputPar[60]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_61_U1 ( .s (reset), .b ({new_AGEMA_signal_1232, keyFF_outputPar[64]}), .a ({key_s1[61], key_s0[61]}), .c ({new_AGEMA_signal_1234, keyFF_inputPar[61]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_62_U1 ( .s (reset), .b ({new_AGEMA_signal_1235, keyFF_outputPar[65]}), .a ({key_s1[62], key_s0[62]}), .c ({new_AGEMA_signal_1237, keyFF_inputPar[62]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_63_U1 ( .s (reset), .b ({new_AGEMA_signal_1238, keyFF_outputPar[66]}), .a ({key_s1[63], key_s0[63]}), .c ({new_AGEMA_signal_1240, keyFF_inputPar[63]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_64_U1 ( .s (reset), .b ({new_AGEMA_signal_1241, keyFF_outputPar[67]}), .a ({key_s1[64], key_s0[64]}), .c ({new_AGEMA_signal_1243, keyFF_inputPar[64]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_65_U1 ( .s (reset), .b ({new_AGEMA_signal_1244, keyFF_outputPar[68]}), .a ({key_s1[65], key_s0[65]}), .c ({new_AGEMA_signal_1246, keyFF_inputPar[65]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_66_U1 ( .s (reset), .b ({new_AGEMA_signal_1247, keyFF_outputPar[69]}), .a ({key_s1[66], key_s0[66]}), .c ({new_AGEMA_signal_1249, keyFF_inputPar[66]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_67_U1 ( .s (reset), .b ({new_AGEMA_signal_1250, keyFF_outputPar[70]}), .a ({key_s1[67], key_s0[67]}), .c ({new_AGEMA_signal_1252, keyFF_inputPar[67]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_68_U1 ( .s (reset), .b ({new_AGEMA_signal_1253, keyFF_outputPar[71]}), .a ({key_s1[68], key_s0[68]}), .c ({new_AGEMA_signal_1255, keyFF_inputPar[68]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_69_U1 ( .s (reset), .b ({new_AGEMA_signal_1256, keyFF_outputPar[72]}), .a ({key_s1[69], key_s0[69]}), .c ({new_AGEMA_signal_1258, keyFF_inputPar[69]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_70_U1 ( .s (reset), .b ({new_AGEMA_signal_1259, keyFF_outputPar[73]}), .a ({key_s1[70], key_s0[70]}), .c ({new_AGEMA_signal_1261, keyFF_inputPar[70]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_71_U1 ( .s (reset), .b ({new_AGEMA_signal_1262, keyFF_outputPar[74]}), .a ({key_s1[71], key_s0[71]}), .c ({new_AGEMA_signal_1264, keyFF_inputPar[71]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_72_U1 ( .s (reset), .b ({new_AGEMA_signal_1265, keyFF_outputPar[75]}), .a ({key_s1[72], key_s0[72]}), .c ({new_AGEMA_signal_1267, keyFF_inputPar[72]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_73_U1 ( .s (reset), .b ({new_AGEMA_signal_856, roundkey[0]}), .a ({key_s1[73], key_s0[73]}), .c ({new_AGEMA_signal_1269, keyFF_inputPar[73]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_74_U1 ( .s (reset), .b ({new_AGEMA_signal_859, roundkey[1]}), .a ({key_s1[74], key_s0[74]}), .c ({new_AGEMA_signal_1271, keyFF_inputPar[74]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_75_U1 ( .s (reset), .b ({new_AGEMA_signal_862, roundkey[2]}), .a ({key_s1[75], key_s0[75]}), .c ({new_AGEMA_signal_1273, keyFF_inputPar[75]}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) sboxInst_U3 ( .a ({new_AGEMA_signal_1295, sboxInst_L0}), .b ({new_AGEMA_signal_1311, sboxInst_n1}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) sboxInst_U2 ( .a ({new_AGEMA_signal_1292, sboxIn[3]}), .b ({new_AGEMA_signal_1293, sboxInst_n2}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) sboxInst_U1 ( .a ({new_AGEMA_signal_1288, sboxIn[1]}), .b ({new_AGEMA_signal_1294, sboxInst_n3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR1_U1 ( .a ({new_AGEMA_signal_1290, sboxIn[2]}), .b ({new_AGEMA_signal_1288, sboxIn[1]}), .c ({new_AGEMA_signal_1295, sboxInst_L0}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR2_U1 ( .a ({new_AGEMA_signal_1288, sboxIn[1]}), .b ({new_AGEMA_signal_1286, sboxIn[0]}), .c ({new_AGEMA_signal_1296, sboxInst_L1}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR3_U1 ( .a ({new_AGEMA_signal_1296, sboxInst_L1}), .b ({new_AGEMA_signal_1292, sboxIn[3]}), .c ({new_AGEMA_signal_1312, sboxInst_L2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR4_U1 ( .a ({new_AGEMA_signal_1292, sboxIn[3]}), .b ({new_AGEMA_signal_1286, sboxIn[0]}), .c ({new_AGEMA_signal_1297, sboxInst_L3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR5_U1 ( .a ({new_AGEMA_signal_1297, sboxInst_L3}), .b ({new_AGEMA_signal_1295, sboxInst_L0}), .c ({new_AGEMA_signal_1313, sboxInst_Q3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR6_U1 ( .a ({new_AGEMA_signal_1292, sboxIn[3]}), .b ({new_AGEMA_signal_1288, sboxIn[1]}), .c ({new_AGEMA_signal_1298, sboxInst_L4}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR9_U1 ( .a ({new_AGEMA_signal_1296, sboxInst_L1}), .b ({new_AGEMA_signal_1290, sboxIn[2]}), .c ({new_AGEMA_signal_1314, sboxInst_Q7}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MUX_sboxin_mux_inst_0_U1 ( .s (selSbox), .b ({new_AGEMA_signal_858, stateXORroundkey[0]}), .a ({new_AGEMA_signal_865, roundkey[3]}), .c ({new_AGEMA_signal_1286, sboxIn[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MUX_sboxin_mux_inst_1_U1 ( .s (selSbox), .b ({new_AGEMA_signal_861, stateXORroundkey[1]}), .a ({new_AGEMA_signal_1287, keyRegKS[1]}), .c ({new_AGEMA_signal_1288, sboxIn[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MUX_sboxin_mux_inst_2_U1 ( .s (selSbox), .b ({new_AGEMA_signal_864, stateXORroundkey[2]}), .a ({new_AGEMA_signal_1289, keyRegKS[2]}), .c ({new_AGEMA_signal_1290, sboxIn[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MUX_sboxin_mux_inst_3_U1 ( .s (selSbox), .b ({new_AGEMA_signal_867, stateXORroundkey[3]}), .a ({new_AGEMA_signal_1291, keyRegKS[3]}), .c ({new_AGEMA_signal_1292, sboxIn[3]}) ) ;

    /* cells in depth 1 */
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_1_MUX_inst1_mux_inst_0_U1 ( .s (new_AGEMA_signal_1480), .b ({new_AGEMA_signal_1446, serialIn[0]}), .a ({new_AGEMA_signal_1482, new_AGEMA_signal_1481}), .c ({new_AGEMA_signal_1447, stateFF_state_gff_1_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_0_U1 ( .s (new_AGEMA_signal_1483), .b ({new_AGEMA_signal_1485, new_AGEMA_signal_1484}), .a ({new_AGEMA_signal_1443, keyFF_inputPar[76]}), .c ({new_AGEMA_signal_1448, keyFF_keystate_gff_20_s_next_state[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_76_U1 ( .s (new_AGEMA_signal_1486), .b ({new_AGEMA_signal_1317, sboxOut[0]}), .a ({new_AGEMA_signal_1488, new_AGEMA_signal_1487}), .c ({new_AGEMA_signal_1443, keyFF_inputPar[76]}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR16_U1 ( .a ({new_AGEMA_signal_1316, sboxInst_T0}), .b ({new_AGEMA_signal_1490, new_AGEMA_signal_1489}), .c ({new_AGEMA_signal_1444, sboxInst_Q2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR7_U1 ( .a ({new_AGEMA_signal_1316, sboxInst_T0}), .b ({new_AGEMA_signal_1315, sboxInst_T2}), .c ({new_AGEMA_signal_1445, sboxInst_L5}) ) ;
    xnor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR8_U1 ( .a ({new_AGEMA_signal_1492, new_AGEMA_signal_1491}), .b ({new_AGEMA_signal_1445, sboxInst_L5}), .c ({new_AGEMA_signal_1449, sboxInst_Q6}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_AND1_U1 ( .a ({new_AGEMA_signal_1311, sboxInst_n1}), .b ({new_AGEMA_signal_1293, sboxInst_n2}), .clk (clk), .r ({Fresh[1], Fresh[0]}), .c ({new_AGEMA_signal_1316, sboxInst_T0}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_AND3_U1 ( .a ({new_AGEMA_signal_1294, sboxInst_n3}), .b ({new_AGEMA_signal_1290, sboxIn[2]}), .clk (clk), .r ({Fresh[3], Fresh[2]}), .c ({new_AGEMA_signal_1315, sboxInst_T2}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR15_U1 ( .a ({new_AGEMA_signal_1494, new_AGEMA_signal_1493}), .b ({new_AGEMA_signal_1315, sboxInst_T2}), .c ({new_AGEMA_signal_1317, sboxOut[0]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MUX_serialIn_mux_inst_0_U1 ( .s (new_AGEMA_signal_1495), .b ({new_AGEMA_signal_1317, sboxOut[0]}), .a ({new_AGEMA_signal_1497, new_AGEMA_signal_1496}), .c ({new_AGEMA_signal_1446, serialIn[0]}) ) ;
    buf_clk new_AGEMA_reg_buffer_704 ( .C (clk), .D (ctrlData_0_), .Q (new_AGEMA_signal_1480) ) ;
    buf_clk new_AGEMA_reg_buffer_705 ( .C (clk), .D (stateFF_inputPar[0]), .Q (new_AGEMA_signal_1481) ) ;
    buf_clk new_AGEMA_reg_buffer_706 ( .C (clk), .D (new_AGEMA_signal_870), .Q (new_AGEMA_signal_1482) ) ;
    buf_clk new_AGEMA_reg_buffer_707 ( .C (clk), .D (keyFF_keystate_n6), .Q (new_AGEMA_signal_1483) ) ;
    buf_clk new_AGEMA_reg_buffer_708 ( .C (clk), .D (keyFF_outputPar[72]), .Q (new_AGEMA_signal_1484) ) ;
    buf_clk new_AGEMA_reg_buffer_709 ( .C (clk), .D (new_AGEMA_signal_1256), .Q (new_AGEMA_signal_1485) ) ;
    buf_clk new_AGEMA_reg_buffer_710 ( .C (clk), .D (reset), .Q (new_AGEMA_signal_1486) ) ;
    buf_clk new_AGEMA_reg_buffer_711 ( .C (clk), .D (key_s0[76]), .Q (new_AGEMA_signal_1487) ) ;
    buf_clk new_AGEMA_reg_buffer_712 ( .C (clk), .D (key_s1[76]), .Q (new_AGEMA_signal_1488) ) ;
    buf_clk new_AGEMA_reg_buffer_713 ( .C (clk), .D (sboxInst_L2), .Q (new_AGEMA_signal_1489) ) ;
    buf_clk new_AGEMA_reg_buffer_714 ( .C (clk), .D (new_AGEMA_signal_1312), .Q (new_AGEMA_signal_1490) ) ;
    buf_clk new_AGEMA_reg_buffer_715 ( .C (clk), .D (sboxInst_L4), .Q (new_AGEMA_signal_1491) ) ;
    buf_clk new_AGEMA_reg_buffer_716 ( .C (clk), .D (new_AGEMA_signal_1298), .Q (new_AGEMA_signal_1492) ) ;
    buf_clk new_AGEMA_reg_buffer_717 ( .C (clk), .D (sboxInst_L3), .Q (new_AGEMA_signal_1493) ) ;
    buf_clk new_AGEMA_reg_buffer_718 ( .C (clk), .D (new_AGEMA_signal_1297), .Q (new_AGEMA_signal_1494) ) ;
    buf_clk new_AGEMA_reg_buffer_719 ( .C (clk), .D (intDone), .Q (new_AGEMA_signal_1495) ) ;
    buf_clk new_AGEMA_reg_buffer_720 ( .C (clk), .D (stateXORroundkey[0]), .Q (new_AGEMA_signal_1496) ) ;
    buf_clk new_AGEMA_reg_buffer_721 ( .C (clk), .D (new_AGEMA_signal_858), .Q (new_AGEMA_signal_1497) ) ;
    buf_clk new_AGEMA_reg_buffer_723 ( .C (clk), .D (stateFF_inputPar[1]), .Q (new_AGEMA_signal_1499) ) ;
    buf_clk new_AGEMA_reg_buffer_725 ( .C (clk), .D (new_AGEMA_signal_873), .Q (new_AGEMA_signal_1501) ) ;
    buf_clk new_AGEMA_reg_buffer_727 ( .C (clk), .D (stateFF_inputPar[2]), .Q (new_AGEMA_signal_1503) ) ;
    buf_clk new_AGEMA_reg_buffer_729 ( .C (clk), .D (new_AGEMA_signal_876), .Q (new_AGEMA_signal_1505) ) ;
    buf_clk new_AGEMA_reg_buffer_731 ( .C (clk), .D (stateFF_inputPar[3]), .Q (new_AGEMA_signal_1507) ) ;
    buf_clk new_AGEMA_reg_buffer_733 ( .C (clk), .D (new_AGEMA_signal_879), .Q (new_AGEMA_signal_1509) ) ;
    buf_clk new_AGEMA_reg_buffer_736 ( .C (clk), .D (keyFF_outputPar[73]), .Q (new_AGEMA_signal_1512) ) ;
    buf_clk new_AGEMA_reg_buffer_738 ( .C (clk), .D (new_AGEMA_signal_1259), .Q (new_AGEMA_signal_1514) ) ;
    buf_clk new_AGEMA_reg_buffer_740 ( .C (clk), .D (keyFF_outputPar[74]), .Q (new_AGEMA_signal_1516) ) ;
    buf_clk new_AGEMA_reg_buffer_742 ( .C (clk), .D (new_AGEMA_signal_1262), .Q (new_AGEMA_signal_1518) ) ;
    buf_clk new_AGEMA_reg_buffer_744 ( .C (clk), .D (keyFF_outputPar[75]), .Q (new_AGEMA_signal_1520) ) ;
    buf_clk new_AGEMA_reg_buffer_746 ( .C (clk), .D (new_AGEMA_signal_1265), .Q (new_AGEMA_signal_1522) ) ;
    buf_clk new_AGEMA_reg_buffer_749 ( .C (clk), .D (key_s0[77]), .Q (new_AGEMA_signal_1525) ) ;
    buf_clk new_AGEMA_reg_buffer_751 ( .C (clk), .D (key_s1[77]), .Q (new_AGEMA_signal_1527) ) ;
    buf_clk new_AGEMA_reg_buffer_753 ( .C (clk), .D (key_s0[78]), .Q (new_AGEMA_signal_1529) ) ;
    buf_clk new_AGEMA_reg_buffer_755 ( .C (clk), .D (key_s1[78]), .Q (new_AGEMA_signal_1531) ) ;
    buf_clk new_AGEMA_reg_buffer_757 ( .C (clk), .D (key_s0[79]), .Q (new_AGEMA_signal_1533) ) ;
    buf_clk new_AGEMA_reg_buffer_759 ( .C (clk), .D (key_s1[79]), .Q (new_AGEMA_signal_1535) ) ;
    buf_clk new_AGEMA_reg_buffer_761 ( .C (clk), .D (sboxInst_Q3), .Q (new_AGEMA_signal_1537) ) ;
    buf_clk new_AGEMA_reg_buffer_762 ( .C (clk), .D (new_AGEMA_signal_1313), .Q (new_AGEMA_signal_1538) ) ;
    buf_clk new_AGEMA_reg_buffer_763 ( .C (clk), .D (sboxInst_Q7), .Q (new_AGEMA_signal_1539) ) ;
    buf_clk new_AGEMA_reg_buffer_764 ( .C (clk), .D (new_AGEMA_signal_1314), .Q (new_AGEMA_signal_1540) ) ;
    buf_clk new_AGEMA_reg_buffer_767 ( .C (clk), .D (sboxIn[0]), .Q (new_AGEMA_signal_1543) ) ;
    buf_clk new_AGEMA_reg_buffer_769 ( .C (clk), .D (new_AGEMA_signal_1286), .Q (new_AGEMA_signal_1545) ) ;
    buf_clk new_AGEMA_reg_buffer_771 ( .C (clk), .D (sboxInst_L1), .Q (new_AGEMA_signal_1547) ) ;
    buf_clk new_AGEMA_reg_buffer_773 ( .C (clk), .D (new_AGEMA_signal_1296), .Q (new_AGEMA_signal_1549) ) ;
    buf_clk new_AGEMA_reg_buffer_778 ( .C (clk), .D (stateXORroundkey[1]), .Q (new_AGEMA_signal_1554) ) ;
    buf_clk new_AGEMA_reg_buffer_780 ( .C (clk), .D (new_AGEMA_signal_861), .Q (new_AGEMA_signal_1556) ) ;
    buf_clk new_AGEMA_reg_buffer_782 ( .C (clk), .D (stateXORroundkey[2]), .Q (new_AGEMA_signal_1558) ) ;
    buf_clk new_AGEMA_reg_buffer_784 ( .C (clk), .D (new_AGEMA_signal_864), .Q (new_AGEMA_signal_1560) ) ;
    buf_clk new_AGEMA_reg_buffer_786 ( .C (clk), .D (stateXORroundkey[3]), .Q (new_AGEMA_signal_1562) ) ;
    buf_clk new_AGEMA_reg_buffer_788 ( .C (clk), .D (new_AGEMA_signal_867), .Q (new_AGEMA_signal_1564) ) ;
    buf_clk new_AGEMA_reg_buffer_790 ( .C (clk), .D (fsm_cnt_rnd_n14), .Q (new_AGEMA_signal_1566) ) ;
    buf_clk new_AGEMA_reg_buffer_792 ( .C (clk), .D (fsm_cnt_rnd_n16), .Q (new_AGEMA_signal_1568) ) ;
    buf_clk new_AGEMA_reg_buffer_794 ( .C (clk), .D (fsm_cnt_rnd_n18), .Q (new_AGEMA_signal_1570) ) ;
    buf_clk new_AGEMA_reg_buffer_796 ( .C (clk), .D (fsm_cnt_rnd_n1), .Q (new_AGEMA_signal_1572) ) ;
    buf_clk new_AGEMA_reg_buffer_798 ( .C (clk), .D (fsm_cnt_rnd_n41), .Q (new_AGEMA_signal_1574) ) ;
    buf_clk new_AGEMA_reg_buffer_800 ( .C (clk), .D (fsm_cnt_ser_n1), .Q (new_AGEMA_signal_1576) ) ;
    buf_clk new_AGEMA_reg_buffer_802 ( .C (clk), .D (fsm_cnt_ser_n3), .Q (new_AGEMA_signal_1578) ) ;
    buf_clk new_AGEMA_reg_buffer_804 ( .C (clk), .D (fsm_cnt_ser_n26), .Q (new_AGEMA_signal_1580) ) ;
    buf_clk new_AGEMA_reg_buffer_806 ( .C (clk), .D (fsm_cnt_ser_n28), .Q (new_AGEMA_signal_1582) ) ;
    buf_clk new_AGEMA_reg_buffer_808 ( .C (clk), .D (fsm_n21), .Q (new_AGEMA_signal_1584) ) ;
    buf_clk new_AGEMA_reg_buffer_810 ( .C (clk), .D (fsm_n20), .Q (new_AGEMA_signal_1586) ) ;
    buf_clk new_AGEMA_reg_buffer_814 ( .C (clk), .D (stateFF_state_gff_2_s_next_state[3]), .Q (new_AGEMA_signal_1590) ) ;
    buf_clk new_AGEMA_reg_buffer_816 ( .C (clk), .D (new_AGEMA_signal_1302), .Q (new_AGEMA_signal_1592) ) ;
    buf_clk new_AGEMA_reg_buffer_818 ( .C (clk), .D (stateFF_state_gff_2_s_next_state[2]), .Q (new_AGEMA_signal_1594) ) ;
    buf_clk new_AGEMA_reg_buffer_820 ( .C (clk), .D (new_AGEMA_signal_1301), .Q (new_AGEMA_signal_1596) ) ;
    buf_clk new_AGEMA_reg_buffer_822 ( .C (clk), .D (stateFF_state_gff_2_s_next_state[1]), .Q (new_AGEMA_signal_1598) ) ;
    buf_clk new_AGEMA_reg_buffer_824 ( .C (clk), .D (new_AGEMA_signal_1300), .Q (new_AGEMA_signal_1600) ) ;
    buf_clk new_AGEMA_reg_buffer_826 ( .C (clk), .D (stateFF_state_gff_2_s_next_state[0]), .Q (new_AGEMA_signal_1602) ) ;
    buf_clk new_AGEMA_reg_buffer_828 ( .C (clk), .D (new_AGEMA_signal_1299), .Q (new_AGEMA_signal_1604) ) ;
    buf_clk new_AGEMA_reg_buffer_830 ( .C (clk), .D (stateFF_state_gff_3_s_next_state[3]), .Q (new_AGEMA_signal_1606) ) ;
    buf_clk new_AGEMA_reg_buffer_832 ( .C (clk), .D (new_AGEMA_signal_1321), .Q (new_AGEMA_signal_1608) ) ;
    buf_clk new_AGEMA_reg_buffer_834 ( .C (clk), .D (stateFF_state_gff_3_s_next_state[2]), .Q (new_AGEMA_signal_1610) ) ;
    buf_clk new_AGEMA_reg_buffer_836 ( .C (clk), .D (new_AGEMA_signal_1320), .Q (new_AGEMA_signal_1612) ) ;
    buf_clk new_AGEMA_reg_buffer_838 ( .C (clk), .D (stateFF_state_gff_3_s_next_state[1]), .Q (new_AGEMA_signal_1614) ) ;
    buf_clk new_AGEMA_reg_buffer_840 ( .C (clk), .D (new_AGEMA_signal_1319), .Q (new_AGEMA_signal_1616) ) ;
    buf_clk new_AGEMA_reg_buffer_842 ( .C (clk), .D (stateFF_state_gff_3_s_next_state[0]), .Q (new_AGEMA_signal_1618) ) ;
    buf_clk new_AGEMA_reg_buffer_844 ( .C (clk), .D (new_AGEMA_signal_1318), .Q (new_AGEMA_signal_1620) ) ;
    buf_clk new_AGEMA_reg_buffer_846 ( .C (clk), .D (stateFF_state_gff_4_s_next_state[3]), .Q (new_AGEMA_signal_1622) ) ;
    buf_clk new_AGEMA_reg_buffer_848 ( .C (clk), .D (new_AGEMA_signal_1325), .Q (new_AGEMA_signal_1624) ) ;
    buf_clk new_AGEMA_reg_buffer_850 ( .C (clk), .D (stateFF_state_gff_4_s_next_state[2]), .Q (new_AGEMA_signal_1626) ) ;
    buf_clk new_AGEMA_reg_buffer_852 ( .C (clk), .D (new_AGEMA_signal_1324), .Q (new_AGEMA_signal_1628) ) ;
    buf_clk new_AGEMA_reg_buffer_854 ( .C (clk), .D (stateFF_state_gff_4_s_next_state[1]), .Q (new_AGEMA_signal_1630) ) ;
    buf_clk new_AGEMA_reg_buffer_856 ( .C (clk), .D (new_AGEMA_signal_1323), .Q (new_AGEMA_signal_1632) ) ;
    buf_clk new_AGEMA_reg_buffer_858 ( .C (clk), .D (stateFF_state_gff_4_s_next_state[0]), .Q (new_AGEMA_signal_1634) ) ;
    buf_clk new_AGEMA_reg_buffer_860 ( .C (clk), .D (new_AGEMA_signal_1322), .Q (new_AGEMA_signal_1636) ) ;
    buf_clk new_AGEMA_reg_buffer_862 ( .C (clk), .D (stateFF_state_gff_5_s_next_state[3]), .Q (new_AGEMA_signal_1638) ) ;
    buf_clk new_AGEMA_reg_buffer_864 ( .C (clk), .D (new_AGEMA_signal_1329), .Q (new_AGEMA_signal_1640) ) ;
    buf_clk new_AGEMA_reg_buffer_866 ( .C (clk), .D (stateFF_state_gff_5_s_next_state[2]), .Q (new_AGEMA_signal_1642) ) ;
    buf_clk new_AGEMA_reg_buffer_868 ( .C (clk), .D (new_AGEMA_signal_1328), .Q (new_AGEMA_signal_1644) ) ;
    buf_clk new_AGEMA_reg_buffer_870 ( .C (clk), .D (stateFF_state_gff_5_s_next_state[1]), .Q (new_AGEMA_signal_1646) ) ;
    buf_clk new_AGEMA_reg_buffer_872 ( .C (clk), .D (new_AGEMA_signal_1327), .Q (new_AGEMA_signal_1648) ) ;
    buf_clk new_AGEMA_reg_buffer_874 ( .C (clk), .D (stateFF_state_gff_5_s_next_state[0]), .Q (new_AGEMA_signal_1650) ) ;
    buf_clk new_AGEMA_reg_buffer_876 ( .C (clk), .D (new_AGEMA_signal_1326), .Q (new_AGEMA_signal_1652) ) ;
    buf_clk new_AGEMA_reg_buffer_878 ( .C (clk), .D (stateFF_state_gff_6_s_next_state[3]), .Q (new_AGEMA_signal_1654) ) ;
    buf_clk new_AGEMA_reg_buffer_880 ( .C (clk), .D (new_AGEMA_signal_1333), .Q (new_AGEMA_signal_1656) ) ;
    buf_clk new_AGEMA_reg_buffer_882 ( .C (clk), .D (stateFF_state_gff_6_s_next_state[2]), .Q (new_AGEMA_signal_1658) ) ;
    buf_clk new_AGEMA_reg_buffer_884 ( .C (clk), .D (new_AGEMA_signal_1332), .Q (new_AGEMA_signal_1660) ) ;
    buf_clk new_AGEMA_reg_buffer_886 ( .C (clk), .D (stateFF_state_gff_6_s_next_state[1]), .Q (new_AGEMA_signal_1662) ) ;
    buf_clk new_AGEMA_reg_buffer_888 ( .C (clk), .D (new_AGEMA_signal_1331), .Q (new_AGEMA_signal_1664) ) ;
    buf_clk new_AGEMA_reg_buffer_890 ( .C (clk), .D (stateFF_state_gff_6_s_next_state[0]), .Q (new_AGEMA_signal_1666) ) ;
    buf_clk new_AGEMA_reg_buffer_892 ( .C (clk), .D (new_AGEMA_signal_1330), .Q (new_AGEMA_signal_1668) ) ;
    buf_clk new_AGEMA_reg_buffer_894 ( .C (clk), .D (stateFF_state_gff_7_s_next_state[3]), .Q (new_AGEMA_signal_1670) ) ;
    buf_clk new_AGEMA_reg_buffer_896 ( .C (clk), .D (new_AGEMA_signal_1337), .Q (new_AGEMA_signal_1672) ) ;
    buf_clk new_AGEMA_reg_buffer_898 ( .C (clk), .D (stateFF_state_gff_7_s_next_state[2]), .Q (new_AGEMA_signal_1674) ) ;
    buf_clk new_AGEMA_reg_buffer_900 ( .C (clk), .D (new_AGEMA_signal_1336), .Q (new_AGEMA_signal_1676) ) ;
    buf_clk new_AGEMA_reg_buffer_902 ( .C (clk), .D (stateFF_state_gff_7_s_next_state[1]), .Q (new_AGEMA_signal_1678) ) ;
    buf_clk new_AGEMA_reg_buffer_904 ( .C (clk), .D (new_AGEMA_signal_1335), .Q (new_AGEMA_signal_1680) ) ;
    buf_clk new_AGEMA_reg_buffer_906 ( .C (clk), .D (stateFF_state_gff_7_s_next_state[0]), .Q (new_AGEMA_signal_1682) ) ;
    buf_clk new_AGEMA_reg_buffer_908 ( .C (clk), .D (new_AGEMA_signal_1334), .Q (new_AGEMA_signal_1684) ) ;
    buf_clk new_AGEMA_reg_buffer_910 ( .C (clk), .D (stateFF_state_gff_8_s_next_state[3]), .Q (new_AGEMA_signal_1686) ) ;
    buf_clk new_AGEMA_reg_buffer_912 ( .C (clk), .D (new_AGEMA_signal_1341), .Q (new_AGEMA_signal_1688) ) ;
    buf_clk new_AGEMA_reg_buffer_914 ( .C (clk), .D (stateFF_state_gff_8_s_next_state[2]), .Q (new_AGEMA_signal_1690) ) ;
    buf_clk new_AGEMA_reg_buffer_916 ( .C (clk), .D (new_AGEMA_signal_1340), .Q (new_AGEMA_signal_1692) ) ;
    buf_clk new_AGEMA_reg_buffer_918 ( .C (clk), .D (stateFF_state_gff_8_s_next_state[1]), .Q (new_AGEMA_signal_1694) ) ;
    buf_clk new_AGEMA_reg_buffer_920 ( .C (clk), .D (new_AGEMA_signal_1339), .Q (new_AGEMA_signal_1696) ) ;
    buf_clk new_AGEMA_reg_buffer_922 ( .C (clk), .D (stateFF_state_gff_8_s_next_state[0]), .Q (new_AGEMA_signal_1698) ) ;
    buf_clk new_AGEMA_reg_buffer_924 ( .C (clk), .D (new_AGEMA_signal_1338), .Q (new_AGEMA_signal_1700) ) ;
    buf_clk new_AGEMA_reg_buffer_926 ( .C (clk), .D (stateFF_state_gff_9_s_next_state[3]), .Q (new_AGEMA_signal_1702) ) ;
    buf_clk new_AGEMA_reg_buffer_928 ( .C (clk), .D (new_AGEMA_signal_1345), .Q (new_AGEMA_signal_1704) ) ;
    buf_clk new_AGEMA_reg_buffer_930 ( .C (clk), .D (stateFF_state_gff_9_s_next_state[2]), .Q (new_AGEMA_signal_1706) ) ;
    buf_clk new_AGEMA_reg_buffer_932 ( .C (clk), .D (new_AGEMA_signal_1344), .Q (new_AGEMA_signal_1708) ) ;
    buf_clk new_AGEMA_reg_buffer_934 ( .C (clk), .D (stateFF_state_gff_9_s_next_state[1]), .Q (new_AGEMA_signal_1710) ) ;
    buf_clk new_AGEMA_reg_buffer_936 ( .C (clk), .D (new_AGEMA_signal_1343), .Q (new_AGEMA_signal_1712) ) ;
    buf_clk new_AGEMA_reg_buffer_938 ( .C (clk), .D (stateFF_state_gff_9_s_next_state[0]), .Q (new_AGEMA_signal_1714) ) ;
    buf_clk new_AGEMA_reg_buffer_940 ( .C (clk), .D (new_AGEMA_signal_1342), .Q (new_AGEMA_signal_1716) ) ;
    buf_clk new_AGEMA_reg_buffer_942 ( .C (clk), .D (stateFF_state_gff_10_s_next_state[3]), .Q (new_AGEMA_signal_1718) ) ;
    buf_clk new_AGEMA_reg_buffer_944 ( .C (clk), .D (new_AGEMA_signal_1349), .Q (new_AGEMA_signal_1720) ) ;
    buf_clk new_AGEMA_reg_buffer_946 ( .C (clk), .D (stateFF_state_gff_10_s_next_state[2]), .Q (new_AGEMA_signal_1722) ) ;
    buf_clk new_AGEMA_reg_buffer_948 ( .C (clk), .D (new_AGEMA_signal_1348), .Q (new_AGEMA_signal_1724) ) ;
    buf_clk new_AGEMA_reg_buffer_950 ( .C (clk), .D (stateFF_state_gff_10_s_next_state[1]), .Q (new_AGEMA_signal_1726) ) ;
    buf_clk new_AGEMA_reg_buffer_952 ( .C (clk), .D (new_AGEMA_signal_1347), .Q (new_AGEMA_signal_1728) ) ;
    buf_clk new_AGEMA_reg_buffer_954 ( .C (clk), .D (stateFF_state_gff_10_s_next_state[0]), .Q (new_AGEMA_signal_1730) ) ;
    buf_clk new_AGEMA_reg_buffer_956 ( .C (clk), .D (new_AGEMA_signal_1346), .Q (new_AGEMA_signal_1732) ) ;
    buf_clk new_AGEMA_reg_buffer_958 ( .C (clk), .D (stateFF_state_gff_11_s_next_state[3]), .Q (new_AGEMA_signal_1734) ) ;
    buf_clk new_AGEMA_reg_buffer_960 ( .C (clk), .D (new_AGEMA_signal_1353), .Q (new_AGEMA_signal_1736) ) ;
    buf_clk new_AGEMA_reg_buffer_962 ( .C (clk), .D (stateFF_state_gff_11_s_next_state[2]), .Q (new_AGEMA_signal_1738) ) ;
    buf_clk new_AGEMA_reg_buffer_964 ( .C (clk), .D (new_AGEMA_signal_1352), .Q (new_AGEMA_signal_1740) ) ;
    buf_clk new_AGEMA_reg_buffer_966 ( .C (clk), .D (stateFF_state_gff_11_s_next_state[1]), .Q (new_AGEMA_signal_1742) ) ;
    buf_clk new_AGEMA_reg_buffer_968 ( .C (clk), .D (new_AGEMA_signal_1351), .Q (new_AGEMA_signal_1744) ) ;
    buf_clk new_AGEMA_reg_buffer_970 ( .C (clk), .D (stateFF_state_gff_11_s_next_state[0]), .Q (new_AGEMA_signal_1746) ) ;
    buf_clk new_AGEMA_reg_buffer_972 ( .C (clk), .D (new_AGEMA_signal_1350), .Q (new_AGEMA_signal_1748) ) ;
    buf_clk new_AGEMA_reg_buffer_974 ( .C (clk), .D (stateFF_state_gff_12_s_next_state[3]), .Q (new_AGEMA_signal_1750) ) ;
    buf_clk new_AGEMA_reg_buffer_976 ( .C (clk), .D (new_AGEMA_signal_1357), .Q (new_AGEMA_signal_1752) ) ;
    buf_clk new_AGEMA_reg_buffer_978 ( .C (clk), .D (stateFF_state_gff_12_s_next_state[2]), .Q (new_AGEMA_signal_1754) ) ;
    buf_clk new_AGEMA_reg_buffer_980 ( .C (clk), .D (new_AGEMA_signal_1356), .Q (new_AGEMA_signal_1756) ) ;
    buf_clk new_AGEMA_reg_buffer_982 ( .C (clk), .D (stateFF_state_gff_12_s_next_state[1]), .Q (new_AGEMA_signal_1758) ) ;
    buf_clk new_AGEMA_reg_buffer_984 ( .C (clk), .D (new_AGEMA_signal_1355), .Q (new_AGEMA_signal_1760) ) ;
    buf_clk new_AGEMA_reg_buffer_986 ( .C (clk), .D (stateFF_state_gff_12_s_next_state[0]), .Q (new_AGEMA_signal_1762) ) ;
    buf_clk new_AGEMA_reg_buffer_988 ( .C (clk), .D (new_AGEMA_signal_1354), .Q (new_AGEMA_signal_1764) ) ;
    buf_clk new_AGEMA_reg_buffer_990 ( .C (clk), .D (stateFF_state_gff_13_s_next_state[3]), .Q (new_AGEMA_signal_1766) ) ;
    buf_clk new_AGEMA_reg_buffer_992 ( .C (clk), .D (new_AGEMA_signal_1361), .Q (new_AGEMA_signal_1768) ) ;
    buf_clk new_AGEMA_reg_buffer_994 ( .C (clk), .D (stateFF_state_gff_13_s_next_state[2]), .Q (new_AGEMA_signal_1770) ) ;
    buf_clk new_AGEMA_reg_buffer_996 ( .C (clk), .D (new_AGEMA_signal_1360), .Q (new_AGEMA_signal_1772) ) ;
    buf_clk new_AGEMA_reg_buffer_998 ( .C (clk), .D (stateFF_state_gff_13_s_next_state[1]), .Q (new_AGEMA_signal_1774) ) ;
    buf_clk new_AGEMA_reg_buffer_1000 ( .C (clk), .D (new_AGEMA_signal_1359), .Q (new_AGEMA_signal_1776) ) ;
    buf_clk new_AGEMA_reg_buffer_1002 ( .C (clk), .D (stateFF_state_gff_13_s_next_state[0]), .Q (new_AGEMA_signal_1778) ) ;
    buf_clk new_AGEMA_reg_buffer_1004 ( .C (clk), .D (new_AGEMA_signal_1358), .Q (new_AGEMA_signal_1780) ) ;
    buf_clk new_AGEMA_reg_buffer_1006 ( .C (clk), .D (stateFF_state_gff_14_s_next_state[3]), .Q (new_AGEMA_signal_1782) ) ;
    buf_clk new_AGEMA_reg_buffer_1008 ( .C (clk), .D (new_AGEMA_signal_1365), .Q (new_AGEMA_signal_1784) ) ;
    buf_clk new_AGEMA_reg_buffer_1010 ( .C (clk), .D (stateFF_state_gff_14_s_next_state[2]), .Q (new_AGEMA_signal_1786) ) ;
    buf_clk new_AGEMA_reg_buffer_1012 ( .C (clk), .D (new_AGEMA_signal_1364), .Q (new_AGEMA_signal_1788) ) ;
    buf_clk new_AGEMA_reg_buffer_1014 ( .C (clk), .D (stateFF_state_gff_14_s_next_state[1]), .Q (new_AGEMA_signal_1790) ) ;
    buf_clk new_AGEMA_reg_buffer_1016 ( .C (clk), .D (new_AGEMA_signal_1363), .Q (new_AGEMA_signal_1792) ) ;
    buf_clk new_AGEMA_reg_buffer_1018 ( .C (clk), .D (stateFF_state_gff_14_s_next_state[0]), .Q (new_AGEMA_signal_1794) ) ;
    buf_clk new_AGEMA_reg_buffer_1020 ( .C (clk), .D (new_AGEMA_signal_1362), .Q (new_AGEMA_signal_1796) ) ;
    buf_clk new_AGEMA_reg_buffer_1022 ( .C (clk), .D (stateFF_state_gff_15_s_next_state[3]), .Q (new_AGEMA_signal_1798) ) ;
    buf_clk new_AGEMA_reg_buffer_1024 ( .C (clk), .D (new_AGEMA_signal_1369), .Q (new_AGEMA_signal_1800) ) ;
    buf_clk new_AGEMA_reg_buffer_1026 ( .C (clk), .D (stateFF_state_gff_15_s_next_state[2]), .Q (new_AGEMA_signal_1802) ) ;
    buf_clk new_AGEMA_reg_buffer_1028 ( .C (clk), .D (new_AGEMA_signal_1368), .Q (new_AGEMA_signal_1804) ) ;
    buf_clk new_AGEMA_reg_buffer_1030 ( .C (clk), .D (stateFF_state_gff_15_s_next_state[1]), .Q (new_AGEMA_signal_1806) ) ;
    buf_clk new_AGEMA_reg_buffer_1032 ( .C (clk), .D (new_AGEMA_signal_1367), .Q (new_AGEMA_signal_1808) ) ;
    buf_clk new_AGEMA_reg_buffer_1034 ( .C (clk), .D (stateFF_state_gff_15_s_next_state[0]), .Q (new_AGEMA_signal_1810) ) ;
    buf_clk new_AGEMA_reg_buffer_1036 ( .C (clk), .D (new_AGEMA_signal_1366), .Q (new_AGEMA_signal_1812) ) ;
    buf_clk new_AGEMA_reg_buffer_1038 ( .C (clk), .D (stateFF_state_gff_16_s_next_state[3]), .Q (new_AGEMA_signal_1814) ) ;
    buf_clk new_AGEMA_reg_buffer_1040 ( .C (clk), .D (new_AGEMA_signal_1373), .Q (new_AGEMA_signal_1816) ) ;
    buf_clk new_AGEMA_reg_buffer_1042 ( .C (clk), .D (stateFF_state_gff_16_s_next_state[2]), .Q (new_AGEMA_signal_1818) ) ;
    buf_clk new_AGEMA_reg_buffer_1044 ( .C (clk), .D (new_AGEMA_signal_1372), .Q (new_AGEMA_signal_1820) ) ;
    buf_clk new_AGEMA_reg_buffer_1046 ( .C (clk), .D (stateFF_state_gff_16_s_next_state[1]), .Q (new_AGEMA_signal_1822) ) ;
    buf_clk new_AGEMA_reg_buffer_1048 ( .C (clk), .D (new_AGEMA_signal_1371), .Q (new_AGEMA_signal_1824) ) ;
    buf_clk new_AGEMA_reg_buffer_1050 ( .C (clk), .D (stateFF_state_gff_16_s_next_state[0]), .Q (new_AGEMA_signal_1826) ) ;
    buf_clk new_AGEMA_reg_buffer_1052 ( .C (clk), .D (new_AGEMA_signal_1370), .Q (new_AGEMA_signal_1828) ) ;
    buf_clk new_AGEMA_reg_buffer_1054 ( .C (clk), .D (keyFF_keystate_gff_1_s_next_state[3]), .Q (new_AGEMA_signal_1830) ) ;
    buf_clk new_AGEMA_reg_buffer_1056 ( .C (clk), .D (new_AGEMA_signal_1377), .Q (new_AGEMA_signal_1832) ) ;
    buf_clk new_AGEMA_reg_buffer_1058 ( .C (clk), .D (keyFF_keystate_gff_1_s_next_state[2]), .Q (new_AGEMA_signal_1834) ) ;
    buf_clk new_AGEMA_reg_buffer_1060 ( .C (clk), .D (new_AGEMA_signal_1376), .Q (new_AGEMA_signal_1836) ) ;
    buf_clk new_AGEMA_reg_buffer_1062 ( .C (clk), .D (keyFF_keystate_gff_1_s_next_state[1]), .Q (new_AGEMA_signal_1838) ) ;
    buf_clk new_AGEMA_reg_buffer_1064 ( .C (clk), .D (new_AGEMA_signal_1375), .Q (new_AGEMA_signal_1840) ) ;
    buf_clk new_AGEMA_reg_buffer_1066 ( .C (clk), .D (keyFF_keystate_gff_1_s_next_state[0]), .Q (new_AGEMA_signal_1842) ) ;
    buf_clk new_AGEMA_reg_buffer_1068 ( .C (clk), .D (new_AGEMA_signal_1374), .Q (new_AGEMA_signal_1844) ) ;
    buf_clk new_AGEMA_reg_buffer_1070 ( .C (clk), .D (keyFF_keystate_gff_2_s_next_state[3]), .Q (new_AGEMA_signal_1846) ) ;
    buf_clk new_AGEMA_reg_buffer_1072 ( .C (clk), .D (new_AGEMA_signal_1381), .Q (new_AGEMA_signal_1848) ) ;
    buf_clk new_AGEMA_reg_buffer_1074 ( .C (clk), .D (keyFF_keystate_gff_2_s_next_state[2]), .Q (new_AGEMA_signal_1850) ) ;
    buf_clk new_AGEMA_reg_buffer_1076 ( .C (clk), .D (new_AGEMA_signal_1380), .Q (new_AGEMA_signal_1852) ) ;
    buf_clk new_AGEMA_reg_buffer_1078 ( .C (clk), .D (keyFF_keystate_gff_2_s_next_state[1]), .Q (new_AGEMA_signal_1854) ) ;
    buf_clk new_AGEMA_reg_buffer_1080 ( .C (clk), .D (new_AGEMA_signal_1379), .Q (new_AGEMA_signal_1856) ) ;
    buf_clk new_AGEMA_reg_buffer_1082 ( .C (clk), .D (keyFF_keystate_gff_2_s_next_state[0]), .Q (new_AGEMA_signal_1858) ) ;
    buf_clk new_AGEMA_reg_buffer_1084 ( .C (clk), .D (new_AGEMA_signal_1378), .Q (new_AGEMA_signal_1860) ) ;
    buf_clk new_AGEMA_reg_buffer_1086 ( .C (clk), .D (keyFF_keystate_gff_3_s_next_state[3]), .Q (new_AGEMA_signal_1862) ) ;
    buf_clk new_AGEMA_reg_buffer_1088 ( .C (clk), .D (new_AGEMA_signal_1385), .Q (new_AGEMA_signal_1864) ) ;
    buf_clk new_AGEMA_reg_buffer_1090 ( .C (clk), .D (keyFF_keystate_gff_3_s_next_state[2]), .Q (new_AGEMA_signal_1866) ) ;
    buf_clk new_AGEMA_reg_buffer_1092 ( .C (clk), .D (new_AGEMA_signal_1384), .Q (new_AGEMA_signal_1868) ) ;
    buf_clk new_AGEMA_reg_buffer_1094 ( .C (clk), .D (keyFF_keystate_gff_3_s_next_state[1]), .Q (new_AGEMA_signal_1870) ) ;
    buf_clk new_AGEMA_reg_buffer_1096 ( .C (clk), .D (new_AGEMA_signal_1383), .Q (new_AGEMA_signal_1872) ) ;
    buf_clk new_AGEMA_reg_buffer_1098 ( .C (clk), .D (keyFF_keystate_gff_3_s_next_state[0]), .Q (new_AGEMA_signal_1874) ) ;
    buf_clk new_AGEMA_reg_buffer_1100 ( .C (clk), .D (new_AGEMA_signal_1382), .Q (new_AGEMA_signal_1876) ) ;
    buf_clk new_AGEMA_reg_buffer_1102 ( .C (clk), .D (keyFF_keystate_gff_4_s_next_state[3]), .Q (new_AGEMA_signal_1878) ) ;
    buf_clk new_AGEMA_reg_buffer_1104 ( .C (clk), .D (new_AGEMA_signal_1389), .Q (new_AGEMA_signal_1880) ) ;
    buf_clk new_AGEMA_reg_buffer_1106 ( .C (clk), .D (keyFF_keystate_gff_4_s_next_state[2]), .Q (new_AGEMA_signal_1882) ) ;
    buf_clk new_AGEMA_reg_buffer_1108 ( .C (clk), .D (new_AGEMA_signal_1388), .Q (new_AGEMA_signal_1884) ) ;
    buf_clk new_AGEMA_reg_buffer_1110 ( .C (clk), .D (keyFF_keystate_gff_4_s_next_state[1]), .Q (new_AGEMA_signal_1886) ) ;
    buf_clk new_AGEMA_reg_buffer_1112 ( .C (clk), .D (new_AGEMA_signal_1387), .Q (new_AGEMA_signal_1888) ) ;
    buf_clk new_AGEMA_reg_buffer_1114 ( .C (clk), .D (keyFF_keystate_gff_4_s_next_state[0]), .Q (new_AGEMA_signal_1890) ) ;
    buf_clk new_AGEMA_reg_buffer_1116 ( .C (clk), .D (new_AGEMA_signal_1386), .Q (new_AGEMA_signal_1892) ) ;
    buf_clk new_AGEMA_reg_buffer_1118 ( .C (clk), .D (keyFF_keystate_gff_5_s_next_state[3]), .Q (new_AGEMA_signal_1894) ) ;
    buf_clk new_AGEMA_reg_buffer_1120 ( .C (clk), .D (new_AGEMA_signal_1306), .Q (new_AGEMA_signal_1896) ) ;
    buf_clk new_AGEMA_reg_buffer_1122 ( .C (clk), .D (keyFF_keystate_gff_5_s_next_state[2]), .Q (new_AGEMA_signal_1898) ) ;
    buf_clk new_AGEMA_reg_buffer_1124 ( .C (clk), .D (new_AGEMA_signal_1305), .Q (new_AGEMA_signal_1900) ) ;
    buf_clk new_AGEMA_reg_buffer_1126 ( .C (clk), .D (keyFF_keystate_gff_5_s_next_state[1]), .Q (new_AGEMA_signal_1902) ) ;
    buf_clk new_AGEMA_reg_buffer_1128 ( .C (clk), .D (new_AGEMA_signal_1304), .Q (new_AGEMA_signal_1904) ) ;
    buf_clk new_AGEMA_reg_buffer_1130 ( .C (clk), .D (keyFF_keystate_gff_5_s_next_state[0]), .Q (new_AGEMA_signal_1906) ) ;
    buf_clk new_AGEMA_reg_buffer_1132 ( .C (clk), .D (new_AGEMA_signal_1303), .Q (new_AGEMA_signal_1908) ) ;
    buf_clk new_AGEMA_reg_buffer_1134 ( .C (clk), .D (keyFF_keystate_gff_6_s_next_state[3]), .Q (new_AGEMA_signal_1910) ) ;
    buf_clk new_AGEMA_reg_buffer_1136 ( .C (clk), .D (new_AGEMA_signal_1310), .Q (new_AGEMA_signal_1912) ) ;
    buf_clk new_AGEMA_reg_buffer_1138 ( .C (clk), .D (keyFF_keystate_gff_6_s_next_state[2]), .Q (new_AGEMA_signal_1914) ) ;
    buf_clk new_AGEMA_reg_buffer_1140 ( .C (clk), .D (new_AGEMA_signal_1309), .Q (new_AGEMA_signal_1916) ) ;
    buf_clk new_AGEMA_reg_buffer_1142 ( .C (clk), .D (keyFF_keystate_gff_6_s_next_state[1]), .Q (new_AGEMA_signal_1918) ) ;
    buf_clk new_AGEMA_reg_buffer_1144 ( .C (clk), .D (new_AGEMA_signal_1308), .Q (new_AGEMA_signal_1920) ) ;
    buf_clk new_AGEMA_reg_buffer_1146 ( .C (clk), .D (keyFF_keystate_gff_6_s_next_state[0]), .Q (new_AGEMA_signal_1922) ) ;
    buf_clk new_AGEMA_reg_buffer_1148 ( .C (clk), .D (new_AGEMA_signal_1307), .Q (new_AGEMA_signal_1924) ) ;
    buf_clk new_AGEMA_reg_buffer_1150 ( .C (clk), .D (keyFF_keystate_gff_7_s_next_state[3]), .Q (new_AGEMA_signal_1926) ) ;
    buf_clk new_AGEMA_reg_buffer_1152 ( .C (clk), .D (new_AGEMA_signal_1393), .Q (new_AGEMA_signal_1928) ) ;
    buf_clk new_AGEMA_reg_buffer_1154 ( .C (clk), .D (keyFF_keystate_gff_7_s_next_state[2]), .Q (new_AGEMA_signal_1930) ) ;
    buf_clk new_AGEMA_reg_buffer_1156 ( .C (clk), .D (new_AGEMA_signal_1392), .Q (new_AGEMA_signal_1932) ) ;
    buf_clk new_AGEMA_reg_buffer_1158 ( .C (clk), .D (keyFF_keystate_gff_7_s_next_state[1]), .Q (new_AGEMA_signal_1934) ) ;
    buf_clk new_AGEMA_reg_buffer_1160 ( .C (clk), .D (new_AGEMA_signal_1391), .Q (new_AGEMA_signal_1936) ) ;
    buf_clk new_AGEMA_reg_buffer_1162 ( .C (clk), .D (keyFF_keystate_gff_7_s_next_state[0]), .Q (new_AGEMA_signal_1938) ) ;
    buf_clk new_AGEMA_reg_buffer_1164 ( .C (clk), .D (new_AGEMA_signal_1390), .Q (new_AGEMA_signal_1940) ) ;
    buf_clk new_AGEMA_reg_buffer_1166 ( .C (clk), .D (keyFF_keystate_gff_8_s_next_state[3]), .Q (new_AGEMA_signal_1942) ) ;
    buf_clk new_AGEMA_reg_buffer_1168 ( .C (clk), .D (new_AGEMA_signal_1397), .Q (new_AGEMA_signal_1944) ) ;
    buf_clk new_AGEMA_reg_buffer_1170 ( .C (clk), .D (keyFF_keystate_gff_8_s_next_state[2]), .Q (new_AGEMA_signal_1946) ) ;
    buf_clk new_AGEMA_reg_buffer_1172 ( .C (clk), .D (new_AGEMA_signal_1396), .Q (new_AGEMA_signal_1948) ) ;
    buf_clk new_AGEMA_reg_buffer_1174 ( .C (clk), .D (keyFF_keystate_gff_8_s_next_state[1]), .Q (new_AGEMA_signal_1950) ) ;
    buf_clk new_AGEMA_reg_buffer_1176 ( .C (clk), .D (new_AGEMA_signal_1395), .Q (new_AGEMA_signal_1952) ) ;
    buf_clk new_AGEMA_reg_buffer_1178 ( .C (clk), .D (keyFF_keystate_gff_8_s_next_state[0]), .Q (new_AGEMA_signal_1954) ) ;
    buf_clk new_AGEMA_reg_buffer_1180 ( .C (clk), .D (new_AGEMA_signal_1394), .Q (new_AGEMA_signal_1956) ) ;
    buf_clk new_AGEMA_reg_buffer_1182 ( .C (clk), .D (keyFF_keystate_gff_9_s_next_state[3]), .Q (new_AGEMA_signal_1958) ) ;
    buf_clk new_AGEMA_reg_buffer_1184 ( .C (clk), .D (new_AGEMA_signal_1401), .Q (new_AGEMA_signal_1960) ) ;
    buf_clk new_AGEMA_reg_buffer_1186 ( .C (clk), .D (keyFF_keystate_gff_9_s_next_state[2]), .Q (new_AGEMA_signal_1962) ) ;
    buf_clk new_AGEMA_reg_buffer_1188 ( .C (clk), .D (new_AGEMA_signal_1400), .Q (new_AGEMA_signal_1964) ) ;
    buf_clk new_AGEMA_reg_buffer_1190 ( .C (clk), .D (keyFF_keystate_gff_9_s_next_state[1]), .Q (new_AGEMA_signal_1966) ) ;
    buf_clk new_AGEMA_reg_buffer_1192 ( .C (clk), .D (new_AGEMA_signal_1399), .Q (new_AGEMA_signal_1968) ) ;
    buf_clk new_AGEMA_reg_buffer_1194 ( .C (clk), .D (keyFF_keystate_gff_9_s_next_state[0]), .Q (new_AGEMA_signal_1970) ) ;
    buf_clk new_AGEMA_reg_buffer_1196 ( .C (clk), .D (new_AGEMA_signal_1398), .Q (new_AGEMA_signal_1972) ) ;
    buf_clk new_AGEMA_reg_buffer_1198 ( .C (clk), .D (keyFF_keystate_gff_10_s_next_state[3]), .Q (new_AGEMA_signal_1974) ) ;
    buf_clk new_AGEMA_reg_buffer_1200 ( .C (clk), .D (new_AGEMA_signal_1405), .Q (new_AGEMA_signal_1976) ) ;
    buf_clk new_AGEMA_reg_buffer_1202 ( .C (clk), .D (keyFF_keystate_gff_10_s_next_state[2]), .Q (new_AGEMA_signal_1978) ) ;
    buf_clk new_AGEMA_reg_buffer_1204 ( .C (clk), .D (new_AGEMA_signal_1404), .Q (new_AGEMA_signal_1980) ) ;
    buf_clk new_AGEMA_reg_buffer_1206 ( .C (clk), .D (keyFF_keystate_gff_10_s_next_state[1]), .Q (new_AGEMA_signal_1982) ) ;
    buf_clk new_AGEMA_reg_buffer_1208 ( .C (clk), .D (new_AGEMA_signal_1403), .Q (new_AGEMA_signal_1984) ) ;
    buf_clk new_AGEMA_reg_buffer_1210 ( .C (clk), .D (keyFF_keystate_gff_10_s_next_state[0]), .Q (new_AGEMA_signal_1986) ) ;
    buf_clk new_AGEMA_reg_buffer_1212 ( .C (clk), .D (new_AGEMA_signal_1402), .Q (new_AGEMA_signal_1988) ) ;
    buf_clk new_AGEMA_reg_buffer_1214 ( .C (clk), .D (keyFF_keystate_gff_11_s_next_state[3]), .Q (new_AGEMA_signal_1990) ) ;
    buf_clk new_AGEMA_reg_buffer_1216 ( .C (clk), .D (new_AGEMA_signal_1409), .Q (new_AGEMA_signal_1992) ) ;
    buf_clk new_AGEMA_reg_buffer_1218 ( .C (clk), .D (keyFF_keystate_gff_11_s_next_state[2]), .Q (new_AGEMA_signal_1994) ) ;
    buf_clk new_AGEMA_reg_buffer_1220 ( .C (clk), .D (new_AGEMA_signal_1408), .Q (new_AGEMA_signal_1996) ) ;
    buf_clk new_AGEMA_reg_buffer_1222 ( .C (clk), .D (keyFF_keystate_gff_11_s_next_state[1]), .Q (new_AGEMA_signal_1998) ) ;
    buf_clk new_AGEMA_reg_buffer_1224 ( .C (clk), .D (new_AGEMA_signal_1407), .Q (new_AGEMA_signal_2000) ) ;
    buf_clk new_AGEMA_reg_buffer_1226 ( .C (clk), .D (keyFF_keystate_gff_11_s_next_state[0]), .Q (new_AGEMA_signal_2002) ) ;
    buf_clk new_AGEMA_reg_buffer_1228 ( .C (clk), .D (new_AGEMA_signal_1406), .Q (new_AGEMA_signal_2004) ) ;
    buf_clk new_AGEMA_reg_buffer_1230 ( .C (clk), .D (keyFF_keystate_gff_12_s_next_state[3]), .Q (new_AGEMA_signal_2006) ) ;
    buf_clk new_AGEMA_reg_buffer_1232 ( .C (clk), .D (new_AGEMA_signal_1413), .Q (new_AGEMA_signal_2008) ) ;
    buf_clk new_AGEMA_reg_buffer_1234 ( .C (clk), .D (keyFF_keystate_gff_12_s_next_state[2]), .Q (new_AGEMA_signal_2010) ) ;
    buf_clk new_AGEMA_reg_buffer_1236 ( .C (clk), .D (new_AGEMA_signal_1412), .Q (new_AGEMA_signal_2012) ) ;
    buf_clk new_AGEMA_reg_buffer_1238 ( .C (clk), .D (keyFF_keystate_gff_12_s_next_state[1]), .Q (new_AGEMA_signal_2014) ) ;
    buf_clk new_AGEMA_reg_buffer_1240 ( .C (clk), .D (new_AGEMA_signal_1411), .Q (new_AGEMA_signal_2016) ) ;
    buf_clk new_AGEMA_reg_buffer_1242 ( .C (clk), .D (keyFF_keystate_gff_12_s_next_state[0]), .Q (new_AGEMA_signal_2018) ) ;
    buf_clk new_AGEMA_reg_buffer_1244 ( .C (clk), .D (new_AGEMA_signal_1410), .Q (new_AGEMA_signal_2020) ) ;
    buf_clk new_AGEMA_reg_buffer_1246 ( .C (clk), .D (keyFF_keystate_gff_13_s_next_state[3]), .Q (new_AGEMA_signal_2022) ) ;
    buf_clk new_AGEMA_reg_buffer_1248 ( .C (clk), .D (new_AGEMA_signal_1417), .Q (new_AGEMA_signal_2024) ) ;
    buf_clk new_AGEMA_reg_buffer_1250 ( .C (clk), .D (keyFF_keystate_gff_13_s_next_state[2]), .Q (new_AGEMA_signal_2026) ) ;
    buf_clk new_AGEMA_reg_buffer_1252 ( .C (clk), .D (new_AGEMA_signal_1416), .Q (new_AGEMA_signal_2028) ) ;
    buf_clk new_AGEMA_reg_buffer_1254 ( .C (clk), .D (keyFF_keystate_gff_13_s_next_state[1]), .Q (new_AGEMA_signal_2030) ) ;
    buf_clk new_AGEMA_reg_buffer_1256 ( .C (clk), .D (new_AGEMA_signal_1415), .Q (new_AGEMA_signal_2032) ) ;
    buf_clk new_AGEMA_reg_buffer_1258 ( .C (clk), .D (keyFF_keystate_gff_13_s_next_state[0]), .Q (new_AGEMA_signal_2034) ) ;
    buf_clk new_AGEMA_reg_buffer_1260 ( .C (clk), .D (new_AGEMA_signal_1414), .Q (new_AGEMA_signal_2036) ) ;
    buf_clk new_AGEMA_reg_buffer_1262 ( .C (clk), .D (keyFF_keystate_gff_14_s_next_state[3]), .Q (new_AGEMA_signal_2038) ) ;
    buf_clk new_AGEMA_reg_buffer_1264 ( .C (clk), .D (new_AGEMA_signal_1421), .Q (new_AGEMA_signal_2040) ) ;
    buf_clk new_AGEMA_reg_buffer_1266 ( .C (clk), .D (keyFF_keystate_gff_14_s_next_state[2]), .Q (new_AGEMA_signal_2042) ) ;
    buf_clk new_AGEMA_reg_buffer_1268 ( .C (clk), .D (new_AGEMA_signal_1420), .Q (new_AGEMA_signal_2044) ) ;
    buf_clk new_AGEMA_reg_buffer_1270 ( .C (clk), .D (keyFF_keystate_gff_14_s_next_state[1]), .Q (new_AGEMA_signal_2046) ) ;
    buf_clk new_AGEMA_reg_buffer_1272 ( .C (clk), .D (new_AGEMA_signal_1419), .Q (new_AGEMA_signal_2048) ) ;
    buf_clk new_AGEMA_reg_buffer_1274 ( .C (clk), .D (keyFF_keystate_gff_14_s_next_state[0]), .Q (new_AGEMA_signal_2050) ) ;
    buf_clk new_AGEMA_reg_buffer_1276 ( .C (clk), .D (new_AGEMA_signal_1418), .Q (new_AGEMA_signal_2052) ) ;
    buf_clk new_AGEMA_reg_buffer_1278 ( .C (clk), .D (keyFF_keystate_gff_15_s_next_state[3]), .Q (new_AGEMA_signal_2054) ) ;
    buf_clk new_AGEMA_reg_buffer_1280 ( .C (clk), .D (new_AGEMA_signal_1425), .Q (new_AGEMA_signal_2056) ) ;
    buf_clk new_AGEMA_reg_buffer_1282 ( .C (clk), .D (keyFF_keystate_gff_15_s_next_state[2]), .Q (new_AGEMA_signal_2058) ) ;
    buf_clk new_AGEMA_reg_buffer_1284 ( .C (clk), .D (new_AGEMA_signal_1424), .Q (new_AGEMA_signal_2060) ) ;
    buf_clk new_AGEMA_reg_buffer_1286 ( .C (clk), .D (keyFF_keystate_gff_15_s_next_state[1]), .Q (new_AGEMA_signal_2062) ) ;
    buf_clk new_AGEMA_reg_buffer_1288 ( .C (clk), .D (new_AGEMA_signal_1423), .Q (new_AGEMA_signal_2064) ) ;
    buf_clk new_AGEMA_reg_buffer_1290 ( .C (clk), .D (keyFF_keystate_gff_15_s_next_state[0]), .Q (new_AGEMA_signal_2066) ) ;
    buf_clk new_AGEMA_reg_buffer_1292 ( .C (clk), .D (new_AGEMA_signal_1422), .Q (new_AGEMA_signal_2068) ) ;
    buf_clk new_AGEMA_reg_buffer_1294 ( .C (clk), .D (keyFF_keystate_gff_16_s_next_state[3]), .Q (new_AGEMA_signal_2070) ) ;
    buf_clk new_AGEMA_reg_buffer_1296 ( .C (clk), .D (new_AGEMA_signal_1429), .Q (new_AGEMA_signal_2072) ) ;
    buf_clk new_AGEMA_reg_buffer_1298 ( .C (clk), .D (keyFF_keystate_gff_16_s_next_state[2]), .Q (new_AGEMA_signal_2074) ) ;
    buf_clk new_AGEMA_reg_buffer_1300 ( .C (clk), .D (new_AGEMA_signal_1428), .Q (new_AGEMA_signal_2076) ) ;
    buf_clk new_AGEMA_reg_buffer_1302 ( .C (clk), .D (keyFF_keystate_gff_16_s_next_state[1]), .Q (new_AGEMA_signal_2078) ) ;
    buf_clk new_AGEMA_reg_buffer_1304 ( .C (clk), .D (new_AGEMA_signal_1427), .Q (new_AGEMA_signal_2080) ) ;
    buf_clk new_AGEMA_reg_buffer_1306 ( .C (clk), .D (keyFF_keystate_gff_16_s_next_state[0]), .Q (new_AGEMA_signal_2082) ) ;
    buf_clk new_AGEMA_reg_buffer_1308 ( .C (clk), .D (new_AGEMA_signal_1426), .Q (new_AGEMA_signal_2084) ) ;
    buf_clk new_AGEMA_reg_buffer_1310 ( .C (clk), .D (keyFF_keystate_gff_17_s_next_state[3]), .Q (new_AGEMA_signal_2086) ) ;
    buf_clk new_AGEMA_reg_buffer_1312 ( .C (clk), .D (new_AGEMA_signal_1433), .Q (new_AGEMA_signal_2088) ) ;
    buf_clk new_AGEMA_reg_buffer_1314 ( .C (clk), .D (keyFF_keystate_gff_17_s_next_state[2]), .Q (new_AGEMA_signal_2090) ) ;
    buf_clk new_AGEMA_reg_buffer_1316 ( .C (clk), .D (new_AGEMA_signal_1432), .Q (new_AGEMA_signal_2092) ) ;
    buf_clk new_AGEMA_reg_buffer_1318 ( .C (clk), .D (keyFF_keystate_gff_17_s_next_state[1]), .Q (new_AGEMA_signal_2094) ) ;
    buf_clk new_AGEMA_reg_buffer_1320 ( .C (clk), .D (new_AGEMA_signal_1431), .Q (new_AGEMA_signal_2096) ) ;
    buf_clk new_AGEMA_reg_buffer_1322 ( .C (clk), .D (keyFF_keystate_gff_17_s_next_state[0]), .Q (new_AGEMA_signal_2098) ) ;
    buf_clk new_AGEMA_reg_buffer_1324 ( .C (clk), .D (new_AGEMA_signal_1430), .Q (new_AGEMA_signal_2100) ) ;
    buf_clk new_AGEMA_reg_buffer_1326 ( .C (clk), .D (keyFF_keystate_gff_18_s_next_state[3]), .Q (new_AGEMA_signal_2102) ) ;
    buf_clk new_AGEMA_reg_buffer_1328 ( .C (clk), .D (new_AGEMA_signal_1437), .Q (new_AGEMA_signal_2104) ) ;
    buf_clk new_AGEMA_reg_buffer_1330 ( .C (clk), .D (keyFF_keystate_gff_18_s_next_state[2]), .Q (new_AGEMA_signal_2106) ) ;
    buf_clk new_AGEMA_reg_buffer_1332 ( .C (clk), .D (new_AGEMA_signal_1436), .Q (new_AGEMA_signal_2108) ) ;
    buf_clk new_AGEMA_reg_buffer_1334 ( .C (clk), .D (keyFF_keystate_gff_18_s_next_state[1]), .Q (new_AGEMA_signal_2110) ) ;
    buf_clk new_AGEMA_reg_buffer_1336 ( .C (clk), .D (new_AGEMA_signal_1435), .Q (new_AGEMA_signal_2112) ) ;
    buf_clk new_AGEMA_reg_buffer_1338 ( .C (clk), .D (keyFF_keystate_gff_18_s_next_state[0]), .Q (new_AGEMA_signal_2114) ) ;
    buf_clk new_AGEMA_reg_buffer_1340 ( .C (clk), .D (new_AGEMA_signal_1434), .Q (new_AGEMA_signal_2116) ) ;
    buf_clk new_AGEMA_reg_buffer_1342 ( .C (clk), .D (keyFF_keystate_gff_19_s_next_state[3]), .Q (new_AGEMA_signal_2118) ) ;
    buf_clk new_AGEMA_reg_buffer_1344 ( .C (clk), .D (new_AGEMA_signal_1441), .Q (new_AGEMA_signal_2120) ) ;
    buf_clk new_AGEMA_reg_buffer_1346 ( .C (clk), .D (keyFF_keystate_gff_19_s_next_state[2]), .Q (new_AGEMA_signal_2122) ) ;
    buf_clk new_AGEMA_reg_buffer_1348 ( .C (clk), .D (new_AGEMA_signal_1440), .Q (new_AGEMA_signal_2124) ) ;
    buf_clk new_AGEMA_reg_buffer_1350 ( .C (clk), .D (keyFF_keystate_gff_19_s_next_state[1]), .Q (new_AGEMA_signal_2126) ) ;
    buf_clk new_AGEMA_reg_buffer_1352 ( .C (clk), .D (new_AGEMA_signal_1439), .Q (new_AGEMA_signal_2128) ) ;
    buf_clk new_AGEMA_reg_buffer_1354 ( .C (clk), .D (keyFF_keystate_gff_19_s_next_state[0]), .Q (new_AGEMA_signal_2130) ) ;
    buf_clk new_AGEMA_reg_buffer_1356 ( .C (clk), .D (new_AGEMA_signal_1438), .Q (new_AGEMA_signal_2132) ) ;

    /* cells in depth 2 */
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_1_MUX_inst1_mux_inst_1_U1 ( .s (new_AGEMA_signal_1498), .b ({new_AGEMA_signal_1461, serialIn[1]}), .a ({new_AGEMA_signal_1502, new_AGEMA_signal_1500}), .c ({new_AGEMA_signal_1463, stateFF_state_gff_1_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_1_MUX_inst1_mux_inst_2_U1 ( .s (new_AGEMA_signal_1498), .b ({new_AGEMA_signal_1462, serialIn[2]}), .a ({new_AGEMA_signal_1506, new_AGEMA_signal_1504}), .c ({new_AGEMA_signal_1464, stateFF_state_gff_1_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_1_MUX_inst1_mux_inst_3_U1 ( .s (new_AGEMA_signal_1498), .b ({new_AGEMA_signal_1469, serialIn[3]}), .a ({new_AGEMA_signal_1510, new_AGEMA_signal_1508}), .c ({new_AGEMA_signal_1470, stateFF_state_gff_1_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_1_U1 ( .s (new_AGEMA_signal_1511), .b ({new_AGEMA_signal_1515, new_AGEMA_signal_1513}), .a ({new_AGEMA_signal_1457, keyFF_inputPar[77]}), .c ({new_AGEMA_signal_1465, keyFF_keystate_gff_20_s_next_state[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_2_U1 ( .s (new_AGEMA_signal_1511), .b ({new_AGEMA_signal_1519, new_AGEMA_signal_1517}), .a ({new_AGEMA_signal_1459, keyFF_inputPar[78]}), .c ({new_AGEMA_signal_1466, keyFF_keystate_gff_20_s_next_state[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_20_MUX_inst1_mux_inst_3_U1 ( .s (new_AGEMA_signal_1511), .b ({new_AGEMA_signal_1523, new_AGEMA_signal_1521}), .a ({new_AGEMA_signal_1468, keyFF_inputPar[79]}), .c ({new_AGEMA_signal_1471, keyFF_keystate_gff_20_s_next_state[3]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_77_U1 ( .s (new_AGEMA_signal_1524), .b ({new_AGEMA_signal_1455, sboxOut[1]}), .a ({new_AGEMA_signal_1528, new_AGEMA_signal_1526}), .c ({new_AGEMA_signal_1457, keyFF_inputPar[77]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_78_U1 ( .s (new_AGEMA_signal_1524), .b ({new_AGEMA_signal_1454, sboxOut[2]}), .a ({new_AGEMA_signal_1532, new_AGEMA_signal_1530}), .c ({new_AGEMA_signal_1459, keyFF_inputPar[78]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) keyFF_MUX_inputPar_mux_inst_79_U1 ( .s (new_AGEMA_signal_1524), .b ({new_AGEMA_signal_1460, sboxOut[3]}), .a ({new_AGEMA_signal_1536, new_AGEMA_signal_1534}), .c ({new_AGEMA_signal_1468, keyFF_inputPar[79]}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_AND2_U1 ( .a ({new_AGEMA_signal_1444, sboxInst_Q2}), .b ({new_AGEMA_signal_1538, new_AGEMA_signal_1537}), .clk (clk), .r ({Fresh[5], Fresh[4]}), .c ({new_AGEMA_signal_1450, sboxInst_T1}) ) ;
    and_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_AND4_U1 ( .a ({new_AGEMA_signal_1449, sboxInst_Q6}), .b ({new_AGEMA_signal_1540, new_AGEMA_signal_1539}), .clk (clk), .r ({Fresh[7], Fresh[6]}), .c ({new_AGEMA_signal_1451, sboxInst_T3}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR10_U1 ( .a ({new_AGEMA_signal_1542, new_AGEMA_signal_1541}), .b ({new_AGEMA_signal_1451, sboxInst_T3}), .c ({new_AGEMA_signal_1453, sboxInst_L7}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR11_U1 ( .a ({new_AGEMA_signal_1546, new_AGEMA_signal_1544}), .b ({new_AGEMA_signal_1453, sboxInst_L7}), .c ({new_AGEMA_signal_1460, sboxOut[3]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR12_U1 ( .a ({new_AGEMA_signal_1542, new_AGEMA_signal_1541}), .b ({new_AGEMA_signal_1450, sboxInst_T1}), .c ({new_AGEMA_signal_1452, sboxInst_L8}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR13_U1 ( .a ({new_AGEMA_signal_1550, new_AGEMA_signal_1548}), .b ({new_AGEMA_signal_1452, sboxInst_L8}), .c ({new_AGEMA_signal_1454, sboxOut[2]}) ) ;
    xor_HPC3 #(.security_order(1), .pipeline(1)) sboxInst_XOR14_U1 ( .a ({new_AGEMA_signal_1552, new_AGEMA_signal_1551}), .b ({new_AGEMA_signal_1451, sboxInst_T3}), .c ({new_AGEMA_signal_1455, sboxOut[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MUX_serialIn_mux_inst_1_U1 ( .s (new_AGEMA_signal_1553), .b ({new_AGEMA_signal_1455, sboxOut[1]}), .a ({new_AGEMA_signal_1557, new_AGEMA_signal_1555}), .c ({new_AGEMA_signal_1461, serialIn[1]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MUX_serialIn_mux_inst_2_U1 ( .s (new_AGEMA_signal_1553), .b ({new_AGEMA_signal_1454, sboxOut[2]}), .a ({new_AGEMA_signal_1561, new_AGEMA_signal_1559}), .c ({new_AGEMA_signal_1462, serialIn[2]}) ) ;
    mux2_masked #(.security_order(1), .pipeline(1)) MUX_serialIn_mux_inst_3_U1 ( .s (new_AGEMA_signal_1553), .b ({new_AGEMA_signal_1460, sboxOut[3]}), .a ({new_AGEMA_signal_1565, new_AGEMA_signal_1563}), .c ({new_AGEMA_signal_1469, serialIn[3]}) ) ;
    buf_clk new_AGEMA_reg_buffer_722 ( .C (clk), .D (new_AGEMA_signal_1480), .Q (new_AGEMA_signal_1498) ) ;
    buf_clk new_AGEMA_reg_buffer_724 ( .C (clk), .D (new_AGEMA_signal_1499), .Q (new_AGEMA_signal_1500) ) ;
    buf_clk new_AGEMA_reg_buffer_726 ( .C (clk), .D (new_AGEMA_signal_1501), .Q (new_AGEMA_signal_1502) ) ;
    buf_clk new_AGEMA_reg_buffer_728 ( .C (clk), .D (new_AGEMA_signal_1503), .Q (new_AGEMA_signal_1504) ) ;
    buf_clk new_AGEMA_reg_buffer_730 ( .C (clk), .D (new_AGEMA_signal_1505), .Q (new_AGEMA_signal_1506) ) ;
    buf_clk new_AGEMA_reg_buffer_732 ( .C (clk), .D (new_AGEMA_signal_1507), .Q (new_AGEMA_signal_1508) ) ;
    buf_clk new_AGEMA_reg_buffer_734 ( .C (clk), .D (new_AGEMA_signal_1509), .Q (new_AGEMA_signal_1510) ) ;
    buf_clk new_AGEMA_reg_buffer_735 ( .C (clk), .D (new_AGEMA_signal_1483), .Q (new_AGEMA_signal_1511) ) ;
    buf_clk new_AGEMA_reg_buffer_737 ( .C (clk), .D (new_AGEMA_signal_1512), .Q (new_AGEMA_signal_1513) ) ;
    buf_clk new_AGEMA_reg_buffer_739 ( .C (clk), .D (new_AGEMA_signal_1514), .Q (new_AGEMA_signal_1515) ) ;
    buf_clk new_AGEMA_reg_buffer_741 ( .C (clk), .D (new_AGEMA_signal_1516), .Q (new_AGEMA_signal_1517) ) ;
    buf_clk new_AGEMA_reg_buffer_743 ( .C (clk), .D (new_AGEMA_signal_1518), .Q (new_AGEMA_signal_1519) ) ;
    buf_clk new_AGEMA_reg_buffer_745 ( .C (clk), .D (new_AGEMA_signal_1520), .Q (new_AGEMA_signal_1521) ) ;
    buf_clk new_AGEMA_reg_buffer_747 ( .C (clk), .D (new_AGEMA_signal_1522), .Q (new_AGEMA_signal_1523) ) ;
    buf_clk new_AGEMA_reg_buffer_748 ( .C (clk), .D (new_AGEMA_signal_1486), .Q (new_AGEMA_signal_1524) ) ;
    buf_clk new_AGEMA_reg_buffer_750 ( .C (clk), .D (new_AGEMA_signal_1525), .Q (new_AGEMA_signal_1526) ) ;
    buf_clk new_AGEMA_reg_buffer_752 ( .C (clk), .D (new_AGEMA_signal_1527), .Q (new_AGEMA_signal_1528) ) ;
    buf_clk new_AGEMA_reg_buffer_754 ( .C (clk), .D (new_AGEMA_signal_1529), .Q (new_AGEMA_signal_1530) ) ;
    buf_clk new_AGEMA_reg_buffer_756 ( .C (clk), .D (new_AGEMA_signal_1531), .Q (new_AGEMA_signal_1532) ) ;
    buf_clk new_AGEMA_reg_buffer_758 ( .C (clk), .D (new_AGEMA_signal_1533), .Q (new_AGEMA_signal_1534) ) ;
    buf_clk new_AGEMA_reg_buffer_760 ( .C (clk), .D (new_AGEMA_signal_1535), .Q (new_AGEMA_signal_1536) ) ;
    buf_clk new_AGEMA_reg_buffer_765 ( .C (clk), .D (sboxInst_L5), .Q (new_AGEMA_signal_1541) ) ;
    buf_clk new_AGEMA_reg_buffer_766 ( .C (clk), .D (new_AGEMA_signal_1445), .Q (new_AGEMA_signal_1542) ) ;
    buf_clk new_AGEMA_reg_buffer_768 ( .C (clk), .D (new_AGEMA_signal_1543), .Q (new_AGEMA_signal_1544) ) ;
    buf_clk new_AGEMA_reg_buffer_770 ( .C (clk), .D (new_AGEMA_signal_1545), .Q (new_AGEMA_signal_1546) ) ;
    buf_clk new_AGEMA_reg_buffer_772 ( .C (clk), .D (new_AGEMA_signal_1547), .Q (new_AGEMA_signal_1548) ) ;
    buf_clk new_AGEMA_reg_buffer_774 ( .C (clk), .D (new_AGEMA_signal_1549), .Q (new_AGEMA_signal_1550) ) ;
    buf_clk new_AGEMA_reg_buffer_775 ( .C (clk), .D (new_AGEMA_signal_1491), .Q (new_AGEMA_signal_1551) ) ;
    buf_clk new_AGEMA_reg_buffer_776 ( .C (clk), .D (new_AGEMA_signal_1492), .Q (new_AGEMA_signal_1552) ) ;
    buf_clk new_AGEMA_reg_buffer_777 ( .C (clk), .D (new_AGEMA_signal_1495), .Q (new_AGEMA_signal_1553) ) ;
    buf_clk new_AGEMA_reg_buffer_779 ( .C (clk), .D (new_AGEMA_signal_1554), .Q (new_AGEMA_signal_1555) ) ;
    buf_clk new_AGEMA_reg_buffer_781 ( .C (clk), .D (new_AGEMA_signal_1556), .Q (new_AGEMA_signal_1557) ) ;
    buf_clk new_AGEMA_reg_buffer_783 ( .C (clk), .D (new_AGEMA_signal_1558), .Q (new_AGEMA_signal_1559) ) ;
    buf_clk new_AGEMA_reg_buffer_785 ( .C (clk), .D (new_AGEMA_signal_1560), .Q (new_AGEMA_signal_1561) ) ;
    buf_clk new_AGEMA_reg_buffer_787 ( .C (clk), .D (new_AGEMA_signal_1562), .Q (new_AGEMA_signal_1563) ) ;
    buf_clk new_AGEMA_reg_buffer_789 ( .C (clk), .D (new_AGEMA_signal_1564), .Q (new_AGEMA_signal_1565) ) ;
    buf_clk new_AGEMA_reg_buffer_791 ( .C (clk), .D (new_AGEMA_signal_1566), .Q (new_AGEMA_signal_1567) ) ;
    buf_clk new_AGEMA_reg_buffer_793 ( .C (clk), .D (new_AGEMA_signal_1568), .Q (new_AGEMA_signal_1569) ) ;
    buf_clk new_AGEMA_reg_buffer_795 ( .C (clk), .D (new_AGEMA_signal_1570), .Q (new_AGEMA_signal_1571) ) ;
    buf_clk new_AGEMA_reg_buffer_797 ( .C (clk), .D (new_AGEMA_signal_1572), .Q (new_AGEMA_signal_1573) ) ;
    buf_clk new_AGEMA_reg_buffer_799 ( .C (clk), .D (new_AGEMA_signal_1574), .Q (new_AGEMA_signal_1575) ) ;
    buf_clk new_AGEMA_reg_buffer_801 ( .C (clk), .D (new_AGEMA_signal_1576), .Q (new_AGEMA_signal_1577) ) ;
    buf_clk new_AGEMA_reg_buffer_803 ( .C (clk), .D (new_AGEMA_signal_1578), .Q (new_AGEMA_signal_1579) ) ;
    buf_clk new_AGEMA_reg_buffer_805 ( .C (clk), .D (new_AGEMA_signal_1580), .Q (new_AGEMA_signal_1581) ) ;
    buf_clk new_AGEMA_reg_buffer_807 ( .C (clk), .D (new_AGEMA_signal_1582), .Q (new_AGEMA_signal_1583) ) ;
    buf_clk new_AGEMA_reg_buffer_809 ( .C (clk), .D (new_AGEMA_signal_1584), .Q (new_AGEMA_signal_1585) ) ;
    buf_clk new_AGEMA_reg_buffer_811 ( .C (clk), .D (new_AGEMA_signal_1586), .Q (new_AGEMA_signal_1587) ) ;
    buf_clk new_AGEMA_reg_buffer_812 ( .C (clk), .D (stateFF_state_gff_1_s_next_state[0]), .Q (new_AGEMA_signal_1588) ) ;
    buf_clk new_AGEMA_reg_buffer_813 ( .C (clk), .D (new_AGEMA_signal_1447), .Q (new_AGEMA_signal_1589) ) ;
    buf_clk new_AGEMA_reg_buffer_815 ( .C (clk), .D (new_AGEMA_signal_1590), .Q (new_AGEMA_signal_1591) ) ;
    buf_clk new_AGEMA_reg_buffer_817 ( .C (clk), .D (new_AGEMA_signal_1592), .Q (new_AGEMA_signal_1593) ) ;
    buf_clk new_AGEMA_reg_buffer_819 ( .C (clk), .D (new_AGEMA_signal_1594), .Q (new_AGEMA_signal_1595) ) ;
    buf_clk new_AGEMA_reg_buffer_821 ( .C (clk), .D (new_AGEMA_signal_1596), .Q (new_AGEMA_signal_1597) ) ;
    buf_clk new_AGEMA_reg_buffer_823 ( .C (clk), .D (new_AGEMA_signal_1598), .Q (new_AGEMA_signal_1599) ) ;
    buf_clk new_AGEMA_reg_buffer_825 ( .C (clk), .D (new_AGEMA_signal_1600), .Q (new_AGEMA_signal_1601) ) ;
    buf_clk new_AGEMA_reg_buffer_827 ( .C (clk), .D (new_AGEMA_signal_1602), .Q (new_AGEMA_signal_1603) ) ;
    buf_clk new_AGEMA_reg_buffer_829 ( .C (clk), .D (new_AGEMA_signal_1604), .Q (new_AGEMA_signal_1605) ) ;
    buf_clk new_AGEMA_reg_buffer_831 ( .C (clk), .D (new_AGEMA_signal_1606), .Q (new_AGEMA_signal_1607) ) ;
    buf_clk new_AGEMA_reg_buffer_833 ( .C (clk), .D (new_AGEMA_signal_1608), .Q (new_AGEMA_signal_1609) ) ;
    buf_clk new_AGEMA_reg_buffer_835 ( .C (clk), .D (new_AGEMA_signal_1610), .Q (new_AGEMA_signal_1611) ) ;
    buf_clk new_AGEMA_reg_buffer_837 ( .C (clk), .D (new_AGEMA_signal_1612), .Q (new_AGEMA_signal_1613) ) ;
    buf_clk new_AGEMA_reg_buffer_839 ( .C (clk), .D (new_AGEMA_signal_1614), .Q (new_AGEMA_signal_1615) ) ;
    buf_clk new_AGEMA_reg_buffer_841 ( .C (clk), .D (new_AGEMA_signal_1616), .Q (new_AGEMA_signal_1617) ) ;
    buf_clk new_AGEMA_reg_buffer_843 ( .C (clk), .D (new_AGEMA_signal_1618), .Q (new_AGEMA_signal_1619) ) ;
    buf_clk new_AGEMA_reg_buffer_845 ( .C (clk), .D (new_AGEMA_signal_1620), .Q (new_AGEMA_signal_1621) ) ;
    buf_clk new_AGEMA_reg_buffer_847 ( .C (clk), .D (new_AGEMA_signal_1622), .Q (new_AGEMA_signal_1623) ) ;
    buf_clk new_AGEMA_reg_buffer_849 ( .C (clk), .D (new_AGEMA_signal_1624), .Q (new_AGEMA_signal_1625) ) ;
    buf_clk new_AGEMA_reg_buffer_851 ( .C (clk), .D (new_AGEMA_signal_1626), .Q (new_AGEMA_signal_1627) ) ;
    buf_clk new_AGEMA_reg_buffer_853 ( .C (clk), .D (new_AGEMA_signal_1628), .Q (new_AGEMA_signal_1629) ) ;
    buf_clk new_AGEMA_reg_buffer_855 ( .C (clk), .D (new_AGEMA_signal_1630), .Q (new_AGEMA_signal_1631) ) ;
    buf_clk new_AGEMA_reg_buffer_857 ( .C (clk), .D (new_AGEMA_signal_1632), .Q (new_AGEMA_signal_1633) ) ;
    buf_clk new_AGEMA_reg_buffer_859 ( .C (clk), .D (new_AGEMA_signal_1634), .Q (new_AGEMA_signal_1635) ) ;
    buf_clk new_AGEMA_reg_buffer_861 ( .C (clk), .D (new_AGEMA_signal_1636), .Q (new_AGEMA_signal_1637) ) ;
    buf_clk new_AGEMA_reg_buffer_863 ( .C (clk), .D (new_AGEMA_signal_1638), .Q (new_AGEMA_signal_1639) ) ;
    buf_clk new_AGEMA_reg_buffer_865 ( .C (clk), .D (new_AGEMA_signal_1640), .Q (new_AGEMA_signal_1641) ) ;
    buf_clk new_AGEMA_reg_buffer_867 ( .C (clk), .D (new_AGEMA_signal_1642), .Q (new_AGEMA_signal_1643) ) ;
    buf_clk new_AGEMA_reg_buffer_869 ( .C (clk), .D (new_AGEMA_signal_1644), .Q (new_AGEMA_signal_1645) ) ;
    buf_clk new_AGEMA_reg_buffer_871 ( .C (clk), .D (new_AGEMA_signal_1646), .Q (new_AGEMA_signal_1647) ) ;
    buf_clk new_AGEMA_reg_buffer_873 ( .C (clk), .D (new_AGEMA_signal_1648), .Q (new_AGEMA_signal_1649) ) ;
    buf_clk new_AGEMA_reg_buffer_875 ( .C (clk), .D (new_AGEMA_signal_1650), .Q (new_AGEMA_signal_1651) ) ;
    buf_clk new_AGEMA_reg_buffer_877 ( .C (clk), .D (new_AGEMA_signal_1652), .Q (new_AGEMA_signal_1653) ) ;
    buf_clk new_AGEMA_reg_buffer_879 ( .C (clk), .D (new_AGEMA_signal_1654), .Q (new_AGEMA_signal_1655) ) ;
    buf_clk new_AGEMA_reg_buffer_881 ( .C (clk), .D (new_AGEMA_signal_1656), .Q (new_AGEMA_signal_1657) ) ;
    buf_clk new_AGEMA_reg_buffer_883 ( .C (clk), .D (new_AGEMA_signal_1658), .Q (new_AGEMA_signal_1659) ) ;
    buf_clk new_AGEMA_reg_buffer_885 ( .C (clk), .D (new_AGEMA_signal_1660), .Q (new_AGEMA_signal_1661) ) ;
    buf_clk new_AGEMA_reg_buffer_887 ( .C (clk), .D (new_AGEMA_signal_1662), .Q (new_AGEMA_signal_1663) ) ;
    buf_clk new_AGEMA_reg_buffer_889 ( .C (clk), .D (new_AGEMA_signal_1664), .Q (new_AGEMA_signal_1665) ) ;
    buf_clk new_AGEMA_reg_buffer_891 ( .C (clk), .D (new_AGEMA_signal_1666), .Q (new_AGEMA_signal_1667) ) ;
    buf_clk new_AGEMA_reg_buffer_893 ( .C (clk), .D (new_AGEMA_signal_1668), .Q (new_AGEMA_signal_1669) ) ;
    buf_clk new_AGEMA_reg_buffer_895 ( .C (clk), .D (new_AGEMA_signal_1670), .Q (new_AGEMA_signal_1671) ) ;
    buf_clk new_AGEMA_reg_buffer_897 ( .C (clk), .D (new_AGEMA_signal_1672), .Q (new_AGEMA_signal_1673) ) ;
    buf_clk new_AGEMA_reg_buffer_899 ( .C (clk), .D (new_AGEMA_signal_1674), .Q (new_AGEMA_signal_1675) ) ;
    buf_clk new_AGEMA_reg_buffer_901 ( .C (clk), .D (new_AGEMA_signal_1676), .Q (new_AGEMA_signal_1677) ) ;
    buf_clk new_AGEMA_reg_buffer_903 ( .C (clk), .D (new_AGEMA_signal_1678), .Q (new_AGEMA_signal_1679) ) ;
    buf_clk new_AGEMA_reg_buffer_905 ( .C (clk), .D (new_AGEMA_signal_1680), .Q (new_AGEMA_signal_1681) ) ;
    buf_clk new_AGEMA_reg_buffer_907 ( .C (clk), .D (new_AGEMA_signal_1682), .Q (new_AGEMA_signal_1683) ) ;
    buf_clk new_AGEMA_reg_buffer_909 ( .C (clk), .D (new_AGEMA_signal_1684), .Q (new_AGEMA_signal_1685) ) ;
    buf_clk new_AGEMA_reg_buffer_911 ( .C (clk), .D (new_AGEMA_signal_1686), .Q (new_AGEMA_signal_1687) ) ;
    buf_clk new_AGEMA_reg_buffer_913 ( .C (clk), .D (new_AGEMA_signal_1688), .Q (new_AGEMA_signal_1689) ) ;
    buf_clk new_AGEMA_reg_buffer_915 ( .C (clk), .D (new_AGEMA_signal_1690), .Q (new_AGEMA_signal_1691) ) ;
    buf_clk new_AGEMA_reg_buffer_917 ( .C (clk), .D (new_AGEMA_signal_1692), .Q (new_AGEMA_signal_1693) ) ;
    buf_clk new_AGEMA_reg_buffer_919 ( .C (clk), .D (new_AGEMA_signal_1694), .Q (new_AGEMA_signal_1695) ) ;
    buf_clk new_AGEMA_reg_buffer_921 ( .C (clk), .D (new_AGEMA_signal_1696), .Q (new_AGEMA_signal_1697) ) ;
    buf_clk new_AGEMA_reg_buffer_923 ( .C (clk), .D (new_AGEMA_signal_1698), .Q (new_AGEMA_signal_1699) ) ;
    buf_clk new_AGEMA_reg_buffer_925 ( .C (clk), .D (new_AGEMA_signal_1700), .Q (new_AGEMA_signal_1701) ) ;
    buf_clk new_AGEMA_reg_buffer_927 ( .C (clk), .D (new_AGEMA_signal_1702), .Q (new_AGEMA_signal_1703) ) ;
    buf_clk new_AGEMA_reg_buffer_929 ( .C (clk), .D (new_AGEMA_signal_1704), .Q (new_AGEMA_signal_1705) ) ;
    buf_clk new_AGEMA_reg_buffer_931 ( .C (clk), .D (new_AGEMA_signal_1706), .Q (new_AGEMA_signal_1707) ) ;
    buf_clk new_AGEMA_reg_buffer_933 ( .C (clk), .D (new_AGEMA_signal_1708), .Q (new_AGEMA_signal_1709) ) ;
    buf_clk new_AGEMA_reg_buffer_935 ( .C (clk), .D (new_AGEMA_signal_1710), .Q (new_AGEMA_signal_1711) ) ;
    buf_clk new_AGEMA_reg_buffer_937 ( .C (clk), .D (new_AGEMA_signal_1712), .Q (new_AGEMA_signal_1713) ) ;
    buf_clk new_AGEMA_reg_buffer_939 ( .C (clk), .D (new_AGEMA_signal_1714), .Q (new_AGEMA_signal_1715) ) ;
    buf_clk new_AGEMA_reg_buffer_941 ( .C (clk), .D (new_AGEMA_signal_1716), .Q (new_AGEMA_signal_1717) ) ;
    buf_clk new_AGEMA_reg_buffer_943 ( .C (clk), .D (new_AGEMA_signal_1718), .Q (new_AGEMA_signal_1719) ) ;
    buf_clk new_AGEMA_reg_buffer_945 ( .C (clk), .D (new_AGEMA_signal_1720), .Q (new_AGEMA_signal_1721) ) ;
    buf_clk new_AGEMA_reg_buffer_947 ( .C (clk), .D (new_AGEMA_signal_1722), .Q (new_AGEMA_signal_1723) ) ;
    buf_clk new_AGEMA_reg_buffer_949 ( .C (clk), .D (new_AGEMA_signal_1724), .Q (new_AGEMA_signal_1725) ) ;
    buf_clk new_AGEMA_reg_buffer_951 ( .C (clk), .D (new_AGEMA_signal_1726), .Q (new_AGEMA_signal_1727) ) ;
    buf_clk new_AGEMA_reg_buffer_953 ( .C (clk), .D (new_AGEMA_signal_1728), .Q (new_AGEMA_signal_1729) ) ;
    buf_clk new_AGEMA_reg_buffer_955 ( .C (clk), .D (new_AGEMA_signal_1730), .Q (new_AGEMA_signal_1731) ) ;
    buf_clk new_AGEMA_reg_buffer_957 ( .C (clk), .D (new_AGEMA_signal_1732), .Q (new_AGEMA_signal_1733) ) ;
    buf_clk new_AGEMA_reg_buffer_959 ( .C (clk), .D (new_AGEMA_signal_1734), .Q (new_AGEMA_signal_1735) ) ;
    buf_clk new_AGEMA_reg_buffer_961 ( .C (clk), .D (new_AGEMA_signal_1736), .Q (new_AGEMA_signal_1737) ) ;
    buf_clk new_AGEMA_reg_buffer_963 ( .C (clk), .D (new_AGEMA_signal_1738), .Q (new_AGEMA_signal_1739) ) ;
    buf_clk new_AGEMA_reg_buffer_965 ( .C (clk), .D (new_AGEMA_signal_1740), .Q (new_AGEMA_signal_1741) ) ;
    buf_clk new_AGEMA_reg_buffer_967 ( .C (clk), .D (new_AGEMA_signal_1742), .Q (new_AGEMA_signal_1743) ) ;
    buf_clk new_AGEMA_reg_buffer_969 ( .C (clk), .D (new_AGEMA_signal_1744), .Q (new_AGEMA_signal_1745) ) ;
    buf_clk new_AGEMA_reg_buffer_971 ( .C (clk), .D (new_AGEMA_signal_1746), .Q (new_AGEMA_signal_1747) ) ;
    buf_clk new_AGEMA_reg_buffer_973 ( .C (clk), .D (new_AGEMA_signal_1748), .Q (new_AGEMA_signal_1749) ) ;
    buf_clk new_AGEMA_reg_buffer_975 ( .C (clk), .D (new_AGEMA_signal_1750), .Q (new_AGEMA_signal_1751) ) ;
    buf_clk new_AGEMA_reg_buffer_977 ( .C (clk), .D (new_AGEMA_signal_1752), .Q (new_AGEMA_signal_1753) ) ;
    buf_clk new_AGEMA_reg_buffer_979 ( .C (clk), .D (new_AGEMA_signal_1754), .Q (new_AGEMA_signal_1755) ) ;
    buf_clk new_AGEMA_reg_buffer_981 ( .C (clk), .D (new_AGEMA_signal_1756), .Q (new_AGEMA_signal_1757) ) ;
    buf_clk new_AGEMA_reg_buffer_983 ( .C (clk), .D (new_AGEMA_signal_1758), .Q (new_AGEMA_signal_1759) ) ;
    buf_clk new_AGEMA_reg_buffer_985 ( .C (clk), .D (new_AGEMA_signal_1760), .Q (new_AGEMA_signal_1761) ) ;
    buf_clk new_AGEMA_reg_buffer_987 ( .C (clk), .D (new_AGEMA_signal_1762), .Q (new_AGEMA_signal_1763) ) ;
    buf_clk new_AGEMA_reg_buffer_989 ( .C (clk), .D (new_AGEMA_signal_1764), .Q (new_AGEMA_signal_1765) ) ;
    buf_clk new_AGEMA_reg_buffer_991 ( .C (clk), .D (new_AGEMA_signal_1766), .Q (new_AGEMA_signal_1767) ) ;
    buf_clk new_AGEMA_reg_buffer_993 ( .C (clk), .D (new_AGEMA_signal_1768), .Q (new_AGEMA_signal_1769) ) ;
    buf_clk new_AGEMA_reg_buffer_995 ( .C (clk), .D (new_AGEMA_signal_1770), .Q (new_AGEMA_signal_1771) ) ;
    buf_clk new_AGEMA_reg_buffer_997 ( .C (clk), .D (new_AGEMA_signal_1772), .Q (new_AGEMA_signal_1773) ) ;
    buf_clk new_AGEMA_reg_buffer_999 ( .C (clk), .D (new_AGEMA_signal_1774), .Q (new_AGEMA_signal_1775) ) ;
    buf_clk new_AGEMA_reg_buffer_1001 ( .C (clk), .D (new_AGEMA_signal_1776), .Q (new_AGEMA_signal_1777) ) ;
    buf_clk new_AGEMA_reg_buffer_1003 ( .C (clk), .D (new_AGEMA_signal_1778), .Q (new_AGEMA_signal_1779) ) ;
    buf_clk new_AGEMA_reg_buffer_1005 ( .C (clk), .D (new_AGEMA_signal_1780), .Q (new_AGEMA_signal_1781) ) ;
    buf_clk new_AGEMA_reg_buffer_1007 ( .C (clk), .D (new_AGEMA_signal_1782), .Q (new_AGEMA_signal_1783) ) ;
    buf_clk new_AGEMA_reg_buffer_1009 ( .C (clk), .D (new_AGEMA_signal_1784), .Q (new_AGEMA_signal_1785) ) ;
    buf_clk new_AGEMA_reg_buffer_1011 ( .C (clk), .D (new_AGEMA_signal_1786), .Q (new_AGEMA_signal_1787) ) ;
    buf_clk new_AGEMA_reg_buffer_1013 ( .C (clk), .D (new_AGEMA_signal_1788), .Q (new_AGEMA_signal_1789) ) ;
    buf_clk new_AGEMA_reg_buffer_1015 ( .C (clk), .D (new_AGEMA_signal_1790), .Q (new_AGEMA_signal_1791) ) ;
    buf_clk new_AGEMA_reg_buffer_1017 ( .C (clk), .D (new_AGEMA_signal_1792), .Q (new_AGEMA_signal_1793) ) ;
    buf_clk new_AGEMA_reg_buffer_1019 ( .C (clk), .D (new_AGEMA_signal_1794), .Q (new_AGEMA_signal_1795) ) ;
    buf_clk new_AGEMA_reg_buffer_1021 ( .C (clk), .D (new_AGEMA_signal_1796), .Q (new_AGEMA_signal_1797) ) ;
    buf_clk new_AGEMA_reg_buffer_1023 ( .C (clk), .D (new_AGEMA_signal_1798), .Q (new_AGEMA_signal_1799) ) ;
    buf_clk new_AGEMA_reg_buffer_1025 ( .C (clk), .D (new_AGEMA_signal_1800), .Q (new_AGEMA_signal_1801) ) ;
    buf_clk new_AGEMA_reg_buffer_1027 ( .C (clk), .D (new_AGEMA_signal_1802), .Q (new_AGEMA_signal_1803) ) ;
    buf_clk new_AGEMA_reg_buffer_1029 ( .C (clk), .D (new_AGEMA_signal_1804), .Q (new_AGEMA_signal_1805) ) ;
    buf_clk new_AGEMA_reg_buffer_1031 ( .C (clk), .D (new_AGEMA_signal_1806), .Q (new_AGEMA_signal_1807) ) ;
    buf_clk new_AGEMA_reg_buffer_1033 ( .C (clk), .D (new_AGEMA_signal_1808), .Q (new_AGEMA_signal_1809) ) ;
    buf_clk new_AGEMA_reg_buffer_1035 ( .C (clk), .D (new_AGEMA_signal_1810), .Q (new_AGEMA_signal_1811) ) ;
    buf_clk new_AGEMA_reg_buffer_1037 ( .C (clk), .D (new_AGEMA_signal_1812), .Q (new_AGEMA_signal_1813) ) ;
    buf_clk new_AGEMA_reg_buffer_1039 ( .C (clk), .D (new_AGEMA_signal_1814), .Q (new_AGEMA_signal_1815) ) ;
    buf_clk new_AGEMA_reg_buffer_1041 ( .C (clk), .D (new_AGEMA_signal_1816), .Q (new_AGEMA_signal_1817) ) ;
    buf_clk new_AGEMA_reg_buffer_1043 ( .C (clk), .D (new_AGEMA_signal_1818), .Q (new_AGEMA_signal_1819) ) ;
    buf_clk new_AGEMA_reg_buffer_1045 ( .C (clk), .D (new_AGEMA_signal_1820), .Q (new_AGEMA_signal_1821) ) ;
    buf_clk new_AGEMA_reg_buffer_1047 ( .C (clk), .D (new_AGEMA_signal_1822), .Q (new_AGEMA_signal_1823) ) ;
    buf_clk new_AGEMA_reg_buffer_1049 ( .C (clk), .D (new_AGEMA_signal_1824), .Q (new_AGEMA_signal_1825) ) ;
    buf_clk new_AGEMA_reg_buffer_1051 ( .C (clk), .D (new_AGEMA_signal_1826), .Q (new_AGEMA_signal_1827) ) ;
    buf_clk new_AGEMA_reg_buffer_1053 ( .C (clk), .D (new_AGEMA_signal_1828), .Q (new_AGEMA_signal_1829) ) ;
    buf_clk new_AGEMA_reg_buffer_1055 ( .C (clk), .D (new_AGEMA_signal_1830), .Q (new_AGEMA_signal_1831) ) ;
    buf_clk new_AGEMA_reg_buffer_1057 ( .C (clk), .D (new_AGEMA_signal_1832), .Q (new_AGEMA_signal_1833) ) ;
    buf_clk new_AGEMA_reg_buffer_1059 ( .C (clk), .D (new_AGEMA_signal_1834), .Q (new_AGEMA_signal_1835) ) ;
    buf_clk new_AGEMA_reg_buffer_1061 ( .C (clk), .D (new_AGEMA_signal_1836), .Q (new_AGEMA_signal_1837) ) ;
    buf_clk new_AGEMA_reg_buffer_1063 ( .C (clk), .D (new_AGEMA_signal_1838), .Q (new_AGEMA_signal_1839) ) ;
    buf_clk new_AGEMA_reg_buffer_1065 ( .C (clk), .D (new_AGEMA_signal_1840), .Q (new_AGEMA_signal_1841) ) ;
    buf_clk new_AGEMA_reg_buffer_1067 ( .C (clk), .D (new_AGEMA_signal_1842), .Q (new_AGEMA_signal_1843) ) ;
    buf_clk new_AGEMA_reg_buffer_1069 ( .C (clk), .D (new_AGEMA_signal_1844), .Q (new_AGEMA_signal_1845) ) ;
    buf_clk new_AGEMA_reg_buffer_1071 ( .C (clk), .D (new_AGEMA_signal_1846), .Q (new_AGEMA_signal_1847) ) ;
    buf_clk new_AGEMA_reg_buffer_1073 ( .C (clk), .D (new_AGEMA_signal_1848), .Q (new_AGEMA_signal_1849) ) ;
    buf_clk new_AGEMA_reg_buffer_1075 ( .C (clk), .D (new_AGEMA_signal_1850), .Q (new_AGEMA_signal_1851) ) ;
    buf_clk new_AGEMA_reg_buffer_1077 ( .C (clk), .D (new_AGEMA_signal_1852), .Q (new_AGEMA_signal_1853) ) ;
    buf_clk new_AGEMA_reg_buffer_1079 ( .C (clk), .D (new_AGEMA_signal_1854), .Q (new_AGEMA_signal_1855) ) ;
    buf_clk new_AGEMA_reg_buffer_1081 ( .C (clk), .D (new_AGEMA_signal_1856), .Q (new_AGEMA_signal_1857) ) ;
    buf_clk new_AGEMA_reg_buffer_1083 ( .C (clk), .D (new_AGEMA_signal_1858), .Q (new_AGEMA_signal_1859) ) ;
    buf_clk new_AGEMA_reg_buffer_1085 ( .C (clk), .D (new_AGEMA_signal_1860), .Q (new_AGEMA_signal_1861) ) ;
    buf_clk new_AGEMA_reg_buffer_1087 ( .C (clk), .D (new_AGEMA_signal_1862), .Q (new_AGEMA_signal_1863) ) ;
    buf_clk new_AGEMA_reg_buffer_1089 ( .C (clk), .D (new_AGEMA_signal_1864), .Q (new_AGEMA_signal_1865) ) ;
    buf_clk new_AGEMA_reg_buffer_1091 ( .C (clk), .D (new_AGEMA_signal_1866), .Q (new_AGEMA_signal_1867) ) ;
    buf_clk new_AGEMA_reg_buffer_1093 ( .C (clk), .D (new_AGEMA_signal_1868), .Q (new_AGEMA_signal_1869) ) ;
    buf_clk new_AGEMA_reg_buffer_1095 ( .C (clk), .D (new_AGEMA_signal_1870), .Q (new_AGEMA_signal_1871) ) ;
    buf_clk new_AGEMA_reg_buffer_1097 ( .C (clk), .D (new_AGEMA_signal_1872), .Q (new_AGEMA_signal_1873) ) ;
    buf_clk new_AGEMA_reg_buffer_1099 ( .C (clk), .D (new_AGEMA_signal_1874), .Q (new_AGEMA_signal_1875) ) ;
    buf_clk new_AGEMA_reg_buffer_1101 ( .C (clk), .D (new_AGEMA_signal_1876), .Q (new_AGEMA_signal_1877) ) ;
    buf_clk new_AGEMA_reg_buffer_1103 ( .C (clk), .D (new_AGEMA_signal_1878), .Q (new_AGEMA_signal_1879) ) ;
    buf_clk new_AGEMA_reg_buffer_1105 ( .C (clk), .D (new_AGEMA_signal_1880), .Q (new_AGEMA_signal_1881) ) ;
    buf_clk new_AGEMA_reg_buffer_1107 ( .C (clk), .D (new_AGEMA_signal_1882), .Q (new_AGEMA_signal_1883) ) ;
    buf_clk new_AGEMA_reg_buffer_1109 ( .C (clk), .D (new_AGEMA_signal_1884), .Q (new_AGEMA_signal_1885) ) ;
    buf_clk new_AGEMA_reg_buffer_1111 ( .C (clk), .D (new_AGEMA_signal_1886), .Q (new_AGEMA_signal_1887) ) ;
    buf_clk new_AGEMA_reg_buffer_1113 ( .C (clk), .D (new_AGEMA_signal_1888), .Q (new_AGEMA_signal_1889) ) ;
    buf_clk new_AGEMA_reg_buffer_1115 ( .C (clk), .D (new_AGEMA_signal_1890), .Q (new_AGEMA_signal_1891) ) ;
    buf_clk new_AGEMA_reg_buffer_1117 ( .C (clk), .D (new_AGEMA_signal_1892), .Q (new_AGEMA_signal_1893) ) ;
    buf_clk new_AGEMA_reg_buffer_1119 ( .C (clk), .D (new_AGEMA_signal_1894), .Q (new_AGEMA_signal_1895) ) ;
    buf_clk new_AGEMA_reg_buffer_1121 ( .C (clk), .D (new_AGEMA_signal_1896), .Q (new_AGEMA_signal_1897) ) ;
    buf_clk new_AGEMA_reg_buffer_1123 ( .C (clk), .D (new_AGEMA_signal_1898), .Q (new_AGEMA_signal_1899) ) ;
    buf_clk new_AGEMA_reg_buffer_1125 ( .C (clk), .D (new_AGEMA_signal_1900), .Q (new_AGEMA_signal_1901) ) ;
    buf_clk new_AGEMA_reg_buffer_1127 ( .C (clk), .D (new_AGEMA_signal_1902), .Q (new_AGEMA_signal_1903) ) ;
    buf_clk new_AGEMA_reg_buffer_1129 ( .C (clk), .D (new_AGEMA_signal_1904), .Q (new_AGEMA_signal_1905) ) ;
    buf_clk new_AGEMA_reg_buffer_1131 ( .C (clk), .D (new_AGEMA_signal_1906), .Q (new_AGEMA_signal_1907) ) ;
    buf_clk new_AGEMA_reg_buffer_1133 ( .C (clk), .D (new_AGEMA_signal_1908), .Q (new_AGEMA_signal_1909) ) ;
    buf_clk new_AGEMA_reg_buffer_1135 ( .C (clk), .D (new_AGEMA_signal_1910), .Q (new_AGEMA_signal_1911) ) ;
    buf_clk new_AGEMA_reg_buffer_1137 ( .C (clk), .D (new_AGEMA_signal_1912), .Q (new_AGEMA_signal_1913) ) ;
    buf_clk new_AGEMA_reg_buffer_1139 ( .C (clk), .D (new_AGEMA_signal_1914), .Q (new_AGEMA_signal_1915) ) ;
    buf_clk new_AGEMA_reg_buffer_1141 ( .C (clk), .D (new_AGEMA_signal_1916), .Q (new_AGEMA_signal_1917) ) ;
    buf_clk new_AGEMA_reg_buffer_1143 ( .C (clk), .D (new_AGEMA_signal_1918), .Q (new_AGEMA_signal_1919) ) ;
    buf_clk new_AGEMA_reg_buffer_1145 ( .C (clk), .D (new_AGEMA_signal_1920), .Q (new_AGEMA_signal_1921) ) ;
    buf_clk new_AGEMA_reg_buffer_1147 ( .C (clk), .D (new_AGEMA_signal_1922), .Q (new_AGEMA_signal_1923) ) ;
    buf_clk new_AGEMA_reg_buffer_1149 ( .C (clk), .D (new_AGEMA_signal_1924), .Q (new_AGEMA_signal_1925) ) ;
    buf_clk new_AGEMA_reg_buffer_1151 ( .C (clk), .D (new_AGEMA_signal_1926), .Q (new_AGEMA_signal_1927) ) ;
    buf_clk new_AGEMA_reg_buffer_1153 ( .C (clk), .D (new_AGEMA_signal_1928), .Q (new_AGEMA_signal_1929) ) ;
    buf_clk new_AGEMA_reg_buffer_1155 ( .C (clk), .D (new_AGEMA_signal_1930), .Q (new_AGEMA_signal_1931) ) ;
    buf_clk new_AGEMA_reg_buffer_1157 ( .C (clk), .D (new_AGEMA_signal_1932), .Q (new_AGEMA_signal_1933) ) ;
    buf_clk new_AGEMA_reg_buffer_1159 ( .C (clk), .D (new_AGEMA_signal_1934), .Q (new_AGEMA_signal_1935) ) ;
    buf_clk new_AGEMA_reg_buffer_1161 ( .C (clk), .D (new_AGEMA_signal_1936), .Q (new_AGEMA_signal_1937) ) ;
    buf_clk new_AGEMA_reg_buffer_1163 ( .C (clk), .D (new_AGEMA_signal_1938), .Q (new_AGEMA_signal_1939) ) ;
    buf_clk new_AGEMA_reg_buffer_1165 ( .C (clk), .D (new_AGEMA_signal_1940), .Q (new_AGEMA_signal_1941) ) ;
    buf_clk new_AGEMA_reg_buffer_1167 ( .C (clk), .D (new_AGEMA_signal_1942), .Q (new_AGEMA_signal_1943) ) ;
    buf_clk new_AGEMA_reg_buffer_1169 ( .C (clk), .D (new_AGEMA_signal_1944), .Q (new_AGEMA_signal_1945) ) ;
    buf_clk new_AGEMA_reg_buffer_1171 ( .C (clk), .D (new_AGEMA_signal_1946), .Q (new_AGEMA_signal_1947) ) ;
    buf_clk new_AGEMA_reg_buffer_1173 ( .C (clk), .D (new_AGEMA_signal_1948), .Q (new_AGEMA_signal_1949) ) ;
    buf_clk new_AGEMA_reg_buffer_1175 ( .C (clk), .D (new_AGEMA_signal_1950), .Q (new_AGEMA_signal_1951) ) ;
    buf_clk new_AGEMA_reg_buffer_1177 ( .C (clk), .D (new_AGEMA_signal_1952), .Q (new_AGEMA_signal_1953) ) ;
    buf_clk new_AGEMA_reg_buffer_1179 ( .C (clk), .D (new_AGEMA_signal_1954), .Q (new_AGEMA_signal_1955) ) ;
    buf_clk new_AGEMA_reg_buffer_1181 ( .C (clk), .D (new_AGEMA_signal_1956), .Q (new_AGEMA_signal_1957) ) ;
    buf_clk new_AGEMA_reg_buffer_1183 ( .C (clk), .D (new_AGEMA_signal_1958), .Q (new_AGEMA_signal_1959) ) ;
    buf_clk new_AGEMA_reg_buffer_1185 ( .C (clk), .D (new_AGEMA_signal_1960), .Q (new_AGEMA_signal_1961) ) ;
    buf_clk new_AGEMA_reg_buffer_1187 ( .C (clk), .D (new_AGEMA_signal_1962), .Q (new_AGEMA_signal_1963) ) ;
    buf_clk new_AGEMA_reg_buffer_1189 ( .C (clk), .D (new_AGEMA_signal_1964), .Q (new_AGEMA_signal_1965) ) ;
    buf_clk new_AGEMA_reg_buffer_1191 ( .C (clk), .D (new_AGEMA_signal_1966), .Q (new_AGEMA_signal_1967) ) ;
    buf_clk new_AGEMA_reg_buffer_1193 ( .C (clk), .D (new_AGEMA_signal_1968), .Q (new_AGEMA_signal_1969) ) ;
    buf_clk new_AGEMA_reg_buffer_1195 ( .C (clk), .D (new_AGEMA_signal_1970), .Q (new_AGEMA_signal_1971) ) ;
    buf_clk new_AGEMA_reg_buffer_1197 ( .C (clk), .D (new_AGEMA_signal_1972), .Q (new_AGEMA_signal_1973) ) ;
    buf_clk new_AGEMA_reg_buffer_1199 ( .C (clk), .D (new_AGEMA_signal_1974), .Q (new_AGEMA_signal_1975) ) ;
    buf_clk new_AGEMA_reg_buffer_1201 ( .C (clk), .D (new_AGEMA_signal_1976), .Q (new_AGEMA_signal_1977) ) ;
    buf_clk new_AGEMA_reg_buffer_1203 ( .C (clk), .D (new_AGEMA_signal_1978), .Q (new_AGEMA_signal_1979) ) ;
    buf_clk new_AGEMA_reg_buffer_1205 ( .C (clk), .D (new_AGEMA_signal_1980), .Q (new_AGEMA_signal_1981) ) ;
    buf_clk new_AGEMA_reg_buffer_1207 ( .C (clk), .D (new_AGEMA_signal_1982), .Q (new_AGEMA_signal_1983) ) ;
    buf_clk new_AGEMA_reg_buffer_1209 ( .C (clk), .D (new_AGEMA_signal_1984), .Q (new_AGEMA_signal_1985) ) ;
    buf_clk new_AGEMA_reg_buffer_1211 ( .C (clk), .D (new_AGEMA_signal_1986), .Q (new_AGEMA_signal_1987) ) ;
    buf_clk new_AGEMA_reg_buffer_1213 ( .C (clk), .D (new_AGEMA_signal_1988), .Q (new_AGEMA_signal_1989) ) ;
    buf_clk new_AGEMA_reg_buffer_1215 ( .C (clk), .D (new_AGEMA_signal_1990), .Q (new_AGEMA_signal_1991) ) ;
    buf_clk new_AGEMA_reg_buffer_1217 ( .C (clk), .D (new_AGEMA_signal_1992), .Q (new_AGEMA_signal_1993) ) ;
    buf_clk new_AGEMA_reg_buffer_1219 ( .C (clk), .D (new_AGEMA_signal_1994), .Q (new_AGEMA_signal_1995) ) ;
    buf_clk new_AGEMA_reg_buffer_1221 ( .C (clk), .D (new_AGEMA_signal_1996), .Q (new_AGEMA_signal_1997) ) ;
    buf_clk new_AGEMA_reg_buffer_1223 ( .C (clk), .D (new_AGEMA_signal_1998), .Q (new_AGEMA_signal_1999) ) ;
    buf_clk new_AGEMA_reg_buffer_1225 ( .C (clk), .D (new_AGEMA_signal_2000), .Q (new_AGEMA_signal_2001) ) ;
    buf_clk new_AGEMA_reg_buffer_1227 ( .C (clk), .D (new_AGEMA_signal_2002), .Q (new_AGEMA_signal_2003) ) ;
    buf_clk new_AGEMA_reg_buffer_1229 ( .C (clk), .D (new_AGEMA_signal_2004), .Q (new_AGEMA_signal_2005) ) ;
    buf_clk new_AGEMA_reg_buffer_1231 ( .C (clk), .D (new_AGEMA_signal_2006), .Q (new_AGEMA_signal_2007) ) ;
    buf_clk new_AGEMA_reg_buffer_1233 ( .C (clk), .D (new_AGEMA_signal_2008), .Q (new_AGEMA_signal_2009) ) ;
    buf_clk new_AGEMA_reg_buffer_1235 ( .C (clk), .D (new_AGEMA_signal_2010), .Q (new_AGEMA_signal_2011) ) ;
    buf_clk new_AGEMA_reg_buffer_1237 ( .C (clk), .D (new_AGEMA_signal_2012), .Q (new_AGEMA_signal_2013) ) ;
    buf_clk new_AGEMA_reg_buffer_1239 ( .C (clk), .D (new_AGEMA_signal_2014), .Q (new_AGEMA_signal_2015) ) ;
    buf_clk new_AGEMA_reg_buffer_1241 ( .C (clk), .D (new_AGEMA_signal_2016), .Q (new_AGEMA_signal_2017) ) ;
    buf_clk new_AGEMA_reg_buffer_1243 ( .C (clk), .D (new_AGEMA_signal_2018), .Q (new_AGEMA_signal_2019) ) ;
    buf_clk new_AGEMA_reg_buffer_1245 ( .C (clk), .D (new_AGEMA_signal_2020), .Q (new_AGEMA_signal_2021) ) ;
    buf_clk new_AGEMA_reg_buffer_1247 ( .C (clk), .D (new_AGEMA_signal_2022), .Q (new_AGEMA_signal_2023) ) ;
    buf_clk new_AGEMA_reg_buffer_1249 ( .C (clk), .D (new_AGEMA_signal_2024), .Q (new_AGEMA_signal_2025) ) ;
    buf_clk new_AGEMA_reg_buffer_1251 ( .C (clk), .D (new_AGEMA_signal_2026), .Q (new_AGEMA_signal_2027) ) ;
    buf_clk new_AGEMA_reg_buffer_1253 ( .C (clk), .D (new_AGEMA_signal_2028), .Q (new_AGEMA_signal_2029) ) ;
    buf_clk new_AGEMA_reg_buffer_1255 ( .C (clk), .D (new_AGEMA_signal_2030), .Q (new_AGEMA_signal_2031) ) ;
    buf_clk new_AGEMA_reg_buffer_1257 ( .C (clk), .D (new_AGEMA_signal_2032), .Q (new_AGEMA_signal_2033) ) ;
    buf_clk new_AGEMA_reg_buffer_1259 ( .C (clk), .D (new_AGEMA_signal_2034), .Q (new_AGEMA_signal_2035) ) ;
    buf_clk new_AGEMA_reg_buffer_1261 ( .C (clk), .D (new_AGEMA_signal_2036), .Q (new_AGEMA_signal_2037) ) ;
    buf_clk new_AGEMA_reg_buffer_1263 ( .C (clk), .D (new_AGEMA_signal_2038), .Q (new_AGEMA_signal_2039) ) ;
    buf_clk new_AGEMA_reg_buffer_1265 ( .C (clk), .D (new_AGEMA_signal_2040), .Q (new_AGEMA_signal_2041) ) ;
    buf_clk new_AGEMA_reg_buffer_1267 ( .C (clk), .D (new_AGEMA_signal_2042), .Q (new_AGEMA_signal_2043) ) ;
    buf_clk new_AGEMA_reg_buffer_1269 ( .C (clk), .D (new_AGEMA_signal_2044), .Q (new_AGEMA_signal_2045) ) ;
    buf_clk new_AGEMA_reg_buffer_1271 ( .C (clk), .D (new_AGEMA_signal_2046), .Q (new_AGEMA_signal_2047) ) ;
    buf_clk new_AGEMA_reg_buffer_1273 ( .C (clk), .D (new_AGEMA_signal_2048), .Q (new_AGEMA_signal_2049) ) ;
    buf_clk new_AGEMA_reg_buffer_1275 ( .C (clk), .D (new_AGEMA_signal_2050), .Q (new_AGEMA_signal_2051) ) ;
    buf_clk new_AGEMA_reg_buffer_1277 ( .C (clk), .D (new_AGEMA_signal_2052), .Q (new_AGEMA_signal_2053) ) ;
    buf_clk new_AGEMA_reg_buffer_1279 ( .C (clk), .D (new_AGEMA_signal_2054), .Q (new_AGEMA_signal_2055) ) ;
    buf_clk new_AGEMA_reg_buffer_1281 ( .C (clk), .D (new_AGEMA_signal_2056), .Q (new_AGEMA_signal_2057) ) ;
    buf_clk new_AGEMA_reg_buffer_1283 ( .C (clk), .D (new_AGEMA_signal_2058), .Q (new_AGEMA_signal_2059) ) ;
    buf_clk new_AGEMA_reg_buffer_1285 ( .C (clk), .D (new_AGEMA_signal_2060), .Q (new_AGEMA_signal_2061) ) ;
    buf_clk new_AGEMA_reg_buffer_1287 ( .C (clk), .D (new_AGEMA_signal_2062), .Q (new_AGEMA_signal_2063) ) ;
    buf_clk new_AGEMA_reg_buffer_1289 ( .C (clk), .D (new_AGEMA_signal_2064), .Q (new_AGEMA_signal_2065) ) ;
    buf_clk new_AGEMA_reg_buffer_1291 ( .C (clk), .D (new_AGEMA_signal_2066), .Q (new_AGEMA_signal_2067) ) ;
    buf_clk new_AGEMA_reg_buffer_1293 ( .C (clk), .D (new_AGEMA_signal_2068), .Q (new_AGEMA_signal_2069) ) ;
    buf_clk new_AGEMA_reg_buffer_1295 ( .C (clk), .D (new_AGEMA_signal_2070), .Q (new_AGEMA_signal_2071) ) ;
    buf_clk new_AGEMA_reg_buffer_1297 ( .C (clk), .D (new_AGEMA_signal_2072), .Q (new_AGEMA_signal_2073) ) ;
    buf_clk new_AGEMA_reg_buffer_1299 ( .C (clk), .D (new_AGEMA_signal_2074), .Q (new_AGEMA_signal_2075) ) ;
    buf_clk new_AGEMA_reg_buffer_1301 ( .C (clk), .D (new_AGEMA_signal_2076), .Q (new_AGEMA_signal_2077) ) ;
    buf_clk new_AGEMA_reg_buffer_1303 ( .C (clk), .D (new_AGEMA_signal_2078), .Q (new_AGEMA_signal_2079) ) ;
    buf_clk new_AGEMA_reg_buffer_1305 ( .C (clk), .D (new_AGEMA_signal_2080), .Q (new_AGEMA_signal_2081) ) ;
    buf_clk new_AGEMA_reg_buffer_1307 ( .C (clk), .D (new_AGEMA_signal_2082), .Q (new_AGEMA_signal_2083) ) ;
    buf_clk new_AGEMA_reg_buffer_1309 ( .C (clk), .D (new_AGEMA_signal_2084), .Q (new_AGEMA_signal_2085) ) ;
    buf_clk new_AGEMA_reg_buffer_1311 ( .C (clk), .D (new_AGEMA_signal_2086), .Q (new_AGEMA_signal_2087) ) ;
    buf_clk new_AGEMA_reg_buffer_1313 ( .C (clk), .D (new_AGEMA_signal_2088), .Q (new_AGEMA_signal_2089) ) ;
    buf_clk new_AGEMA_reg_buffer_1315 ( .C (clk), .D (new_AGEMA_signal_2090), .Q (new_AGEMA_signal_2091) ) ;
    buf_clk new_AGEMA_reg_buffer_1317 ( .C (clk), .D (new_AGEMA_signal_2092), .Q (new_AGEMA_signal_2093) ) ;
    buf_clk new_AGEMA_reg_buffer_1319 ( .C (clk), .D (new_AGEMA_signal_2094), .Q (new_AGEMA_signal_2095) ) ;
    buf_clk new_AGEMA_reg_buffer_1321 ( .C (clk), .D (new_AGEMA_signal_2096), .Q (new_AGEMA_signal_2097) ) ;
    buf_clk new_AGEMA_reg_buffer_1323 ( .C (clk), .D (new_AGEMA_signal_2098), .Q (new_AGEMA_signal_2099) ) ;
    buf_clk new_AGEMA_reg_buffer_1325 ( .C (clk), .D (new_AGEMA_signal_2100), .Q (new_AGEMA_signal_2101) ) ;
    buf_clk new_AGEMA_reg_buffer_1327 ( .C (clk), .D (new_AGEMA_signal_2102), .Q (new_AGEMA_signal_2103) ) ;
    buf_clk new_AGEMA_reg_buffer_1329 ( .C (clk), .D (new_AGEMA_signal_2104), .Q (new_AGEMA_signal_2105) ) ;
    buf_clk new_AGEMA_reg_buffer_1331 ( .C (clk), .D (new_AGEMA_signal_2106), .Q (new_AGEMA_signal_2107) ) ;
    buf_clk new_AGEMA_reg_buffer_1333 ( .C (clk), .D (new_AGEMA_signal_2108), .Q (new_AGEMA_signal_2109) ) ;
    buf_clk new_AGEMA_reg_buffer_1335 ( .C (clk), .D (new_AGEMA_signal_2110), .Q (new_AGEMA_signal_2111) ) ;
    buf_clk new_AGEMA_reg_buffer_1337 ( .C (clk), .D (new_AGEMA_signal_2112), .Q (new_AGEMA_signal_2113) ) ;
    buf_clk new_AGEMA_reg_buffer_1339 ( .C (clk), .D (new_AGEMA_signal_2114), .Q (new_AGEMA_signal_2115) ) ;
    buf_clk new_AGEMA_reg_buffer_1341 ( .C (clk), .D (new_AGEMA_signal_2116), .Q (new_AGEMA_signal_2117) ) ;
    buf_clk new_AGEMA_reg_buffer_1343 ( .C (clk), .D (new_AGEMA_signal_2118), .Q (new_AGEMA_signal_2119) ) ;
    buf_clk new_AGEMA_reg_buffer_1345 ( .C (clk), .D (new_AGEMA_signal_2120), .Q (new_AGEMA_signal_2121) ) ;
    buf_clk new_AGEMA_reg_buffer_1347 ( .C (clk), .D (new_AGEMA_signal_2122), .Q (new_AGEMA_signal_2123) ) ;
    buf_clk new_AGEMA_reg_buffer_1349 ( .C (clk), .D (new_AGEMA_signal_2124), .Q (new_AGEMA_signal_2125) ) ;
    buf_clk new_AGEMA_reg_buffer_1351 ( .C (clk), .D (new_AGEMA_signal_2126), .Q (new_AGEMA_signal_2127) ) ;
    buf_clk new_AGEMA_reg_buffer_1353 ( .C (clk), .D (new_AGEMA_signal_2128), .Q (new_AGEMA_signal_2129) ) ;
    buf_clk new_AGEMA_reg_buffer_1355 ( .C (clk), .D (new_AGEMA_signal_2130), .Q (new_AGEMA_signal_2131) ) ;
    buf_clk new_AGEMA_reg_buffer_1357 ( .C (clk), .D (new_AGEMA_signal_2132), .Q (new_AGEMA_signal_2133) ) ;
    buf_clk new_AGEMA_reg_buffer_1358 ( .C (clk), .D (keyFF_keystate_gff_20_s_next_state[0]), .Q (new_AGEMA_signal_2134) ) ;
    buf_clk new_AGEMA_reg_buffer_1359 ( .C (clk), .D (new_AGEMA_signal_1448), .Q (new_AGEMA_signal_2135) ) ;

    /* register cells */
    DFF_X1 fsm_cnt_rnd_count_reg_reg_4__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1567), .Q (counter[4]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1569), .Q (counter[2]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1571), .Q (counter[0]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1573), .Q (counter[3]), .QN () ) ;
    DFF_X1 fsm_cnt_rnd_count_reg_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1575), .Q (fsm_cnt_rnd_n24), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_2__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1577), .Q (fsm_countSerial[2]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1579), .Q (fsm_countSerial[0]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_3__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1581), .Q (fsm_countSerial[3]), .QN () ) ;
    DFF_X1 fsm_cnt_ser_count_reg_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1583), .Q (fsm_countSerial[1]), .QN () ) ;
    DFF_X1 fsm_ps_state_reg_0__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1585), .Q (fsm_ps_state_0_), .QN () ) ;
    DFF_X1 fsm_ps_state_reg_1__FF_FF ( .CK (clk), .D (new_AGEMA_signal_1587), .Q (fsm_ps_state_1_), .QN () ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_1_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1589, new_AGEMA_signal_1588}), .Q ({data_out_s1[0], data_out_s0[0]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_1_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1464, stateFF_state_gff_1_s_next_state[2]}), .Q ({data_out_s1[2], data_out_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_1_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1463, stateFF_state_gff_1_s_next_state[1]}), .Q ({data_out_s1[1], data_out_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_1_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1470, stateFF_state_gff_1_s_next_state[3]}), .Q ({data_out_s1[3], data_out_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_2_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1593, new_AGEMA_signal_1591}), .Q ({data_out_s1[7], data_out_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_2_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1597, new_AGEMA_signal_1595}), .Q ({data_out_s1[6], data_out_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_2_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1601, new_AGEMA_signal_1599}), .Q ({data_out_s1[5], data_out_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_2_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1605, new_AGEMA_signal_1603}), .Q ({data_out_s1[4], data_out_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_3_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1609, new_AGEMA_signal_1607}), .Q ({data_out_s1[11], data_out_s0[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_3_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1613, new_AGEMA_signal_1611}), .Q ({data_out_s1[10], data_out_s0[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_3_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1617, new_AGEMA_signal_1615}), .Q ({data_out_s1[9], data_out_s0[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_3_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1621, new_AGEMA_signal_1619}), .Q ({data_out_s1[8], data_out_s0[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_4_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1625, new_AGEMA_signal_1623}), .Q ({data_out_s1[15], data_out_s0[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_4_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1629, new_AGEMA_signal_1627}), .Q ({data_out_s1[14], data_out_s0[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_4_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1633, new_AGEMA_signal_1631}), .Q ({data_out_s1[13], data_out_s0[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_4_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1637, new_AGEMA_signal_1635}), .Q ({data_out_s1[12], data_out_s0[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_5_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1641, new_AGEMA_signal_1639}), .Q ({data_out_s1[19], data_out_s0[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_5_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1645, new_AGEMA_signal_1643}), .Q ({data_out_s1[18], data_out_s0[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_5_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1649, new_AGEMA_signal_1647}), .Q ({data_out_s1[17], data_out_s0[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_5_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1653, new_AGEMA_signal_1651}), .Q ({data_out_s1[16], data_out_s0[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_6_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1657, new_AGEMA_signal_1655}), .Q ({data_out_s1[23], data_out_s0[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_6_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1661, new_AGEMA_signal_1659}), .Q ({data_out_s1[22], data_out_s0[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_6_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1665, new_AGEMA_signal_1663}), .Q ({data_out_s1[21], data_out_s0[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_6_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1669, new_AGEMA_signal_1667}), .Q ({data_out_s1[20], data_out_s0[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_7_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1673, new_AGEMA_signal_1671}), .Q ({data_out_s1[27], data_out_s0[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_7_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1677, new_AGEMA_signal_1675}), .Q ({data_out_s1[26], data_out_s0[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_7_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1681, new_AGEMA_signal_1679}), .Q ({data_out_s1[25], data_out_s0[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_7_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1685, new_AGEMA_signal_1683}), .Q ({data_out_s1[24], data_out_s0[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_8_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1689, new_AGEMA_signal_1687}), .Q ({data_out_s1[31], data_out_s0[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_8_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1693, new_AGEMA_signal_1691}), .Q ({data_out_s1[30], data_out_s0[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_8_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1697, new_AGEMA_signal_1695}), .Q ({data_out_s1[29], data_out_s0[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_8_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1701, new_AGEMA_signal_1699}), .Q ({data_out_s1[28], data_out_s0[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_9_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1705, new_AGEMA_signal_1703}), .Q ({data_out_s1[35], data_out_s0[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_9_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1709, new_AGEMA_signal_1707}), .Q ({data_out_s1[34], data_out_s0[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_9_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1713, new_AGEMA_signal_1711}), .Q ({data_out_s1[33], data_out_s0[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_9_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1717, new_AGEMA_signal_1715}), .Q ({data_out_s1[32], data_out_s0[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_10_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1721, new_AGEMA_signal_1719}), .Q ({data_out_s1[39], data_out_s0[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_10_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1725, new_AGEMA_signal_1723}), .Q ({data_out_s1[38], data_out_s0[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_10_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1729, new_AGEMA_signal_1727}), .Q ({data_out_s1[37], data_out_s0[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_10_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1733, new_AGEMA_signal_1731}), .Q ({data_out_s1[36], data_out_s0[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_11_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1737, new_AGEMA_signal_1735}), .Q ({data_out_s1[43], data_out_s0[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_11_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1741, new_AGEMA_signal_1739}), .Q ({data_out_s1[42], data_out_s0[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_11_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1745, new_AGEMA_signal_1743}), .Q ({data_out_s1[41], data_out_s0[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_11_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1749, new_AGEMA_signal_1747}), .Q ({data_out_s1[40], data_out_s0[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_12_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1753, new_AGEMA_signal_1751}), .Q ({data_out_s1[47], data_out_s0[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_12_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1757, new_AGEMA_signal_1755}), .Q ({data_out_s1[46], data_out_s0[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_12_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1761, new_AGEMA_signal_1759}), .Q ({data_out_s1[45], data_out_s0[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_12_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1765, new_AGEMA_signal_1763}), .Q ({data_out_s1[44], data_out_s0[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_13_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1769, new_AGEMA_signal_1767}), .Q ({data_out_s1[51], data_out_s0[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_13_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1773, new_AGEMA_signal_1771}), .Q ({data_out_s1[50], data_out_s0[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_13_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1777, new_AGEMA_signal_1775}), .Q ({data_out_s1[49], data_out_s0[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_13_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1781, new_AGEMA_signal_1779}), .Q ({data_out_s1[48], data_out_s0[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_14_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1785, new_AGEMA_signal_1783}), .Q ({data_out_s1[55], data_out_s0[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_14_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1789, new_AGEMA_signal_1787}), .Q ({data_out_s1[54], data_out_s0[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_14_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1793, new_AGEMA_signal_1791}), .Q ({data_out_s1[53], data_out_s0[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_14_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1797, new_AGEMA_signal_1795}), .Q ({data_out_s1[52], data_out_s0[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_15_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1801, new_AGEMA_signal_1799}), .Q ({data_out_s1[59], data_out_s0[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_15_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1805, new_AGEMA_signal_1803}), .Q ({data_out_s1[58], data_out_s0[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_15_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1809, new_AGEMA_signal_1807}), .Q ({data_out_s1[57], data_out_s0[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_15_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1813, new_AGEMA_signal_1811}), .Q ({data_out_s1[56], data_out_s0[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_16_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1817, new_AGEMA_signal_1815}), .Q ({data_out_s1[63], data_out_s0[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_16_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1821, new_AGEMA_signal_1819}), .Q ({data_out_s1[62], data_out_s0[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_16_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1825, new_AGEMA_signal_1823}), .Q ({data_out_s1[61], data_out_s0[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) stateFF_state_gff_16_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1829, new_AGEMA_signal_1827}), .Q ({data_out_s1[60], data_out_s0[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_1_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1833, new_AGEMA_signal_1831}), .Q ({new_AGEMA_signal_1064, keyFF_outputPar[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_1_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1837, new_AGEMA_signal_1835}), .Q ({new_AGEMA_signal_1291, keyRegKS[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_1_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1841, new_AGEMA_signal_1839}), .Q ({new_AGEMA_signal_1289, keyRegKS[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_1_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1845, new_AGEMA_signal_1843}), .Q ({new_AGEMA_signal_1287, keyRegKS[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_2_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1849, new_AGEMA_signal_1847}), .Q ({new_AGEMA_signal_1076, keyFF_outputPar[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_2_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1853, new_AGEMA_signal_1851}), .Q ({new_AGEMA_signal_1073, keyFF_outputPar[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_2_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1857, new_AGEMA_signal_1855}), .Q ({new_AGEMA_signal_1070, keyFF_outputPar[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_2_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1861, new_AGEMA_signal_1859}), .Q ({new_AGEMA_signal_1067, keyFF_outputPar[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_3_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1865, new_AGEMA_signal_1863}), .Q ({new_AGEMA_signal_1088, keyFF_outputPar[11]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_3_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1869, new_AGEMA_signal_1867}), .Q ({new_AGEMA_signal_1085, keyFF_outputPar[10]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_3_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1873, new_AGEMA_signal_1871}), .Q ({new_AGEMA_signal_1082, keyFF_outputPar[9]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_3_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1877, new_AGEMA_signal_1875}), .Q ({new_AGEMA_signal_1079, keyFF_outputPar[8]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_4_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1881, new_AGEMA_signal_1879}), .Q ({new_AGEMA_signal_1100, keyFF_outputPar[15]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_4_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1885, new_AGEMA_signal_1883}), .Q ({new_AGEMA_signal_1097, keyFF_outputPar[14]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_4_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1889, new_AGEMA_signal_1887}), .Q ({new_AGEMA_signal_1094, keyFF_outputPar[13]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_4_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1893, new_AGEMA_signal_1891}), .Q ({new_AGEMA_signal_1091, keyFF_outputPar[12]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_5_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1897, new_AGEMA_signal_1895}), .Q ({new_AGEMA_signal_1274, keyFF_outputPar[19]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_5_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1901, new_AGEMA_signal_1899}), .Q ({new_AGEMA_signal_1062, keyFF_outputPar[18]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_5_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1905, new_AGEMA_signal_1903}), .Q ({new_AGEMA_signal_1106, keyFF_outputPar[17]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_5_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1909, new_AGEMA_signal_1907}), .Q ({new_AGEMA_signal_1103, keyFF_outputPar[16]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_6_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1913, new_AGEMA_signal_1911}), .Q ({new_AGEMA_signal_1109, keyFF_outputPar[23]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_6_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1917, new_AGEMA_signal_1915}), .Q ({new_AGEMA_signal_1056, keyFF_outputPar[22]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_6_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1921, new_AGEMA_signal_1919}), .Q ({new_AGEMA_signal_1058, keyFF_outputPar[21]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_6_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1925, new_AGEMA_signal_1923}), .Q ({new_AGEMA_signal_1060, keyFF_outputPar[20]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_7_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1929, new_AGEMA_signal_1927}), .Q ({new_AGEMA_signal_1121, keyFF_outputPar[27]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_7_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1933, new_AGEMA_signal_1931}), .Q ({new_AGEMA_signal_1118, keyFF_outputPar[26]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_7_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1937, new_AGEMA_signal_1935}), .Q ({new_AGEMA_signal_1115, keyFF_outputPar[25]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_7_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1941, new_AGEMA_signal_1939}), .Q ({new_AGEMA_signal_1112, keyFF_outputPar[24]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_8_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1945, new_AGEMA_signal_1943}), .Q ({new_AGEMA_signal_1133, keyFF_outputPar[31]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_8_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1949, new_AGEMA_signal_1947}), .Q ({new_AGEMA_signal_1130, keyFF_outputPar[30]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_8_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1953, new_AGEMA_signal_1951}), .Q ({new_AGEMA_signal_1127, keyFF_outputPar[29]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_8_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1957, new_AGEMA_signal_1955}), .Q ({new_AGEMA_signal_1124, keyFF_outputPar[28]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_9_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1961, new_AGEMA_signal_1959}), .Q ({new_AGEMA_signal_1145, keyFF_outputPar[35]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_9_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1965, new_AGEMA_signal_1963}), .Q ({new_AGEMA_signal_1142, keyFF_outputPar[34]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_9_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1969, new_AGEMA_signal_1967}), .Q ({new_AGEMA_signal_1139, keyFF_outputPar[33]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_9_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1973, new_AGEMA_signal_1971}), .Q ({new_AGEMA_signal_1136, keyFF_outputPar[32]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_10_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1977, new_AGEMA_signal_1975}), .Q ({new_AGEMA_signal_1157, keyFF_outputPar[39]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_10_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1981, new_AGEMA_signal_1979}), .Q ({new_AGEMA_signal_1154, keyFF_outputPar[38]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_10_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1985, new_AGEMA_signal_1983}), .Q ({new_AGEMA_signal_1151, keyFF_outputPar[37]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_10_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1989, new_AGEMA_signal_1987}), .Q ({new_AGEMA_signal_1148, keyFF_outputPar[36]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_11_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1993, new_AGEMA_signal_1991}), .Q ({new_AGEMA_signal_1169, keyFF_outputPar[43]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_11_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1997, new_AGEMA_signal_1995}), .Q ({new_AGEMA_signal_1166, keyFF_outputPar[42]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_11_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2001, new_AGEMA_signal_1999}), .Q ({new_AGEMA_signal_1163, keyFF_outputPar[41]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_11_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2005, new_AGEMA_signal_2003}), .Q ({new_AGEMA_signal_1160, keyFF_outputPar[40]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_12_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2009, new_AGEMA_signal_2007}), .Q ({new_AGEMA_signal_1181, keyFF_outputPar[47]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_12_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2013, new_AGEMA_signal_2011}), .Q ({new_AGEMA_signal_1178, keyFF_outputPar[46]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_12_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2017, new_AGEMA_signal_2015}), .Q ({new_AGEMA_signal_1175, keyFF_outputPar[45]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_12_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2021, new_AGEMA_signal_2019}), .Q ({new_AGEMA_signal_1172, keyFF_outputPar[44]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_13_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2025, new_AGEMA_signal_2023}), .Q ({new_AGEMA_signal_1193, keyFF_outputPar[51]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_13_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2029, new_AGEMA_signal_2027}), .Q ({new_AGEMA_signal_1190, keyFF_outputPar[50]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_13_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2033, new_AGEMA_signal_2031}), .Q ({new_AGEMA_signal_1187, keyFF_outputPar[49]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_13_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2037, new_AGEMA_signal_2035}), .Q ({new_AGEMA_signal_1184, keyFF_outputPar[48]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_14_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2041, new_AGEMA_signal_2039}), .Q ({new_AGEMA_signal_1205, keyFF_outputPar[55]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_14_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2045, new_AGEMA_signal_2043}), .Q ({new_AGEMA_signal_1202, keyFF_outputPar[54]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_14_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2049, new_AGEMA_signal_2047}), .Q ({new_AGEMA_signal_1199, keyFF_outputPar[53]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_14_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2053, new_AGEMA_signal_2051}), .Q ({new_AGEMA_signal_1196, keyFF_outputPar[52]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_15_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2057, new_AGEMA_signal_2055}), .Q ({new_AGEMA_signal_1217, keyFF_outputPar[59]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_15_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2061, new_AGEMA_signal_2059}), .Q ({new_AGEMA_signal_1214, keyFF_outputPar[58]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_15_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2065, new_AGEMA_signal_2063}), .Q ({new_AGEMA_signal_1211, keyFF_outputPar[57]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_15_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2069, new_AGEMA_signal_2067}), .Q ({new_AGEMA_signal_1208, keyFF_outputPar[56]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_16_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2073, new_AGEMA_signal_2071}), .Q ({new_AGEMA_signal_1229, keyFF_outputPar[63]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_16_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2077, new_AGEMA_signal_2075}), .Q ({new_AGEMA_signal_1226, keyFF_outputPar[62]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_16_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2081, new_AGEMA_signal_2079}), .Q ({new_AGEMA_signal_1223, keyFF_outputPar[61]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_16_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2085, new_AGEMA_signal_2083}), .Q ({new_AGEMA_signal_1220, keyFF_outputPar[60]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_17_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2089, new_AGEMA_signal_2087}), .Q ({new_AGEMA_signal_1241, keyFF_outputPar[67]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_17_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2093, new_AGEMA_signal_2091}), .Q ({new_AGEMA_signal_1238, keyFF_outputPar[66]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_17_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2097, new_AGEMA_signal_2095}), .Q ({new_AGEMA_signal_1235, keyFF_outputPar[65]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_17_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2101, new_AGEMA_signal_2099}), .Q ({new_AGEMA_signal_1232, keyFF_outputPar[64]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_18_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2105, new_AGEMA_signal_2103}), .Q ({new_AGEMA_signal_1253, keyFF_outputPar[71]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_18_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2109, new_AGEMA_signal_2107}), .Q ({new_AGEMA_signal_1250, keyFF_outputPar[70]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_18_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2113, new_AGEMA_signal_2111}), .Q ({new_AGEMA_signal_1247, keyFF_outputPar[69]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_18_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2117, new_AGEMA_signal_2115}), .Q ({new_AGEMA_signal_1244, keyFF_outputPar[68]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_19_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2121, new_AGEMA_signal_2119}), .Q ({new_AGEMA_signal_1265, keyFF_outputPar[75]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_19_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2125, new_AGEMA_signal_2123}), .Q ({new_AGEMA_signal_1262, keyFF_outputPar[74]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_19_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2129, new_AGEMA_signal_2127}), .Q ({new_AGEMA_signal_1259, keyFF_outputPar[73]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_19_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2133, new_AGEMA_signal_2131}), .Q ({new_AGEMA_signal_1256, keyFF_outputPar[72]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_20_s_current_state_reg_3__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1471, keyFF_keystate_gff_20_s_next_state[3]}), .Q ({new_AGEMA_signal_865, roundkey[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_20_s_current_state_reg_2__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1466, keyFF_keystate_gff_20_s_next_state[2]}), .Q ({new_AGEMA_signal_862, roundkey[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_20_s_current_state_reg_1__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_1465, keyFF_keystate_gff_20_s_next_state[1]}), .Q ({new_AGEMA_signal_859, roundkey[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) keyFF_keystate_gff_20_s_current_state_reg_0__FF_FF ( .clk (clk), .D ({new_AGEMA_signal_2135, new_AGEMA_signal_2134}), .Q ({new_AGEMA_signal_856, roundkey[0]}) ) ;
endmodule
