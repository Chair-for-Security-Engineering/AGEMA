/* modified netlist. Source: module sbox in file Designs/SkinnySbox/AGEMA/sbox_opt_correct/sbox.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d1 (X_s0, clk, X_s1, Fresh, Y_s0, Y_s1);
    input [3:0] X_s0 ;
    input clk ;
    input [3:0] X_s1 ;
    input [3:0] Fresh ;
    output [3:0] Y_s0 ;
    output [3:0] Y_s1 ;
    wire signal_33 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_47 ;
    wire signal_48 ;
    wire signal_49 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_56 ;
    wire signal_58 ;
    wire signal_60 ;
    wire signal_62 ;
    wire signal_64 ;
    wire signal_65 ;
    wire signal_66 ;
    wire signal_67 ;
    wire signal_68 ;
    wire signal_69 ;
    wire signal_70 ;
    wire signal_71 ;
    wire signal_72 ;
    wire signal_73 ;
    wire signal_74 ;
    wire signal_75 ;
    wire signal_76 ;
    wire signal_77 ;
    wire signal_78 ;
    wire signal_79 ;
    wire signal_80 ;
    wire signal_81 ;
    wire signal_82 ;
    wire signal_83 ;
    wire signal_84 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_95 ;
    wire signal_96 ;
    wire signal_97 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_104 ;
    wire signal_105 ;
    wire signal_106 ;
    wire signal_107 ;
    wire signal_108 ;
    wire signal_109 ;
    wire signal_110 ;
    wire signal_111 ;
    wire signal_112 ;
    wire signal_113 ;
    wire signal_114 ;
    wire signal_115 ;
    wire signal_116 ;
    wire signal_117 ;
    wire signal_118 ;
    wire signal_119 ;
    wire signal_120 ;
    wire signal_121 ;
    wire signal_122 ;
    wire signal_123 ;
    wire signal_124 ;
    wire signal_125 ;
    wire signal_126 ;
    wire signal_127 ;
    wire signal_128 ;
    wire signal_129 ;
    wire signal_130 ;
    wire signal_131 ;
    wire signal_132 ;
    wire signal_133 ;
    wire signal_134 ;
    wire signal_135 ;
    wire signal_136 ;
    wire signal_137 ;
    wire signal_138 ;
    wire signal_139 ;
    wire signal_140 ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(1)) cell_26 ( .a ({X_s1[2], X_s0[2]}), .b ({signal_58, signal_37}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_27 ( .a ({X_s1[3], X_s0[3]}), .b ({X_s1[2], X_s0[2]}), .c ({signal_60, signal_38}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_28 ( .a ({X_s1[2], X_s0[2]}), .b ({X_s1[0], X_s0[0]}), .c ({signal_62, signal_39}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_29 ( .a ({X_s1[2], X_s0[2]}), .b ({X_s1[1], X_s0[1]}), .c ({signal_64, signal_40}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_31 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_62, signal_39}), .c ({signal_66, signal_42}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_32 ( .a ({X_s1[1], X_s0[1]}), .b ({signal_60, signal_38}), .c ({signal_67, signal_43}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_33 ( .a ({X_s1[2], X_s0[2]}), .b ({signal_62, signal_39}), .c ({signal_68, signal_44}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_34 ( .a ({signal_68, signal_44}), .b ({signal_69, signal_45}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_36 ( .a ({signal_67, signal_43}), .b ({signal_68, signal_44}), .c ({signal_71, signal_47}) ) ;

    /* cells in depth 1 */
    buf_clk cell_50 ( .C (clk), .D (signal_38), .Q (signal_93) ) ;
    buf_clk cell_52 ( .C (clk), .D (signal_60), .Q (signal_95) ) ;
    buf_clk cell_54 ( .C (clk), .D (signal_42), .Q (signal_97) ) ;
    buf_clk cell_56 ( .C (clk), .D (signal_66), .Q (signal_99) ) ;
    buf_clk cell_58 ( .C (clk), .D (signal_47), .Q (signal_101) ) ;
    buf_clk cell_60 ( .C (clk), .D (signal_71), .Q (signal_103) ) ;
    buf_clk cell_62 ( .C (clk), .D (signal_39), .Q (signal_105) ) ;
    buf_clk cell_64 ( .C (clk), .D (signal_62), .Q (signal_107) ) ;
    buf_clk cell_66 ( .C (clk), .D (X_s0[1]), .Q (signal_109) ) ;
    buf_clk cell_68 ( .C (clk), .D (X_s1[1]), .Q (signal_111) ) ;
    buf_clk cell_70 ( .C (clk), .D (signal_45), .Q (signal_113) ) ;
    buf_clk cell_72 ( .C (clk), .D (signal_69), .Q (signal_115) ) ;
    buf_clk cell_78 ( .C (clk), .D (signal_40), .Q (signal_121) ) ;
    buf_clk cell_82 ( .C (clk), .D (signal_64), .Q (signal_125) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_30 ( .a ({signal_58, signal_37}), .b ({signal_64, signal_40}), .clk (clk), .r (Fresh[0]), .c ({signal_65, signal_41}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_35 ( .a ({signal_58, signal_37}), .b ({signal_67, signal_43}), .clk (clk), .r (Fresh[1]), .c ({signal_70, signal_46}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_37 ( .a ({signal_96, signal_94}), .b ({signal_65, signal_41}), .c ({signal_72, signal_48}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_38 ( .a ({signal_72, signal_48}), .b ({signal_73, signal_36}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_39 ( .a ({signal_100, signal_98}), .b ({signal_70, signal_46}), .c ({signal_74, signal_49}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_40 ( .a ({signal_65, signal_41}), .b ({signal_104, signal_102}), .c ({signal_75, signal_50}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_41 ( .a ({signal_108, signal_106}), .b ({signal_70, signal_46}), .c ({signal_76, signal_51}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_44 ( .a ({signal_65, signal_41}), .b ({signal_76, signal_51}), .c ({signal_79, signal_54}) ) ;
    not_masked #(.security_order(1), .pipeline(1)) cell_45 ( .a ({signal_79, signal_54}), .b ({signal_80, signal_35}) ) ;
    buf_clk cell_51 ( .C (clk), .D (signal_93), .Q (signal_94) ) ;
    buf_clk cell_53 ( .C (clk), .D (signal_95), .Q (signal_96) ) ;
    buf_clk cell_55 ( .C (clk), .D (signal_97), .Q (signal_98) ) ;
    buf_clk cell_57 ( .C (clk), .D (signal_99), .Q (signal_100) ) ;
    buf_clk cell_59 ( .C (clk), .D (signal_101), .Q (signal_102) ) ;
    buf_clk cell_61 ( .C (clk), .D (signal_103), .Q (signal_104) ) ;
    buf_clk cell_63 ( .C (clk), .D (signal_105), .Q (signal_106) ) ;
    buf_clk cell_65 ( .C (clk), .D (signal_107), .Q (signal_108) ) ;
    buf_clk cell_67 ( .C (clk), .D (signal_109), .Q (signal_110) ) ;
    buf_clk cell_69 ( .C (clk), .D (signal_111), .Q (signal_112) ) ;
    buf_clk cell_71 ( .C (clk), .D (signal_113), .Q (signal_114) ) ;
    buf_clk cell_73 ( .C (clk), .D (signal_115), .Q (signal_116) ) ;
    buf_clk cell_79 ( .C (clk), .D (signal_121), .Q (signal_122) ) ;
    buf_clk cell_83 ( .C (clk), .D (signal_125), .Q (signal_126) ) ;

    /* cells in depth 3 */
    buf_clk cell_74 ( .C (clk), .D (signal_41), .Q (signal_117) ) ;
    buf_clk cell_76 ( .C (clk), .D (signal_65), .Q (signal_119) ) ;
    buf_clk cell_80 ( .C (clk), .D (signal_122), .Q (signal_123) ) ;
    buf_clk cell_84 ( .C (clk), .D (signal_126), .Q (signal_127) ) ;
    buf_clk cell_86 ( .C (clk), .D (signal_51), .Q (signal_129) ) ;
    buf_clk cell_88 ( .C (clk), .D (signal_76), .Q (signal_131) ) ;
    buf_clk cell_90 ( .C (clk), .D (signal_35), .Q (signal_133) ) ;
    buf_clk cell_92 ( .C (clk), .D (signal_80), .Q (signal_135) ) ;
    buf_clk cell_94 ( .C (clk), .D (signal_36), .Q (signal_137) ) ;
    buf_clk cell_96 ( .C (clk), .D (signal_73), .Q (signal_139) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_42 ( .a ({signal_112, signal_110}), .b ({signal_74, signal_49}), .clk (clk), .r (Fresh[2]), .c ({signal_77, signal_52}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(1)) cell_43 ( .a ({signal_116, signal_114}), .b ({signal_75, signal_50}), .clk (clk), .r (Fresh[3]), .c ({signal_78, signal_53}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_46 ( .a ({signal_120, signal_118}), .b ({signal_77, signal_52}), .c ({signal_81, signal_55}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_47 ( .a ({signal_128, signal_124}), .b ({signal_77, signal_52}), .c ({signal_82, signal_56}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_48 ( .a ({signal_132, signal_130}), .b ({signal_82, signal_56}), .c ({signal_83, signal_33}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(1)) cell_49 ( .a ({signal_78, signal_53}), .b ({signal_81, signal_55}), .c ({signal_84, signal_34}) ) ;
    buf_clk cell_75 ( .C (clk), .D (signal_117), .Q (signal_118) ) ;
    buf_clk cell_77 ( .C (clk), .D (signal_119), .Q (signal_120) ) ;
    buf_clk cell_81 ( .C (clk), .D (signal_123), .Q (signal_124) ) ;
    buf_clk cell_85 ( .C (clk), .D (signal_127), .Q (signal_128) ) ;
    buf_clk cell_87 ( .C (clk), .D (signal_129), .Q (signal_130) ) ;
    buf_clk cell_89 ( .C (clk), .D (signal_131), .Q (signal_132) ) ;
    buf_clk cell_91 ( .C (clk), .D (signal_133), .Q (signal_134) ) ;
    buf_clk cell_93 ( .C (clk), .D (signal_135), .Q (signal_136) ) ;
    buf_clk cell_95 ( .C (clk), .D (signal_137), .Q (signal_138) ) ;
    buf_clk cell_97 ( .C (clk), .D (signal_139), .Q (signal_140) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_136, signal_134}), .Q ({Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_140, signal_138}), .Q ({Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_83, signal_33}), .Q ({Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_84, signal_34}), .Q ({Y_s1[0], Y_s0[0]}) ) ;
endmodule
