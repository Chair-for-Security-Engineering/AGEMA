/* modified netlist. Source: module sbox in file Designs/AESSbox//lookup/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 34 time(s)  */

module sbox_HPC2_AIG_ClockGating_d1 (SI_s0, clk, SI_s1, Fresh, rst, SO_s0, SO_s1, Synch);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input rst ;
    input [878:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output Synch ;
    wire signal_23 ;
    wire signal_24 ;
    wire signal_25 ;
    wire signal_26 ;
    wire signal_27 ;
    wire signal_28 ;
    wire signal_29 ;
    wire signal_30 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;
    wire signal_1069 ;
    wire signal_1070 ;
    wire signal_1071 ;
    wire signal_1072 ;
    wire signal_1073 ;
    wire signal_1074 ;
    wire signal_1075 ;
    wire signal_1076 ;
    wire signal_1077 ;
    wire signal_1078 ;
    wire signal_1079 ;
    wire signal_1080 ;
    wire signal_1081 ;
    wire signal_1082 ;
    wire signal_1083 ;
    wire signal_1084 ;
    wire signal_1085 ;
    wire signal_1086 ;
    wire signal_1087 ;
    wire signal_1088 ;
    wire signal_1089 ;
    wire signal_1090 ;
    wire signal_1091 ;
    wire signal_1092 ;
    wire signal_1093 ;
    wire signal_1094 ;
    wire signal_1095 ;
    wire signal_1096 ;
    wire signal_1097 ;
    wire signal_1098 ;
    wire signal_1099 ;
    wire signal_1100 ;
    wire signal_1101 ;
    wire signal_1102 ;
    wire signal_1103 ;
    wire signal_1104 ;
    wire signal_1105 ;
    wire signal_1106 ;
    wire signal_1107 ;
    wire signal_1108 ;
    wire signal_1109 ;
    wire signal_1110 ;
    wire signal_1111 ;
    wire signal_1112 ;
    wire signal_1113 ;
    wire signal_1114 ;
    wire signal_1115 ;
    wire signal_1116 ;
    wire signal_1117 ;
    wire signal_1118 ;
    wire signal_1119 ;
    wire signal_1120 ;
    wire signal_1121 ;
    wire signal_1122 ;
    wire signal_1123 ;
    wire signal_1124 ;
    wire signal_1125 ;
    wire signal_1126 ;
    wire signal_1127 ;
    wire signal_1128 ;
    wire signal_1129 ;
    wire signal_1130 ;
    wire signal_1131 ;
    wire signal_1132 ;
    wire signal_1133 ;
    wire signal_1134 ;
    wire signal_1135 ;
    wire signal_1136 ;
    wire signal_1137 ;
    wire signal_1138 ;
    wire signal_1139 ;
    wire signal_1140 ;
    wire signal_1141 ;
    wire signal_1142 ;
    wire signal_1143 ;
    wire signal_1144 ;
    wire signal_1145 ;
    wire signal_1146 ;
    wire signal_1147 ;
    wire signal_1148 ;
    wire signal_1149 ;
    wire signal_1150 ;
    wire signal_1151 ;
    wire signal_1152 ;
    wire signal_1153 ;
    wire signal_1154 ;
    wire signal_1155 ;
    wire signal_1156 ;
    wire signal_1157 ;
    wire signal_1158 ;
    wire signal_1159 ;
    wire signal_1160 ;
    wire signal_1161 ;
    wire signal_1162 ;
    wire signal_1163 ;
    wire signal_1164 ;
    wire signal_1165 ;
    wire signal_1166 ;
    wire signal_1167 ;
    wire signal_1168 ;
    wire signal_1169 ;
    wire signal_1170 ;
    wire signal_1171 ;
    wire signal_1172 ;
    wire signal_1173 ;
    wire signal_1174 ;
    wire signal_1175 ;
    wire signal_1176 ;
    wire signal_1177 ;
    wire signal_1178 ;
    wire signal_1179 ;
    wire signal_1180 ;
    wire signal_1181 ;
    wire signal_1182 ;
    wire signal_1183 ;
    wire signal_1184 ;
    wire signal_1185 ;
    wire signal_1186 ;
    wire signal_1187 ;
    wire signal_1188 ;
    wire signal_1189 ;
    wire signal_1190 ;
    wire signal_1191 ;
    wire signal_1192 ;
    wire signal_1193 ;
    wire signal_1194 ;
    wire signal_1195 ;
    wire signal_1196 ;
    wire signal_1197 ;
    wire signal_1198 ;
    wire signal_1199 ;
    wire signal_1200 ;
    wire signal_1201 ;
    wire signal_1202 ;
    wire signal_1203 ;
    wire signal_1204 ;
    wire signal_1205 ;
    wire signal_1206 ;
    wire signal_1207 ;
    wire signal_1208 ;
    wire signal_1209 ;
    wire signal_1210 ;
    wire signal_1211 ;
    wire signal_1212 ;
    wire signal_1213 ;
    wire signal_1214 ;
    wire signal_1215 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1228 ;
    wire signal_1229 ;
    wire signal_1230 ;
    wire signal_1231 ;
    wire signal_1232 ;
    wire signal_1233 ;
    wire signal_1234 ;
    wire signal_1235 ;
    wire signal_1236 ;
    wire signal_1237 ;
    wire signal_1238 ;
    wire signal_1239 ;
    wire signal_1240 ;
    wire signal_1241 ;
    wire signal_1242 ;
    wire signal_1243 ;
    wire signal_1244 ;
    wire signal_1245 ;
    wire signal_1246 ;
    wire signal_1247 ;
    wire signal_1248 ;
    wire signal_1249 ;
    wire signal_1250 ;
    wire signal_1251 ;
    wire signal_1252 ;
    wire signal_1253 ;
    wire signal_1254 ;
    wire signal_1255 ;
    wire signal_1256 ;
    wire signal_1257 ;
    wire signal_1258 ;
    wire signal_1259 ;
    wire signal_1260 ;
    wire signal_1261 ;
    wire signal_1262 ;
    wire signal_1263 ;
    wire signal_1264 ;
    wire signal_1265 ;
    wire signal_1266 ;
    wire signal_1267 ;
    wire signal_1268 ;
    wire signal_1269 ;
    wire signal_1270 ;
    wire signal_1271 ;
    wire signal_1272 ;
    wire signal_1273 ;
    wire signal_1274 ;
    wire signal_1275 ;
    wire signal_1276 ;
    wire signal_1277 ;
    wire signal_1278 ;
    wire signal_1279 ;
    wire signal_1280 ;
    wire signal_1281 ;
    wire signal_1282 ;
    wire signal_1283 ;
    wire signal_1284 ;
    wire signal_1285 ;
    wire signal_1286 ;
    wire signal_1287 ;
    wire signal_1288 ;
    wire signal_1289 ;
    wire signal_1290 ;
    wire signal_1291 ;
    wire signal_1292 ;
    wire signal_1293 ;
    wire signal_1294 ;
    wire signal_1295 ;
    wire signal_1296 ;
    wire signal_1297 ;
    wire signal_1298 ;
    wire signal_1299 ;
    wire signal_1300 ;
    wire signal_1301 ;
    wire signal_1302 ;
    wire signal_1303 ;
    wire signal_1304 ;
    wire signal_1305 ;
    wire signal_1306 ;
    wire signal_1307 ;
    wire signal_1308 ;
    wire signal_1309 ;
    wire signal_1310 ;
    wire signal_1311 ;
    wire signal_1312 ;
    wire signal_1313 ;
    wire signal_1314 ;
    wire signal_1315 ;
    wire signal_1316 ;
    wire signal_1317 ;
    wire signal_1318 ;
    wire signal_1319 ;
    wire signal_1320 ;
    wire signal_1321 ;
    wire signal_1322 ;
    wire signal_1323 ;
    wire signal_1324 ;
    wire signal_1325 ;
    wire signal_1326 ;
    wire signal_1327 ;
    wire signal_1328 ;
    wire signal_1329 ;
    wire signal_1330 ;
    wire signal_1331 ;
    wire signal_1332 ;
    wire signal_1333 ;
    wire signal_1334 ;
    wire signal_1335 ;
    wire signal_1336 ;
    wire signal_1337 ;
    wire signal_1338 ;
    wire signal_1339 ;
    wire signal_1340 ;
    wire signal_1341 ;
    wire signal_1342 ;
    wire signal_1343 ;
    wire signal_1344 ;
    wire signal_1345 ;
    wire signal_1346 ;
    wire signal_1347 ;
    wire signal_1348 ;
    wire signal_1349 ;
    wire signal_1350 ;
    wire signal_1351 ;
    wire signal_1352 ;
    wire signal_1353 ;
    wire signal_1354 ;
    wire signal_1355 ;
    wire signal_1356 ;
    wire signal_1357 ;
    wire signal_1358 ;
    wire signal_1359 ;
    wire signal_1360 ;
    wire signal_1361 ;
    wire signal_1362 ;
    wire signal_1363 ;
    wire signal_1364 ;
    wire signal_1365 ;
    wire signal_1366 ;
    wire signal_1367 ;
    wire signal_1368 ;
    wire signal_1369 ;
    wire signal_1370 ;
    wire signal_1371 ;
    wire signal_1372 ;
    wire signal_1373 ;
    wire signal_1374 ;
    wire signal_1375 ;
    wire signal_1376 ;
    wire signal_1377 ;
    wire signal_1378 ;
    wire signal_1379 ;
    wire signal_1380 ;
    wire signal_1381 ;
    wire signal_1382 ;
    wire signal_1383 ;
    wire signal_1384 ;
    wire signal_1385 ;
    wire signal_1386 ;
    wire signal_1387 ;
    wire signal_1388 ;
    wire signal_1389 ;
    wire signal_1390 ;
    wire signal_1391 ;
    wire signal_1392 ;
    wire signal_1393 ;
    wire signal_1394 ;
    wire signal_1395 ;
    wire signal_1396 ;
    wire signal_1397 ;
    wire signal_1398 ;
    wire signal_1399 ;
    wire signal_1400 ;
    wire signal_1401 ;
    wire signal_1402 ;
    wire signal_1403 ;
    wire signal_1404 ;
    wire signal_1405 ;
    wire signal_1406 ;
    wire signal_1407 ;
    wire signal_1408 ;
    wire signal_1409 ;
    wire signal_1410 ;
    wire signal_1411 ;
    wire signal_1412 ;
    wire signal_1413 ;
    wire signal_1414 ;
    wire signal_1415 ;
    wire signal_1416 ;
    wire signal_1417 ;
    wire signal_1418 ;
    wire signal_1419 ;
    wire signal_1420 ;
    wire signal_1421 ;
    wire signal_1422 ;
    wire signal_1423 ;
    wire signal_1424 ;
    wire signal_1425 ;
    wire signal_1426 ;
    wire signal_1427 ;
    wire signal_1428 ;
    wire signal_1429 ;
    wire signal_1430 ;
    wire signal_1431 ;
    wire signal_1432 ;
    wire signal_1433 ;
    wire signal_1434 ;
    wire signal_1435 ;
    wire signal_1436 ;
    wire signal_1437 ;
    wire signal_1438 ;
    wire signal_1439 ;
    wire signal_1440 ;
    wire signal_1441 ;
    wire signal_1442 ;
    wire signal_1443 ;
    wire signal_1444 ;
    wire signal_1445 ;
    wire signal_1446 ;
    wire signal_1447 ;
    wire signal_1448 ;
    wire signal_1449 ;
    wire signal_1450 ;
    wire signal_1451 ;
    wire signal_1452 ;
    wire signal_1453 ;
    wire signal_1454 ;
    wire signal_1455 ;
    wire signal_1456 ;
    wire signal_1457 ;
    wire signal_1458 ;
    wire signal_1459 ;
    wire signal_1460 ;
    wire signal_1461 ;
    wire signal_1462 ;
    wire signal_1463 ;
    wire signal_1464 ;
    wire signal_1465 ;
    wire signal_1466 ;
    wire signal_1467 ;
    wire signal_1468 ;
    wire signal_1469 ;
    wire signal_1470 ;
    wire signal_1471 ;
    wire signal_1472 ;
    wire signal_1473 ;
    wire signal_1474 ;
    wire signal_1475 ;
    wire signal_1476 ;
    wire signal_1477 ;
    wire signal_1478 ;
    wire signal_1479 ;
    wire signal_1480 ;
    wire signal_1481 ;
    wire signal_1482 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1503 ;
    wire signal_1504 ;
    wire signal_1505 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1521 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1844 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2277 ;
    wire signal_2278 ;
    wire signal_2279 ;
    wire signal_2280 ;
    wire signal_2281 ;
    wire signal_2282 ;
    wire signal_2283 ;
    wire signal_2284 ;
    wire signal_2285 ;
    wire signal_2286 ;
    wire signal_2287 ;
    wire signal_2288 ;
    wire signal_2289 ;
    wire signal_2290 ;
    wire signal_2291 ;
    wire signal_2292 ;
    wire signal_2293 ;
    wire signal_2294 ;
    wire signal_2295 ;
    wire signal_2296 ;
    wire signal_2297 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2301 ;
    wire signal_2302 ;
    wire signal_2303 ;
    wire signal_2304 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2338 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2341 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2344 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2347 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2350 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2353 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2356 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2359 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2362 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2365 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2368 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2371 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2374 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2377 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2380 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2383 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2386 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2389 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2393 ;
    wire signal_2395 ;
    wire signal_2397 ;
    wire signal_2399 ;
    wire signal_2401 ;
    wire signal_2403 ;
    wire signal_2405 ;
    wire signal_2407 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2410 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2413 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2416 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2419 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2422 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2425 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2428 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2431 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2434 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2437 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2440 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2443 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2446 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2449 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2452 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2455 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2458 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2461 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2464 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2467 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2470 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2473 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2476 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2479 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2482 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2485 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2488 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2491 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2494 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2497 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2500 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2503 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2506 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2509 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2512 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2515 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2518 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2521 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2524 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2527 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2530 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2533 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2536 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2539 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2542 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2545 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2548 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2551 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2554 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2557 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2560 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2563 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2566 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2569 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2572 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2575 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2578 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2581 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2584 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2587 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2590 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2593 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2596 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2599 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2602 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2605 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2608 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2611 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2614 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2617 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2620 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2623 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2626 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2629 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2632 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2635 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2638 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2641 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2644 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2647 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2650 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2653 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2656 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2659 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2662 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2665 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2668 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2671 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2674 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2677 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2680 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2683 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2686 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2689 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2692 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2695 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2698 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2701 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2704 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2707 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2710 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2713 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2716 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2719 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2850 ;
    wire signal_2851 ;
    wire signal_2852 ;
    wire signal_2853 ;
    wire signal_2854 ;
    wire signal_2855 ;
    wire signal_2856 ;
    wire signal_2857 ;
    wire signal_2858 ;
    wire signal_2859 ;
    wire signal_2860 ;
    wire signal_2861 ;
    wire signal_2862 ;
    wire signal_2863 ;
    wire signal_2864 ;
    wire signal_2865 ;
    wire signal_2866 ;
    wire signal_2867 ;
    wire signal_2868 ;
    wire signal_2869 ;
    wire signal_2870 ;
    wire signal_2871 ;
    wire signal_2872 ;
    wire signal_2873 ;
    wire signal_2874 ;
    wire signal_2875 ;
    wire signal_2876 ;
    wire signal_2877 ;
    wire signal_2878 ;
    wire signal_2879 ;
    wire signal_2880 ;
    wire signal_2881 ;
    wire signal_2882 ;
    wire signal_2883 ;
    wire signal_2884 ;
    wire signal_2885 ;
    wire signal_2886 ;
    wire signal_2887 ;
    wire signal_2888 ;
    wire signal_2889 ;
    wire signal_2890 ;
    wire signal_2891 ;
    wire signal_2892 ;
    wire signal_2893 ;
    wire signal_2894 ;
    wire signal_2895 ;
    wire signal_2896 ;
    wire signal_2897 ;
    wire signal_2898 ;
    wire signal_2899 ;
    wire signal_2900 ;
    wire signal_2901 ;
    wire signal_2902 ;
    wire signal_2903 ;
    wire signal_2904 ;
    wire signal_2905 ;
    wire signal_2906 ;
    wire signal_2907 ;
    wire signal_2908 ;
    wire signal_2909 ;
    wire signal_2910 ;
    wire signal_2911 ;
    wire signal_2912 ;
    wire signal_2913 ;
    wire signal_2914 ;
    wire signal_2915 ;
    wire signal_2916 ;
    wire signal_2917 ;
    wire signal_2918 ;
    wire signal_2919 ;
    wire signal_2920 ;
    wire signal_2921 ;
    wire signal_2922 ;
    wire signal_2923 ;
    wire signal_2924 ;
    wire signal_2925 ;
    wire signal_2926 ;
    wire signal_2927 ;
    wire signal_2928 ;
    wire signal_2929 ;
    wire signal_2930 ;
    wire signal_2931 ;
    wire signal_2932 ;
    wire signal_2933 ;
    wire signal_2934 ;
    wire signal_2935 ;
    wire signal_2936 ;
    wire signal_2937 ;
    wire signal_2938 ;
    wire signal_2939 ;
    wire signal_2940 ;
    wire signal_2941 ;
    wire signal_2942 ;
    wire signal_2943 ;
    wire signal_2944 ;
    wire signal_2945 ;
    wire signal_2946 ;
    wire signal_2947 ;
    wire signal_2948 ;
    wire signal_2949 ;
    wire signal_2950 ;
    wire signal_2951 ;
    wire signal_2952 ;
    wire signal_2953 ;
    wire signal_2954 ;
    wire signal_2955 ;
    wire signal_2956 ;
    wire signal_2957 ;
    wire signal_2958 ;
    wire signal_2959 ;
    wire signal_2960 ;
    wire signal_2961 ;
    wire signal_2962 ;
    wire signal_2963 ;
    wire signal_2964 ;
    wire signal_2965 ;
    wire signal_2966 ;
    wire signal_2967 ;
    wire signal_2968 ;
    wire signal_2969 ;
    wire signal_2970 ;
    wire signal_2971 ;
    wire signal_2972 ;
    wire signal_2973 ;
    wire signal_2974 ;
    wire signal_2975 ;
    wire signal_2976 ;
    wire signal_2977 ;
    wire signal_2978 ;
    wire signal_2979 ;
    wire signal_2980 ;
    wire signal_2981 ;
    wire signal_2982 ;
    wire signal_2983 ;
    wire signal_2984 ;
    wire signal_2985 ;
    wire signal_2986 ;
    wire signal_2987 ;
    wire signal_2988 ;
    wire signal_2989 ;
    wire signal_2990 ;
    wire signal_2991 ;
    wire signal_2992 ;
    wire signal_2993 ;
    wire signal_2994 ;
    wire signal_2995 ;
    wire signal_2996 ;
    wire signal_2997 ;
    wire signal_2998 ;
    wire signal_2999 ;
    wire signal_3000 ;
    wire signal_3001 ;
    wire signal_3002 ;
    wire signal_3003 ;
    wire signal_3004 ;
    wire signal_3005 ;
    wire signal_3006 ;
    wire signal_3007 ;
    wire signal_3008 ;
    wire signal_3009 ;
    wire signal_3010 ;
    wire signal_3011 ;
    wire signal_3012 ;
    wire signal_3013 ;
    wire signal_3014 ;
    wire signal_3015 ;
    wire signal_3016 ;
    wire signal_3017 ;
    wire signal_3018 ;
    wire signal_3019 ;
    wire signal_3020 ;
    wire signal_3021 ;
    wire signal_3022 ;
    wire signal_3023 ;
    wire signal_3024 ;
    wire signal_3025 ;
    wire signal_3026 ;
    wire signal_3027 ;
    wire signal_3028 ;
    wire signal_3029 ;
    wire signal_3030 ;
    wire signal_3031 ;
    wire signal_3032 ;
    wire signal_3033 ;
    wire signal_3034 ;
    wire signal_3035 ;
    wire signal_3036 ;
    wire signal_3037 ;
    wire signal_3038 ;
    wire signal_3039 ;
    wire signal_3040 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3262 ;
    wire signal_3263 ;
    wire signal_3264 ;
    wire signal_3265 ;
    wire signal_3266 ;
    wire signal_3267 ;
    wire signal_3268 ;
    wire signal_3269 ;
    wire signal_3270 ;
    wire signal_3271 ;
    wire signal_3272 ;
    wire signal_3273 ;
    wire signal_3274 ;
    wire signal_3275 ;
    wire signal_3276 ;
    wire signal_3277 ;
    wire signal_3278 ;
    wire signal_3279 ;
    wire signal_3280 ;
    wire signal_3281 ;
    wire signal_3282 ;
    wire signal_3283 ;
    wire signal_3284 ;
    wire signal_3285 ;
    wire signal_3286 ;
    wire signal_3287 ;
    wire signal_3288 ;
    wire signal_3289 ;
    wire signal_3290 ;
    wire signal_3291 ;
    wire signal_3292 ;
    wire signal_3293 ;
    wire signal_3294 ;
    wire signal_3295 ;
    wire signal_3296 ;
    wire signal_3297 ;
    wire signal_3298 ;
    wire signal_3299 ;
    wire signal_3300 ;
    wire signal_3301 ;
    wire signal_3302 ;
    wire signal_3303 ;
    wire signal_3304 ;
    wire signal_3305 ;
    wire signal_3306 ;
    wire signal_3307 ;
    wire signal_3308 ;
    wire signal_3309 ;
    wire signal_3310 ;
    wire signal_3311 ;
    wire signal_3312 ;
    wire signal_3313 ;
    wire signal_3314 ;
    wire signal_3315 ;
    wire signal_3316 ;
    wire signal_3317 ;
    wire signal_3318 ;
    wire signal_3319 ;
    wire signal_3320 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3324 ;
    wire signal_3325 ;
    wire signal_3326 ;
    wire signal_3327 ;
    wire signal_3328 ;
    wire signal_3329 ;
    wire signal_3330 ;
    wire signal_3331 ;
    wire signal_3332 ;
    wire signal_3333 ;
    wire signal_3334 ;
    wire signal_3335 ;
    wire signal_3336 ;
    wire signal_3337 ;
    wire signal_3338 ;
    wire signal_3339 ;
    wire signal_3340 ;
    wire signal_3341 ;
    wire signal_3342 ;
    wire signal_3343 ;
    wire signal_3344 ;
    wire signal_3345 ;
    wire signal_3346 ;
    wire signal_3347 ;
    wire signal_3348 ;
    wire signal_3349 ;
    wire signal_3350 ;
    wire signal_3351 ;
    wire signal_3352 ;
    wire signal_3353 ;
    wire signal_3354 ;
    wire signal_3355 ;
    wire signal_3356 ;
    wire signal_3357 ;
    wire signal_3358 ;
    wire signal_3359 ;
    wire signal_3360 ;
    wire signal_3361 ;
    wire signal_3362 ;
    wire signal_3363 ;
    wire signal_3364 ;
    wire signal_3365 ;
    wire signal_3366 ;
    wire signal_3367 ;
    wire signal_3368 ;
    wire signal_3369 ;
    wire signal_3370 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3436 ;
    wire signal_3437 ;
    wire signal_3438 ;
    wire signal_3439 ;
    wire signal_3440 ;
    wire signal_3441 ;
    wire signal_3442 ;
    wire signal_3443 ;
    wire signal_3444 ;
    wire signal_3445 ;
    wire signal_3446 ;
    wire signal_3447 ;
    wire signal_3448 ;
    wire signal_3449 ;
    wire signal_3450 ;
    wire signal_3451 ;
    wire signal_3452 ;
    wire signal_3453 ;
    wire signal_3454 ;
    wire signal_3455 ;
    wire signal_3456 ;
    wire signal_3457 ;
    wire signal_3458 ;
    wire signal_3459 ;
    wire signal_3460 ;
    wire signal_3461 ;
    wire signal_3462 ;
    wire signal_3463 ;
    wire signal_3464 ;
    wire signal_3465 ;
    wire signal_3466 ;
    wire signal_3467 ;
    wire signal_3468 ;
    wire signal_3469 ;
    wire signal_3470 ;
    wire signal_3471 ;
    wire signal_3472 ;
    wire signal_3473 ;
    wire signal_3474 ;
    wire signal_3475 ;
    wire signal_3476 ;
    wire signal_3477 ;
    wire signal_3478 ;
    wire signal_3479 ;
    wire signal_3480 ;
    wire signal_3481 ;
    wire signal_3482 ;
    wire signal_3483 ;
    wire signal_3484 ;
    wire signal_3485 ;
    wire signal_3486 ;
    wire signal_3487 ;
    wire signal_3488 ;
    wire signal_3489 ;
    wire signal_3490 ;
    wire signal_3491 ;
    wire signal_3492 ;
    wire signal_3493 ;
    wire signal_3494 ;
    wire signal_3495 ;
    wire signal_3496 ;
    wire signal_3497 ;
    wire signal_3498 ;
    wire signal_3499 ;
    wire signal_3500 ;
    wire signal_3501 ;
    wire signal_3502 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3568 ;
    wire signal_3569 ;
    wire signal_3570 ;
    wire signal_3571 ;
    wire signal_3572 ;
    wire signal_3573 ;
    wire signal_3574 ;
    wire signal_3575 ;
    wire signal_3576 ;
    wire signal_3577 ;
    wire signal_3578 ;
    wire signal_3579 ;
    wire signal_3580 ;
    wire signal_3581 ;
    wire signal_3582 ;
    wire signal_3583 ;
    wire signal_3584 ;
    wire signal_3585 ;
    wire signal_3586 ;
    wire signal_3587 ;
    wire signal_3588 ;
    wire signal_3589 ;
    wire signal_3590 ;
    wire signal_3591 ;
    wire signal_3592 ;
    wire signal_3593 ;
    wire signal_3594 ;
    wire signal_3595 ;
    wire signal_3596 ;
    wire signal_3597 ;
    wire signal_3598 ;
    wire signal_3599 ;
    wire signal_3600 ;
    wire signal_3601 ;
    wire signal_3602 ;
    wire signal_3603 ;
    wire signal_3604 ;
    wire signal_3605 ;
    wire signal_3606 ;
    wire signal_3607 ;
    wire signal_3608 ;
    wire signal_3609 ;
    wire signal_3610 ;
    wire signal_3611 ;
    wire signal_3612 ;
    wire signal_3613 ;
    wire signal_3614 ;
    wire signal_3615 ;
    wire signal_3616 ;
    wire signal_3617 ;
    wire signal_3618 ;
    wire signal_3619 ;
    wire signal_3620 ;
    wire signal_3621 ;
    wire signal_3622 ;
    wire signal_3623 ;
    wire signal_3624 ;
    wire signal_3625 ;
    wire signal_3626 ;
    wire signal_3627 ;
    wire signal_3628 ;
    wire signal_3629 ;
    wire signal_3630 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3672 ;
    wire signal_3673 ;
    wire signal_3674 ;
    wire signal_3675 ;
    wire signal_3676 ;
    wire signal_3677 ;
    wire signal_3678 ;
    wire signal_3679 ;
    wire signal_3680 ;
    wire signal_3681 ;
    wire signal_3682 ;
    wire signal_3683 ;
    wire signal_3684 ;
    wire signal_3685 ;
    wire signal_3686 ;
    wire signal_3687 ;
    wire signal_3688 ;
    wire signal_3689 ;
    wire signal_3690 ;
    wire signal_3691 ;
    wire signal_3692 ;
    wire signal_3693 ;
    wire signal_3694 ;
    wire signal_3695 ;
    wire signal_3696 ;
    wire signal_3697 ;
    wire signal_3698 ;
    wire signal_3699 ;
    wire signal_3700 ;
    wire signal_3701 ;
    wire signal_3702 ;
    wire signal_3703 ;
    wire signal_3704 ;
    wire signal_3705 ;
    wire signal_3706 ;
    wire signal_3707 ;
    wire signal_3708 ;
    wire signal_3709 ;
    wire signal_3710 ;
    wire signal_3711 ;
    wire signal_3712 ;
    wire signal_3713 ;
    wire signal_3714 ;
    wire signal_3715 ;
    wire signal_3716 ;
    wire signal_3717 ;
    wire signal_3718 ;
    wire signal_3719 ;
    wire signal_3720 ;
    wire signal_3721 ;
    wire signal_3722 ;
    wire signal_3723 ;
    wire signal_3724 ;
    wire signal_3725 ;
    wire signal_3726 ;
    wire signal_3727 ;
    wire signal_3728 ;
    wire signal_3729 ;
    wire signal_3730 ;
    wire signal_3731 ;
    wire signal_3732 ;
    wire signal_3733 ;
    wire signal_3734 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3744 ;
    wire signal_3745 ;
    wire signal_3746 ;
    wire signal_3747 ;
    wire signal_3748 ;
    wire signal_3749 ;
    wire signal_3750 ;
    wire signal_3751 ;
    wire signal_3752 ;
    wire signal_3753 ;
    wire signal_3754 ;
    wire signal_3755 ;
    wire signal_3756 ;
    wire signal_3757 ;
    wire signal_3758 ;
    wire signal_3759 ;
    wire signal_3760 ;
    wire signal_3761 ;
    wire signal_3762 ;
    wire signal_3763 ;
    wire signal_3764 ;
    wire signal_3765 ;
    wire signal_3766 ;
    wire signal_3767 ;
    wire signal_3768 ;
    wire signal_3769 ;
    wire signal_3770 ;
    wire signal_3771 ;
    wire signal_3772 ;
    wire signal_3773 ;
    wire signal_3774 ;
    wire signal_3775 ;
    wire signal_3776 ;
    wire signal_3777 ;
    wire signal_3778 ;
    wire signal_3779 ;
    wire signal_3780 ;
    wire signal_3781 ;
    wire signal_3782 ;
    wire signal_3783 ;
    wire signal_3784 ;
    wire signal_3785 ;
    wire signal_3786 ;
    wire signal_3787 ;
    wire signal_3788 ;
    wire signal_3789 ;
    wire signal_3790 ;
    wire signal_3791 ;
    wire signal_3792 ;
    wire signal_3793 ;
    wire signal_3794 ;
    wire signal_3795 ;
    wire signal_3796 ;
    wire signal_3797 ;
    wire signal_3798 ;
    wire signal_3799 ;
    wire signal_3800 ;
    wire signal_3801 ;
    wire signal_3802 ;
    wire signal_3803 ;
    wire signal_3804 ;
    wire signal_3805 ;
    wire signal_3806 ;
    wire signal_3807 ;
    wire signal_3808 ;
    wire signal_3809 ;
    wire signal_3810 ;
    wire signal_3811 ;
    wire signal_3812 ;
    wire signal_3813 ;
    wire signal_3814 ;
    wire signal_3815 ;
    wire signal_3816 ;
    wire signal_3817 ;
    wire signal_3818 ;
    wire signal_3819 ;
    wire signal_3820 ;
    wire signal_3821 ;
    wire signal_3822 ;
    wire signal_3823 ;
    wire signal_3824 ;
    wire signal_3825 ;
    wire signal_3826 ;
    wire signal_3827 ;
    wire signal_3828 ;
    wire signal_3829 ;
    wire signal_3830 ;
    wire signal_3831 ;
    wire signal_3832 ;
    wire signal_3833 ;
    wire signal_3834 ;
    wire signal_3835 ;
    wire signal_3836 ;
    wire signal_3837 ;
    wire signal_3838 ;
    wire signal_3839 ;
    wire signal_3840 ;
    wire signal_3841 ;
    wire signal_3842 ;
    wire signal_3843 ;
    wire signal_3844 ;
    wire signal_3845 ;
    wire signal_3846 ;
    wire signal_3847 ;
    wire signal_3848 ;
    wire signal_3849 ;
    wire signal_3850 ;
    wire signal_3851 ;
    wire signal_3852 ;
    wire signal_3853 ;
    wire signal_3854 ;
    wire signal_3855 ;
    wire signal_3856 ;
    wire signal_3857 ;
    wire signal_4746 ;

    /* cells in depth 0 */
    not_masked #(.security_order(1), .pipeline(0)) cell_927 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2393, signal_942}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_928 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2395, signal_943}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_929 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2397, signal_944}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_930 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2399, signal_945}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_931 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2401, signal_946}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_932 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_2403, signal_947}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_933 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2405, signal_948}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_934 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2407, signal_949}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_949 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .c ({signal_2422, signal_964}) ) ;
    xor_HPC2 #(.security_order(1), .pipeline(0)) cell_950 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[0], SI_s0[0]}), .c ({signal_2423, signal_965}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_962 ( .a ({signal_2422, signal_964}), .b ({signal_2435, signal_977}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_963 ( .a ({signal_2423, signal_965}), .b ({signal_2436, signal_978}) ) ;
    ClockGatingController #(35) cell_2385 ( .clk ( clk ), .rst ( rst ), .GatedClk ( signal_4746 ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_935 ( .a ({SI_s1[3], SI_s0[3]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[0] ), .c ({signal_2408, signal_950}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_936 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ( Fresh[1] ), .c ({signal_2409, signal_951}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_937 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[2] ), .c ({signal_2410, signal_952}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_938 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[3] ), .c ({signal_2411, signal_953}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_939 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[4] ), .c ({signal_2412, signal_954}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_940 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[5] ), .c ({signal_2413, signal_955}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_941 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[6] ), .c ({signal_2414, signal_956}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_942 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[7] ), .c ({signal_2415, signal_957}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_943 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[8] ), .c ({signal_2416, signal_958}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_944 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[9] ), .c ({signal_2417, signal_959}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_945 ( .a ({SI_s1[3], SI_s0[3]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[10] ), .c ({signal_2418, signal_960}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_946 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[11] ), .c ({signal_2419, signal_961}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_947 ( .a ({SI_s1[1], SI_s0[1]}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[12] ), .c ({signal_2420, signal_962}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_948 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[13] ), .c ({signal_2421, signal_963}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_951 ( .a ({signal_2408, signal_950}), .b ({signal_2424, signal_966}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_952 ( .a ({signal_2409, signal_951}), .b ({signal_2425, signal_967}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_953 ( .a ({signal_2410, signal_952}), .b ({signal_2426, signal_968}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_954 ( .a ({signal_2411, signal_953}), .b ({signal_2427, signal_969}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_955 ( .a ({signal_2412, signal_954}), .b ({signal_2428, signal_970}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_956 ( .a ({signal_2414, signal_956}), .b ({signal_2429, signal_971}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_957 ( .a ({signal_2415, signal_957}), .b ({signal_2430, signal_972}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_958 ( .a ({signal_2417, signal_959}), .b ({signal_2431, signal_973}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_959 ( .a ({signal_2418, signal_960}), .b ({signal_2432, signal_974}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_960 ( .a ({signal_2419, signal_961}), .b ({signal_2433, signal_975}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_961 ( .a ({signal_2420, signal_962}), .b ({signal_2434, signal_976}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_964 ( .a ({signal_2395, signal_943}), .b ({signal_2397, signal_944}), .clk ( clk ), .r ( Fresh[14] ), .c ({signal_2437, signal_979}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_965 ( .a ({signal_2405, signal_948}), .b ({signal_2407, signal_949}), .clk ( clk ), .r ( Fresh[15] ), .c ({signal_2438, signal_980}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_966 ( .a ({signal_2399, signal_945}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[16] ), .c ({signal_2439, signal_981}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_967 ( .a ({signal_2397, signal_944}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[17] ), .c ({signal_2440, signal_982}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_968 ( .a ({signal_2397, signal_944}), .b ({signal_2399, signal_945}), .clk ( clk ), .r ( Fresh[18] ), .c ({signal_2441, signal_983}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_969 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2395, signal_943}), .clk ( clk ), .r ( Fresh[19] ), .c ({signal_2442, signal_984}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_970 ( .a ({signal_2393, signal_942}), .b ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ( Fresh[20] ), .c ({signal_2443, signal_985}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_971 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[21] ), .c ({signal_2444, signal_986}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_972 ( .a ({signal_2403, signal_947}), .b ({signal_2407, signal_949}), .clk ( clk ), .r ( Fresh[22] ), .c ({signal_2445, signal_987}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_973 ( .a ({signal_2403, signal_947}), .b ({signal_2405, signal_948}), .clk ( clk ), .r ( Fresh[23] ), .c ({signal_2446, signal_988}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_974 ( .a ({signal_2403, signal_947}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[24] ), .c ({signal_2447, signal_989}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_975 ( .a ({signal_2395, signal_943}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[25] ), .c ({signal_2448, signal_990}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_976 ( .a ({signal_2399, signal_945}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[26] ), .c ({signal_2449, signal_991}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_977 ( .a ({signal_2405, signal_948}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[27] ), .c ({signal_2450, signal_992}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_978 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2397, signal_944}), .clk ( clk ), .r ( Fresh[28] ), .c ({signal_2451, signal_993}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_979 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[29] ), .c ({signal_2452, signal_994}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_980 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2397, signal_944}), .clk ( clk ), .r ( Fresh[30] ), .c ({signal_2453, signal_995}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_981 ( .a ({signal_2397, signal_944}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[31] ), .c ({signal_2454, signal_996}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_982 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2403, signal_947}), .clk ( clk ), .r ( Fresh[32] ), .c ({signal_2455, signal_997}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_983 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2407, signal_949}), .clk ( clk ), .r ( Fresh[33] ), .c ({signal_2456, signal_998}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_984 ( .a ({signal_2393, signal_942}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[34] ), .c ({signal_2457, signal_999}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_985 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_2405, signal_948}), .clk ( clk ), .r ( Fresh[35] ), .c ({signal_2458, signal_1000}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_986 ( .a ({signal_2393, signal_942}), .b ({signal_2395, signal_943}), .clk ( clk ), .r ( Fresh[36] ), .c ({signal_2459, signal_1001}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_987 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2399, signal_945}), .clk ( clk ), .r ( Fresh[37] ), .c ({signal_2460, signal_1002}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_989 ( .a ({signal_2401, signal_946}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[38] ), .c ({signal_2462, signal_1004}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_990 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2399, signal_945}), .clk ( clk ), .r ( Fresh[39] ), .c ({signal_2463, signal_1005}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_991 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2403, signal_947}), .clk ( clk ), .r ( Fresh[40] ), .c ({signal_2464, signal_1006}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_992 ( .a ({signal_2397, signal_944}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[41] ), .c ({signal_2465, signal_1007}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_993 ( .a ({signal_2403, signal_947}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[42] ), .c ({signal_2466, signal_1008}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_994 ( .a ({signal_2401, signal_946}), .b ({signal_2403, signal_947}), .clk ( clk ), .r ( Fresh[43] ), .c ({signal_2467, signal_1009}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_995 ( .a ({signal_2393, signal_942}), .b ({signal_2397, signal_944}), .clk ( clk ), .r ( Fresh[44] ), .c ({signal_2468, signal_1010}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_996 ( .a ({signal_2397, signal_944}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[45] ), .c ({signal_2469, signal_1011}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_997 ( .a ({signal_2399, signal_945}), .b ({signal_2403, signal_947}), .clk ( clk ), .r ( Fresh[46] ), .c ({signal_2470, signal_1012}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_998 ( .a ({signal_2399, signal_945}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[47] ), .c ({signal_2471, signal_1013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1000 ( .a ({signal_2399, signal_945}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[48] ), .c ({signal_2473, signal_1015}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1001 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2405, signal_948}), .clk ( clk ), .r ( Fresh[49] ), .c ({signal_2474, signal_1016}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1002 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2401, signal_946}), .clk ( clk ), .r ( Fresh[50] ), .c ({signal_2475, signal_1017}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1003 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2407, signal_949}), .clk ( clk ), .r ( Fresh[51] ), .c ({signal_2476, signal_1018}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1016 ( .a ({signal_2437, signal_979}), .b ({signal_2489, signal_1031}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1017 ( .a ({signal_2438, signal_980}), .b ({signal_2490, signal_1032}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1018 ( .a ({signal_2441, signal_983}), .b ({signal_2491, signal_1033}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1019 ( .a ({signal_2442, signal_984}), .b ({signal_2492, signal_1034}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1020 ( .a ({signal_2444, signal_986}), .b ({signal_2493, signal_1035}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1021 ( .a ({signal_2445, signal_987}), .b ({signal_2494, signal_1036}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1022 ( .a ({signal_2446, signal_988}), .b ({signal_2495, signal_1037}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1023 ( .a ({signal_2447, signal_989}), .b ({signal_2496, signal_1038}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1024 ( .a ({signal_2448, signal_990}), .b ({signal_2497, signal_1039}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1025 ( .a ({signal_2449, signal_991}), .b ({signal_2498, signal_1040}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1026 ( .a ({signal_2450, signal_992}), .b ({signal_2499, signal_1041}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1027 ( .a ({signal_2451, signal_993}), .b ({signal_2500, signal_1042}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1028 ( .a ({signal_2453, signal_995}), .b ({signal_2501, signal_1043}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1029 ( .a ({signal_2454, signal_996}), .b ({signal_2502, signal_1044}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1030 ( .a ({signal_2455, signal_997}), .b ({signal_2503, signal_1045}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1031 ( .a ({signal_2456, signal_998}), .b ({signal_2504, signal_1046}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1032 ( .a ({signal_2458, signal_1000}), .b ({signal_2505, signal_1047}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1034 ( .a ({signal_2462, signal_1004}), .b ({signal_2507, signal_1049}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1035 ( .a ({signal_2463, signal_1005}), .b ({signal_2508, signal_1050}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1036 ( .a ({signal_2464, signal_1006}), .b ({signal_2509, signal_1051}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1037 ( .a ({signal_2466, signal_1008}), .b ({signal_2510, signal_1052}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1038 ( .a ({signal_2467, signal_1009}), .b ({signal_2511, signal_1053}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1039 ( .a ({signal_2471, signal_1013}), .b ({signal_2512, signal_1054}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1041 ( .a ({signal_2473, signal_1015}), .b ({signal_2514, signal_1056}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1042 ( .a ({signal_2474, signal_1016}), .b ({signal_2515, signal_1057}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1043 ( .a ({signal_2475, signal_1017}), .b ({signal_2516, signal_1058}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_988 ( .a ({signal_2409, signal_951}), .b ({signal_2411, signal_953}), .clk ( clk ), .r ( Fresh[52] ), .c ({signal_2461, signal_1003}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_999 ( .a ({signal_2410, signal_952}), .b ({signal_2413, signal_955}), .clk ( clk ), .r ( Fresh[53] ), .c ({signal_2472, signal_1014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1004 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2411, signal_953}), .clk ( clk ), .r ( Fresh[54] ), .c ({signal_2477, signal_1019}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1005 ( .a ({signal_2409, signal_951}), .b ({signal_2416, signal_958}), .clk ( clk ), .r ( Fresh[55] ), .c ({signal_2478, signal_1020}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1006 ( .a ({signal_2407, signal_949}), .b ({signal_2411, signal_953}), .clk ( clk ), .r ( Fresh[56] ), .c ({signal_2479, signal_1021}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1007 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2418, signal_960}), .clk ( clk ), .r ( Fresh[57] ), .c ({signal_2480, signal_1022}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1008 ( .a ({signal_2415, signal_957}), .b ({signal_2417, signal_959}), .clk ( clk ), .r ( Fresh[58] ), .c ({signal_2481, signal_1023}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1009 ( .a ({signal_2409, signal_951}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[59] ), .c ({signal_2482, signal_1024}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1010 ( .a ({signal_2409, signal_951}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[60] ), .c ({signal_2483, signal_1025}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1011 ( .a ({signal_2413, signal_955}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[61] ), .c ({signal_2484, signal_1026}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1012 ( .a ({signal_2411, signal_953}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[62] ), .c ({signal_2485, signal_1027}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1013 ( .a ({signal_2408, signal_950}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[63] ), .c ({signal_2486, signal_1028}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1014 ( .a ({signal_2397, signal_944}), .b ({signal_2418, signal_960}), .clk ( clk ), .r ( Fresh[64] ), .c ({signal_2487, signal_1029}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1015 ( .a ({signal_2414, signal_956}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[65] ), .c ({signal_2488, signal_1030}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1033 ( .a ({signal_2461, signal_1003}), .b ({signal_2506, signal_1048}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1040 ( .a ({signal_2472, signal_1014}), .b ({signal_2513, signal_1055}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1044 ( .a ({signal_2478, signal_1020}), .b ({signal_2517, signal_1059}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1045 ( .a ({signal_2481, signal_1023}), .b ({signal_2518, signal_1060}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1046 ( .a ({signal_2483, signal_1025}), .b ({signal_2519, signal_1061}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1047 ( .a ({signal_2484, signal_1026}), .b ({signal_2520, signal_1062}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1048 ( .a ({signal_2485, signal_1027}), .b ({signal_2521, signal_1063}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1049 ( .a ({signal_2486, signal_1028}), .b ({signal_2522, signal_1064}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1050 ( .a ({signal_2487, signal_1029}), .b ({signal_2523, signal_1065}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1051 ( .a ({signal_2488, signal_1030}), .b ({signal_2524, signal_1066}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1052 ( .a ({signal_2407, signal_949}), .b ({signal_2437, signal_979}), .clk ( clk ), .r ( Fresh[66] ), .c ({signal_2525, signal_1067}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1053 ( .a ({signal_2393, signal_942}), .b ({signal_2441, signal_983}), .clk ( clk ), .r ( Fresh[67] ), .c ({signal_2526, signal_1068}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1054 ( .a ({signal_2425, signal_967}), .b ({signal_2426, signal_968}), .clk ( clk ), .r ( Fresh[68] ), .c ({signal_2527, signal_1069}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1055 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2424, signal_966}), .clk ( clk ), .r ( Fresh[69] ), .c ({signal_2528, signal_1070}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1056 ( .a ({signal_2401, signal_946}), .b ({signal_2438, signal_980}), .clk ( clk ), .r ( Fresh[70] ), .c ({signal_2529, signal_1071}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1057 ( .a ({signal_2410, signal_952}), .b ({signal_2438, signal_980}), .clk ( clk ), .r ( Fresh[71] ), .c ({signal_2530, signal_1072}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1058 ( .a ({signal_2443, signal_985}), .b ({signal_2416, signal_958}), .clk ( clk ), .r ( Fresh[72] ), .c ({signal_2531, signal_1073}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1059 ( .a ({signal_2409, signal_951}), .b ({signal_2439, signal_981}), .clk ( clk ), .r ( Fresh[73] ), .c ({signal_2532, signal_1074}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1060 ( .a ({signal_2409, signal_951}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[74] ), .c ({signal_2533, signal_1075}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1061 ( .a ({signal_2452, signal_994}), .b ({signal_2457, signal_999}), .clk ( clk ), .r ( Fresh[75] ), .c ({signal_2534, signal_1076}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1062 ( .a ({signal_2393, signal_942}), .b ({signal_2437, signal_979}), .clk ( clk ), .r ( Fresh[76] ), .c ({signal_2535, signal_1077}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1063 ( .a ({signal_2441, signal_983}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[77] ), .c ({signal_2536, signal_1078}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1064 ( .a ({signal_2446, signal_988}), .b ({signal_2460, signal_1002}), .clk ( clk ), .r ( Fresh[78] ), .c ({signal_2537, signal_1079}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1065 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[79] ), .c ({signal_2538, signal_1080}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1066 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2462, signal_1004}), .clk ( clk ), .r ( Fresh[80] ), .c ({signal_2539, signal_1081}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1067 ( .a ({signal_2441, signal_983}), .b ({signal_2443, signal_985}), .clk ( clk ), .r ( Fresh[81] ), .c ({signal_2540, signal_1082}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1068 ( .a ({signal_2409, signal_951}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[82] ), .c ({signal_2541, signal_1083}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1069 ( .a ({signal_2409, signal_951}), .b ({signal_2441, signal_983}), .clk ( clk ), .r ( Fresh[83] ), .c ({signal_2542, signal_1084}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1070 ( .a ({signal_2442, signal_984}), .b ({signal_2456, signal_998}), .clk ( clk ), .r ( Fresh[84] ), .c ({signal_2543, signal_1085}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1071 ( .a ({signal_2410, signal_952}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[85] ), .c ({signal_2544, signal_1086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1072 ( .a ({signal_2458, signal_1000}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[86] ), .c ({signal_2545, signal_1087}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1073 ( .a ({signal_2438, signal_980}), .b ({signal_2442, signal_984}), .clk ( clk ), .r ( Fresh[87] ), .c ({signal_2546, signal_1088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1074 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[88] ), .c ({signal_2547, signal_1089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1075 ( .a ({signal_2411, signal_953}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[89] ), .c ({signal_2548, signal_1090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1076 ( .a ({signal_2442, signal_984}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[90] ), .c ({signal_2549, signal_1091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1077 ( .a ({signal_2409, signal_951}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[91] ), .c ({signal_2550, signal_1092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1078 ( .a ({signal_2437, signal_979}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[92] ), .c ({signal_2551, signal_1093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1079 ( .a ({signal_2408, signal_950}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[93] ), .c ({signal_2552, signal_1094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1080 ( .a ({signal_2442, signal_984}), .b ({signal_2416, signal_958}), .clk ( clk ), .r ( Fresh[94] ), .c ({signal_2553, signal_1095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1081 ( .a ({signal_2437, signal_979}), .b ({signal_2470, signal_1012}), .clk ( clk ), .r ( Fresh[95] ), .c ({signal_2554, signal_1096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1082 ( .a ({signal_2439, signal_981}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[96] ), .c ({signal_2555, signal_1097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1083 ( .a ({signal_2410, signal_952}), .b ({signal_2439, signal_981}), .clk ( clk ), .r ( Fresh[97] ), .c ({signal_2556, signal_1098}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1084 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[98] ), .c ({signal_2557, signal_1099}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1086 ( .a ({signal_2440, signal_982}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[99] ), .c ({signal_2559, signal_1101}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1087 ( .a ({signal_2409, signal_951}), .b ({signal_2440, signal_982}), .clk ( clk ), .r ( Fresh[100] ), .c ({signal_2560, signal_1102}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1088 ( .a ({signal_2411, signal_953}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[101] ), .c ({signal_2561, signal_1103}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1089 ( .a ({signal_2407, signal_949}), .b ({signal_2446, signal_988}), .clk ( clk ), .r ( Fresh[102] ), .c ({signal_2562, signal_1104}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1090 ( .a ({signal_2441, signal_983}), .b ({signal_2418, signal_960}), .clk ( clk ), .r ( Fresh[103] ), .c ({signal_2563, signal_1105}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1091 ( .a ({signal_2410, signal_952}), .b ({signal_2474, signal_1016}), .clk ( clk ), .r ( Fresh[104] ), .c ({signal_2564, signal_1106}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1092 ( .a ({signal_2393, signal_942}), .b ({signal_2462, signal_1004}), .clk ( clk ), .r ( Fresh[105] ), .c ({signal_2565, signal_1107}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1093 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2438, signal_980}), .clk ( clk ), .r ( Fresh[106] ), .c ({signal_2566, signal_1108}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1094 ( .a ({signal_2410, signal_952}), .b ({signal_2470, signal_1012}), .clk ( clk ), .r ( Fresh[107] ), .c ({signal_2567, signal_1109}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1095 ( .a ({signal_2448, signal_990}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[108] ), .c ({signal_2568, signal_1110}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1096 ( .a ({signal_2439, signal_981}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[109] ), .c ({signal_2569, signal_1111}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1097 ( .a ({signal_2419, signal_961}), .b ({signal_2471, signal_1013}), .clk ( clk ), .r ( Fresh[110] ), .c ({signal_2570, signal_1112}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1098 ( .a ({signal_2439, signal_981}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[111] ), .c ({signal_2571, signal_1113}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1099 ( .a ({signal_2399, signal_945}), .b ({signal_2468, signal_1010}), .clk ( clk ), .r ( Fresh[112] ), .c ({signal_2572, signal_1114}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1100 ( .a ({signal_2401, signal_946}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[113] ), .c ({signal_2573, signal_1115}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1101 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2468, signal_1010}), .clk ( clk ), .r ( Fresh[114] ), .c ({signal_2574, signal_1116}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1102 ( .a ({signal_2444, signal_986}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[115] ), .c ({signal_2575, signal_1117}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1103 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2460, signal_1002}), .clk ( clk ), .r ( Fresh[116] ), .c ({signal_2576, signal_1118}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1104 ( .a ({signal_2439, signal_981}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[117] ), .c ({signal_2577, signal_1119}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1105 ( .a ({signal_2405, signal_948}), .b ({signal_2441, signal_983}), .clk ( clk ), .r ( Fresh[118] ), .c ({signal_2578, signal_1120}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1106 ( .a ({signal_2447, signal_989}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[119] ), .c ({signal_2579, signal_1121}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1107 ( .a ({signal_2418, signal_960}), .b ({signal_2476, signal_1018}), .clk ( clk ), .r ( Fresh[120] ), .c ({signal_2580, signal_1122}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1108 ( .a ({signal_2463, signal_1005}), .b ({signal_2466, signal_1008}), .clk ( clk ), .r ( Fresh[121] ), .c ({signal_2581, signal_1123}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1109 ( .a ({signal_2438, signal_980}), .b ({signal_2457, signal_999}), .clk ( clk ), .r ( Fresh[122] ), .c ({signal_2582, signal_1124}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1110 ( .a ({signal_2439, signal_981}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[123] ), .c ({signal_2583, signal_1125}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1111 ( .a ({signal_2444, signal_986}), .b ({signal_2466, signal_1008}), .clk ( clk ), .r ( Fresh[124] ), .c ({signal_2584, signal_1126}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1112 ( .a ({signal_2438, signal_980}), .b ({signal_2414, signal_956}), .clk ( clk ), .r ( Fresh[125] ), .c ({signal_2585, signal_1127}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1113 ( .a ({signal_2437, signal_979}), .b ({signal_2421, signal_963}), .clk ( clk ), .r ( Fresh[126] ), .c ({signal_2586, signal_1128}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1114 ( .a ({signal_2441, signal_983}), .b ({signal_2474, signal_1016}), .clk ( clk ), .r ( Fresh[127] ), .c ({signal_2587, signal_1129}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1115 ( .a ({signal_2412, signal_954}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[128] ), .c ({signal_2588, signal_1130}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1116 ( .a ({signal_2446, signal_988}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[129] ), .c ({signal_2589, signal_1131}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1117 ( .a ({signal_2409, signal_951}), .b ({signal_2444, signal_986}), .clk ( clk ), .r ( Fresh[130] ), .c ({signal_2590, signal_1132}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1118 ( .a ({signal_2447, signal_989}), .b ({signal_2448, signal_990}), .clk ( clk ), .r ( Fresh[131] ), .c ({signal_2591, signal_1133}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1119 ( .a ({signal_2448, signal_990}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[132] ), .c ({signal_2592, signal_1134}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1120 ( .a ({signal_2446, signal_988}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[133] ), .c ({signal_2593, signal_1135}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1121 ( .a ({signal_2448, signal_990}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[134] ), .c ({signal_2594, signal_1136}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1122 ( .a ({signal_2449, signal_991}), .b ({signal_2453, signal_995}), .clk ( clk ), .r ( Fresh[135] ), .c ({signal_2595, signal_1137}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1123 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[136] ), .c ({signal_2596, signal_1138}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1125 ( .a ({signal_2440, signal_982}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[137] ), .c ({signal_2598, signal_1140}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1126 ( .a ({signal_2415, signal_957}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[138] ), .c ({signal_2599, signal_1141}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1127 ( .a ({signal_2416, signal_958}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[139] ), .c ({signal_2600, signal_1142}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1128 ( .a ({signal_2459, signal_1001}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[140] ), .c ({signal_2601, signal_1143}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1129 ( .a ({signal_2442, signal_984}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[141] ), .c ({signal_2602, signal_1144}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1130 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[142] ), .c ({signal_2603, signal_1145}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1131 ( .a ({signal_2450, signal_992}), .b ({signal_2464, signal_1006}), .clk ( clk ), .r ( Fresh[143] ), .c ({signal_2604, signal_1146}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1133 ( .a ({signal_2412, signal_954}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[144] ), .c ({signal_2606, signal_1148}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1134 ( .a ({signal_2447, signal_989}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[145] ), .c ({signal_2607, signal_1149}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1135 ( .a ({signal_2462, signal_1004}), .b ({signal_2420, signal_962}), .clk ( clk ), .r ( Fresh[146] ), .c ({signal_2608, signal_1150}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1136 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2466, signal_1008}), .clk ( clk ), .r ( Fresh[147] ), .c ({signal_2609, signal_1151}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1137 ( .a ({signal_2463, signal_1005}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[148] ), .c ({signal_2610, signal_1152}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1138 ( .a ({signal_2407, signal_949}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[149] ), .c ({signal_2611, signal_1153}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1139 ( .a ({signal_2411, signal_953}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[150] ), .c ({signal_2612, signal_1154}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1141 ( .a ({signal_2458, signal_1000}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[151] ), .c ({signal_2614, signal_1156}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1142 ( .a ({signal_2449, signal_991}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[152] ), .c ({signal_2615, signal_1157}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1143 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2446, signal_988}), .clk ( clk ), .r ( Fresh[153] ), .c ({signal_2616, signal_1158}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1144 ( .a ({signal_2443, signal_985}), .b ({signal_2415, signal_957}), .clk ( clk ), .r ( Fresh[154] ), .c ({signal_2617, signal_1159}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1145 ( .a ({signal_2449, signal_991}), .b ({signal_2451, signal_993}), .clk ( clk ), .r ( Fresh[155] ), .c ({signal_2618, signal_1160}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1146 ( .a ({signal_2410, signal_952}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[156] ), .c ({signal_2619, signal_1161}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1147 ( .a ({signal_2443, signal_985}), .b ({signal_2454, signal_996}), .clk ( clk ), .r ( Fresh[157] ), .c ({signal_2620, signal_1162}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1148 ( .a ({signal_2424, signal_966}), .b ({signal_2431, signal_973}), .clk ( clk ), .r ( Fresh[158] ), .c ({signal_2621, signal_1163}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1149 ( .a ({signal_2446, signal_988}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[159] ), .c ({signal_2622, signal_1164}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1150 ( .a ({signal_2450, signal_992}), .b ({signal_2469, signal_1011}), .clk ( clk ), .r ( Fresh[160] ), .c ({signal_2623, signal_1165}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1151 ( .a ({signal_2440, signal_982}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[161] ), .c ({signal_2624, signal_1166}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1152 ( .a ({signal_2438, signal_980}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[162] ), .c ({signal_2625, signal_1167}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1153 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2452, signal_994}), .clk ( clk ), .r ( Fresh[163] ), .c ({signal_2626, signal_1168}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1154 ( .a ({signal_2415, signal_957}), .b ({signal_2468, signal_1010}), .clk ( clk ), .r ( Fresh[164] ), .c ({signal_2627, signal_1169}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1156 ( .a ({signal_2464, signal_1006}), .b ({signal_2468, signal_1010}), .clk ( clk ), .r ( Fresh[165] ), .c ({signal_2629, signal_1171}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1157 ( .a ({signal_2442, signal_984}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[166] ), .c ({signal_2630, signal_1172}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1158 ( .a ({signal_2455, signal_997}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[167] ), .c ({signal_2631, signal_1173}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1159 ( .a ({signal_2449, signal_991}), .b ({signal_2466, signal_1008}), .clk ( clk ), .r ( Fresh[168] ), .c ({signal_2632, signal_1174}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1160 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2446, signal_988}), .clk ( clk ), .r ( Fresh[169] ), .c ({signal_2633, signal_1175}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1161 ( .a ({signal_2401, signal_946}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[170] ), .c ({signal_2634, signal_1176}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1162 ( .a ({signal_2393, signal_942}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[171] ), .c ({signal_2635, signal_1177}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1163 ( .a ({signal_2453, signal_995}), .b ({signal_2473, signal_1015}), .clk ( clk ), .r ( Fresh[172] ), .c ({signal_2636, signal_1178}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1164 ( .a ({signal_2424, signal_966}), .b ({signal_2430, signal_972}), .clk ( clk ), .r ( Fresh[173] ), .c ({signal_2637, signal_1179}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1165 ( .a ({signal_2429, signal_971}), .b ({signal_2430, signal_972}), .clk ( clk ), .r ( Fresh[174] ), .c ({signal_2638, signal_1180}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1166 ( .a ({signal_2420, signal_962}), .b ({signal_2470, signal_1012}), .clk ( clk ), .r ( Fresh[175] ), .c ({signal_2639, signal_1181}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1167 ( .a ({signal_2438, signal_980}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[176] ), .c ({signal_2640, signal_1182}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1168 ( .a ({signal_2413, signal_955}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[177] ), .c ({signal_2641, signal_1183}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1169 ( .a ({signal_2397, signal_944}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[178] ), .c ({signal_2642, signal_1184}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1170 ( .a ({signal_2444, signal_986}), .b ({signal_2458, signal_1000}), .clk ( clk ), .r ( Fresh[179] ), .c ({signal_2643, signal_1185}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1171 ( .a ({signal_2420, signal_962}), .b ({signal_2473, signal_1015}), .clk ( clk ), .r ( Fresh[180] ), .c ({signal_2644, signal_1186}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1172 ( .a ({signal_2446, signal_988}), .b ({signal_2453, signal_995}), .clk ( clk ), .r ( Fresh[181] ), .c ({signal_2645, signal_1187}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1174 ( .a ({signal_2441, signal_983}), .b ({signal_2442, signal_984}), .clk ( clk ), .r ( Fresh[182] ), .c ({signal_2647, signal_1189}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1175 ( .a ({signal_2441, signal_983}), .b ({signal_2462, signal_1004}), .clk ( clk ), .r ( Fresh[183] ), .c ({signal_2648, signal_1190}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1176 ( .a ({signal_2409, signal_951}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[184] ), .c ({signal_2649, signal_1191}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1177 ( .a ({signal_2454, signal_996}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[185] ), .c ({signal_2650, signal_1192}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1178 ( .a ({signal_2427, signal_969}), .b ({signal_2434, signal_976}), .clk ( clk ), .r ( Fresh[186] ), .c ({signal_2651, signal_1193}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1179 ( .a ({signal_2411, signal_953}), .b ({signal_2449, signal_991}), .clk ( clk ), .r ( Fresh[187] ), .c ({signal_2652, signal_1194}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1180 ( .a ({signal_2445, signal_987}), .b ({signal_2415, signal_957}), .clk ( clk ), .r ( Fresh[188] ), .c ({signal_2653, signal_1195}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1181 ( .a ({signal_2420, signal_962}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[189] ), .c ({signal_2654, signal_1196}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1182 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[190] ), .c ({signal_2655, signal_1197}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1183 ( .a ({signal_2438, signal_980}), .b ({signal_2419, signal_961}), .clk ( clk ), .r ( Fresh[191] ), .c ({signal_2656, signal_1198}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1185 ( .a ({signal_2442, signal_984}), .b ({signal_2473, signal_1015}), .clk ( clk ), .r ( Fresh[192] ), .c ({signal_2658, signal_1200}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1186 ( .a ({signal_2456, signal_998}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[193] ), .c ({signal_2659, signal_1201}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1187 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2443, signal_985}), .clk ( clk ), .r ( Fresh[194] ), .c ({signal_2660, signal_1202}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1188 ( .a ({signal_2444, signal_986}), .b ({signal_2417, signal_959}), .clk ( clk ), .r ( Fresh[195] ), .c ({signal_2661, signal_1203}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1191 ( .a ({signal_2439, signal_981}), .b ({signal_2445, signal_987}), .clk ( clk ), .r ( Fresh[196] ), .c ({signal_2664, signal_1206}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1192 ( .a ({signal_2456, signal_998}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[197] ), .c ({signal_2665, signal_1207}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1193 ( .a ({signal_2415, signal_957}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[198] ), .c ({signal_2666, signal_1208}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1194 ( .a ({signal_2444, signal_986}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[199] ), .c ({signal_2667, signal_1209}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1195 ( .a ({signal_2446, signal_988}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[200] ), .c ({signal_2668, signal_1210}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1196 ( .a ({signal_2447, signal_989}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[201] ), .c ({signal_2669, signal_1211}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1197 ( .a ({signal_2443, signal_985}), .b ({signal_2444, signal_986}), .clk ( clk ), .r ( Fresh[202] ), .c ({signal_2670, signal_1212}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1199 ( .a ({signal_2449, signal_991}), .b ({signal_2450, signal_992}), .clk ( clk ), .r ( Fresh[203] ), .c ({signal_2672, signal_1214}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1200 ( .a ({signal_2411, signal_953}), .b ({signal_2465, signal_1007}), .clk ( clk ), .r ( Fresh[204] ), .c ({signal_2673, signal_1215}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1201 ( .a ({signal_2451, signal_993}), .b ({signal_2456, signal_998}), .clk ( clk ), .r ( Fresh[205] ), .c ({signal_2674, signal_1216}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1202 ( .a ({signal_2446, signal_988}), .b ({signal_2459, signal_1001}), .clk ( clk ), .r ( Fresh[206] ), .c ({signal_2675, signal_1217}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1203 ( .a ({signal_2453, signal_995}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[207] ), .c ({signal_2676, signal_1218}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1204 ( .a ({signal_2437, signal_979}), .b ({signal_2447, signal_989}), .clk ( clk ), .r ( Fresh[208] ), .c ({signal_2677, signal_1219}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1205 ( .a ({signal_2399, signal_945}), .b ({signal_2455, signal_997}), .clk ( clk ), .r ( Fresh[209] ), .c ({signal_2678, signal_1220}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1206 ( .a ({signal_2397, signal_944}), .b ({signal_2467, signal_1009}), .clk ( clk ), .r ( Fresh[210] ), .c ({signal_2679, signal_1221}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1208 ( .a ({signal_2462, signal_1004}), .b ({signal_2463, signal_1005}), .clk ( clk ), .r ( Fresh[211] ), .c ({signal_2681, signal_1223}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1210 ( .a ({signal_2405, signal_948}), .b ({signal_2428, signal_970}), .clk ( clk ), .r ( Fresh[212] ), .c ({signal_2683, signal_1225}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1213 ( .a ({signal_2437, signal_979}), .b ({signal_2436, signal_978}), .clk ( clk ), .r ( Fresh[213] ), .c ({signal_2686, signal_1228}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1214 ( .a ({signal_2405, signal_948}), .b ({signal_2430, signal_972}), .clk ( clk ), .r ( Fresh[214] ), .c ({signal_2687, signal_1229}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1215 ( .a ({signal_2527, signal_1069}), .b ({signal_2688, signal_1230}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1216 ( .a ({signal_2528, signal_1070}), .b ({signal_2689, signal_1231}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1217 ( .a ({signal_2530, signal_1072}), .b ({signal_2690, signal_1232}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1218 ( .a ({signal_2531, signal_1073}), .b ({signal_2691, signal_1233}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1219 ( .a ({signal_2532, signal_1074}), .b ({signal_2692, signal_1234}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1220 ( .a ({signal_2533, signal_1075}), .b ({signal_2693, signal_1235}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1221 ( .a ({signal_2534, signal_1076}), .b ({signal_2694, signal_1236}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1222 ( .a ({signal_2535, signal_1077}), .b ({signal_2695, signal_1237}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1223 ( .a ({signal_2536, signal_1078}), .b ({signal_2696, signal_1238}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1224 ( .a ({signal_2537, signal_1079}), .b ({signal_2697, signal_1239}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1225 ( .a ({signal_2538, signal_1080}), .b ({signal_2698, signal_1240}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1226 ( .a ({signal_2539, signal_1081}), .b ({signal_2699, signal_1241}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1227 ( .a ({signal_2540, signal_1082}), .b ({signal_2700, signal_1242}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1228 ( .a ({signal_2541, signal_1083}), .b ({signal_2701, signal_1243}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1229 ( .a ({signal_2542, signal_1084}), .b ({signal_2702, signal_1244}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1230 ( .a ({signal_2544, signal_1086}), .b ({signal_2703, signal_1245}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1231 ( .a ({signal_2545, signal_1087}), .b ({signal_2704, signal_1246}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1232 ( .a ({signal_2546, signal_1088}), .b ({signal_2705, signal_1247}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1233 ( .a ({signal_2548, signal_1090}), .b ({signal_2706, signal_1248}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1234 ( .a ({signal_2549, signal_1091}), .b ({signal_2707, signal_1249}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1235 ( .a ({signal_2550, signal_1092}), .b ({signal_2708, signal_1250}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1236 ( .a ({signal_2551, signal_1093}), .b ({signal_2709, signal_1251}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1237 ( .a ({signal_2552, signal_1094}), .b ({signal_2710, signal_1252}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1238 ( .a ({signal_2553, signal_1095}), .b ({signal_2711, signal_1253}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1239 ( .a ({signal_2554, signal_1096}), .b ({signal_2712, signal_1254}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1240 ( .a ({signal_2555, signal_1097}), .b ({signal_2713, signal_1255}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1241 ( .a ({signal_2556, signal_1098}), .b ({signal_2714, signal_1256}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1242 ( .a ({signal_2557, signal_1099}), .b ({signal_2715, signal_1257}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1244 ( .a ({signal_2559, signal_1101}), .b ({signal_2717, signal_1259}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1245 ( .a ({signal_2561, signal_1103}), .b ({signal_2718, signal_1260}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1246 ( .a ({signal_2563, signal_1105}), .b ({signal_2719, signal_1261}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1247 ( .a ({signal_2564, signal_1106}), .b ({signal_2720, signal_1262}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1248 ( .a ({signal_2566, signal_1108}), .b ({signal_2721, signal_1263}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1249 ( .a ({signal_2567, signal_1109}), .b ({signal_2722, signal_1264}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1250 ( .a ({signal_2568, signal_1110}), .b ({signal_2723, signal_1265}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1251 ( .a ({signal_2569, signal_1111}), .b ({signal_2724, signal_1266}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1252 ( .a ({signal_2570, signal_1112}), .b ({signal_2725, signal_1267}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1253 ( .a ({signal_2571, signal_1113}), .b ({signal_2726, signal_1268}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1254 ( .a ({signal_2573, signal_1115}), .b ({signal_2727, signal_1269}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1255 ( .a ({signal_2574, signal_1116}), .b ({signal_2728, signal_1270}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1256 ( .a ({signal_2575, signal_1117}), .b ({signal_2729, signal_1271}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1257 ( .a ({signal_2576, signal_1118}), .b ({signal_2730, signal_1272}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1258 ( .a ({signal_2578, signal_1120}), .b ({signal_2731, signal_1273}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1259 ( .a ({signal_2579, signal_1121}), .b ({signal_2732, signal_1274}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1260 ( .a ({signal_2580, signal_1122}), .b ({signal_2733, signal_1275}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1261 ( .a ({signal_2582, signal_1124}), .b ({signal_2734, signal_1276}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1262 ( .a ({signal_2583, signal_1125}), .b ({signal_2735, signal_1277}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1263 ( .a ({signal_2584, signal_1126}), .b ({signal_2736, signal_1278}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1264 ( .a ({signal_2585, signal_1127}), .b ({signal_2737, signal_1279}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1265 ( .a ({signal_2587, signal_1129}), .b ({signal_2738, signal_1280}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1266 ( .a ({signal_2588, signal_1130}), .b ({signal_2739, signal_1281}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1267 ( .a ({signal_2589, signal_1131}), .b ({signal_2740, signal_1282}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1268 ( .a ({signal_2592, signal_1134}), .b ({signal_2741, signal_1283}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1269 ( .a ({signal_2593, signal_1135}), .b ({signal_2742, signal_1284}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1270 ( .a ({signal_2594, signal_1136}), .b ({signal_2743, signal_1285}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1271 ( .a ({signal_2595, signal_1137}), .b ({signal_2744, signal_1286}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1273 ( .a ({signal_2599, signal_1141}), .b ({signal_2746, signal_1288}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1274 ( .a ({signal_2601, signal_1143}), .b ({signal_2747, signal_1289}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1275 ( .a ({signal_2602, signal_1144}), .b ({signal_2748, signal_1290}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1276 ( .a ({signal_2604, signal_1146}), .b ({signal_2749, signal_1291}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1278 ( .a ({signal_2606, signal_1148}), .b ({signal_2751, signal_1293}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1279 ( .a ({signal_2607, signal_1149}), .b ({signal_2752, signal_1294}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1280 ( .a ({signal_2608, signal_1150}), .b ({signal_2753, signal_1295}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1281 ( .a ({signal_2610, signal_1152}), .b ({signal_2754, signal_1296}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1282 ( .a ({signal_2611, signal_1153}), .b ({signal_2755, signal_1297}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1283 ( .a ({signal_2612, signal_1154}), .b ({signal_2756, signal_1298}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1285 ( .a ({signal_2614, signal_1156}), .b ({signal_2758, signal_1300}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1286 ( .a ({signal_2615, signal_1157}), .b ({signal_2759, signal_1301}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1287 ( .a ({signal_2617, signal_1159}), .b ({signal_2760, signal_1302}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1288 ( .a ({signal_2618, signal_1160}), .b ({signal_2761, signal_1303}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1289 ( .a ({signal_2619, signal_1161}), .b ({signal_2762, signal_1304}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1290 ( .a ({signal_2620, signal_1162}), .b ({signal_2763, signal_1305}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1291 ( .a ({signal_2621, signal_1163}), .b ({signal_2764, signal_1306}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1292 ( .a ({signal_2622, signal_1164}), .b ({signal_2765, signal_1307}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1293 ( .a ({signal_2623, signal_1165}), .b ({signal_2766, signal_1308}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1294 ( .a ({signal_2624, signal_1166}), .b ({signal_2767, signal_1309}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1295 ( .a ({signal_2625, signal_1167}), .b ({signal_2768, signal_1310}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1296 ( .a ({signal_2627, signal_1169}), .b ({signal_2769, signal_1311}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1298 ( .a ({signal_2629, signal_1171}), .b ({signal_2771, signal_1313}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1299 ( .a ({signal_2630, signal_1172}), .b ({signal_2772, signal_1314}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1300 ( .a ({signal_2631, signal_1173}), .b ({signal_2773, signal_1315}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1301 ( .a ({signal_2632, signal_1174}), .b ({signal_2774, signal_1316}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1302 ( .a ({signal_2633, signal_1175}), .b ({signal_2775, signal_1317}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1303 ( .a ({signal_2634, signal_1176}), .b ({signal_2776, signal_1318}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1304 ( .a ({signal_2635, signal_1177}), .b ({signal_2777, signal_1319}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1305 ( .a ({signal_2637, signal_1179}), .b ({signal_2778, signal_1320}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1306 ( .a ({signal_2638, signal_1180}), .b ({signal_2779, signal_1321}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1307 ( .a ({signal_2639, signal_1181}), .b ({signal_2780, signal_1322}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1308 ( .a ({signal_2640, signal_1182}), .b ({signal_2781, signal_1323}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1309 ( .a ({signal_2641, signal_1183}), .b ({signal_2782, signal_1324}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1310 ( .a ({signal_2642, signal_1184}), .b ({signal_2783, signal_1325}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1311 ( .a ({signal_2643, signal_1185}), .b ({signal_2784, signal_1326}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1312 ( .a ({signal_2644, signal_1186}), .b ({signal_2785, signal_1327}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1313 ( .a ({signal_2645, signal_1187}), .b ({signal_2786, signal_1328}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1315 ( .a ({signal_2647, signal_1189}), .b ({signal_2788, signal_1330}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1316 ( .a ({signal_2649, signal_1191}), .b ({signal_2789, signal_1331}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1317 ( .a ({signal_2650, signal_1192}), .b ({signal_2790, signal_1332}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1318 ( .a ({signal_2651, signal_1193}), .b ({signal_2791, signal_1333}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1319 ( .a ({signal_2652, signal_1194}), .b ({signal_2792, signal_1334}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1320 ( .a ({signal_2653, signal_1195}), .b ({signal_2793, signal_1335}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1321 ( .a ({signal_2654, signal_1196}), .b ({signal_2794, signal_1336}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1322 ( .a ({signal_2655, signal_1197}), .b ({signal_2795, signal_1337}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1324 ( .a ({signal_2658, signal_1200}), .b ({signal_2797, signal_1339}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1325 ( .a ({signal_2659, signal_1201}), .b ({signal_2798, signal_1340}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1326 ( .a ({signal_2660, signal_1202}), .b ({signal_2799, signal_1341}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1327 ( .a ({signal_2661, signal_1203}), .b ({signal_2800, signal_1342}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1330 ( .a ({signal_2665, signal_1207}), .b ({signal_2803, signal_1345}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1331 ( .a ({signal_2667, signal_1209}), .b ({signal_2804, signal_1346}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1332 ( .a ({signal_2668, signal_1210}), .b ({signal_2805, signal_1347}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1333 ( .a ({signal_2669, signal_1211}), .b ({signal_2806, signal_1348}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1334 ( .a ({signal_2670, signal_1212}), .b ({signal_2807, signal_1349}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1336 ( .a ({signal_2672, signal_1214}), .b ({signal_2809, signal_1351}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1337 ( .a ({signal_2673, signal_1215}), .b ({signal_2810, signal_1352}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1338 ( .a ({signal_2674, signal_1216}), .b ({signal_2811, signal_1353}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1339 ( .a ({signal_2676, signal_1218}), .b ({signal_2812, signal_1354}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1340 ( .a ({signal_2677, signal_1219}), .b ({signal_2813, signal_1355}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1341 ( .a ({signal_2678, signal_1220}), .b ({signal_2814, signal_1356}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1342 ( .a ({signal_2679, signal_1221}), .b ({signal_2815, signal_1357}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1344 ( .a ({signal_2681, signal_1223}), .b ({signal_2817, signal_1359}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1346 ( .a ({signal_2683, signal_1225}), .b ({signal_2819, signal_1361}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1349 ( .a ({signal_2686, signal_1228}), .b ({signal_2822, signal_1364}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1350 ( .a ({signal_2687, signal_1229}), .b ({signal_2823, signal_1365}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1353 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_2504, signal_1046}), .clk ( clk ), .r ( Fresh[215] ), .c ({signal_2826, signal_1368}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1354 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2500, signal_1042}), .clk ( clk ), .r ( Fresh[216] ), .c ({signal_2827, signal_1369}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1355 ( .a ({signal_2489, signal_1031}), .b ({signal_2516, signal_1058}), .clk ( clk ), .r ( Fresh[217] ), .c ({signal_2828, signal_1370}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1356 ( .a ({signal_2503, signal_1045}), .b ({signal_2515, signal_1057}), .clk ( clk ), .r ( Fresh[218] ), .c ({signal_2829, signal_1371}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1357 ( .a ({signal_2494, signal_1036}), .b ({signal_2495, signal_1037}), .clk ( clk ), .r ( Fresh[219] ), .c ({signal_2830, signal_1372}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1360 ( .a ({signal_2494, signal_1036}), .b ({signal_2503, signal_1045}), .clk ( clk ), .r ( Fresh[220] ), .c ({signal_2833, signal_1375}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1361 ( .a ({signal_2499, signal_1041}), .b ({signal_2510, signal_1052}), .clk ( clk ), .r ( Fresh[221] ), .c ({signal_2834, signal_1376}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1362 ( .a ({signal_2509, signal_1051}), .b ({signal_2511, signal_1053}), .clk ( clk ), .r ( Fresh[222] ), .c ({signal_2835, signal_1377}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1365 ( .a ({signal_2489, signal_1031}), .b ({signal_2502, signal_1044}), .clk ( clk ), .r ( Fresh[223] ), .c ({signal_2838, signal_1380}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1366 ( .a ({signal_2490, signal_1032}), .b ({signal_2510, signal_1052}), .clk ( clk ), .r ( Fresh[224] ), .c ({signal_2839, signal_1381}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1367 ( .a ({signal_2500, signal_1042}), .b ({signal_2501, signal_1043}), .clk ( clk ), .r ( Fresh[225] ), .c ({signal_2840, signal_1382}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1368 ( .a ({signal_2495, signal_1037}), .b ({signal_2503, signal_1045}), .clk ( clk ), .r ( Fresh[226] ), .c ({signal_2841, signal_1383}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1369 ( .a ({signal_2432, signal_974}), .b ({signal_2511, signal_1053}), .clk ( clk ), .r ( Fresh[227] ), .c ({signal_2842, signal_1384}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1375 ( .a ({signal_2498, signal_1040}), .b ({signal_2514, signal_1056}), .clk ( clk ), .r ( Fresh[228] ), .c ({signal_2848, signal_1390}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1376 ( .a ({signal_2503, signal_1045}), .b ({signal_2508, signal_1050}), .clk ( clk ), .r ( Fresh[229] ), .c ({signal_2849, signal_1391}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1383 ( .a ({signal_2491, signal_1033}), .b ({signal_2493, signal_1035}), .clk ( clk ), .r ( Fresh[230] ), .c ({signal_2856, signal_1398}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1395 ( .a ({signal_2429, signal_971}), .b ({signal_2507, signal_1049}), .clk ( clk ), .r ( Fresh[231] ), .c ({signal_2868, signal_1410}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1396 ( .a ({signal_2490, signal_1032}), .b ({signal_2505, signal_1047}), .clk ( clk ), .r ( Fresh[232] ), .c ({signal_2869, signal_1411}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1401 ( .a ({signal_2425, signal_967}), .b ({signal_2501, signal_1043}), .clk ( clk ), .r ( Fresh[233] ), .c ({signal_2874, signal_1416}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1402 ( .a ({signal_2508, signal_1050}), .b ({signal_2433, signal_975}), .clk ( clk ), .r ( Fresh[234] ), .c ({signal_2875, signal_1417}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1403 ( .a ({signal_2430, signal_972}), .b ({signal_2503, signal_1045}), .clk ( clk ), .r ( Fresh[235] ), .c ({signal_2876, signal_1418}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1407 ( .a ({signal_2496, signal_1038}), .b ({signal_2504, signal_1046}), .clk ( clk ), .r ( Fresh[236] ), .c ({signal_2880, signal_1422}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1408 ( .a ({signal_2498, signal_1040}), .b ({signal_2433, signal_975}), .clk ( clk ), .r ( Fresh[237] ), .c ({signal_2881, signal_1423}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1492 ( .a ({signal_2826, signal_1368}), .b ({signal_2965, signal_1507}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1493 ( .a ({signal_2827, signal_1369}), .b ({signal_2966, signal_1508}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1494 ( .a ({signal_2828, signal_1370}), .b ({signal_2967, signal_1509}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1495 ( .a ({signal_2829, signal_1371}), .b ({signal_2968, signal_1510}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1496 ( .a ({signal_2830, signal_1372}), .b ({signal_2969, signal_1511}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1499 ( .a ({signal_2833, signal_1375}), .b ({signal_2972, signal_1514}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1500 ( .a ({signal_2834, signal_1376}), .b ({signal_2973, signal_1515}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1501 ( .a ({signal_2835, signal_1377}), .b ({signal_2974, signal_1516}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1504 ( .a ({signal_2838, signal_1380}), .b ({signal_2977, signal_1519}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1505 ( .a ({signal_2839, signal_1381}), .b ({signal_2978, signal_1520}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1506 ( .a ({signal_2840, signal_1382}), .b ({signal_2979, signal_1521}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1507 ( .a ({signal_2842, signal_1384}), .b ({signal_2980, signal_1522}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1513 ( .a ({signal_2849, signal_1391}), .b ({signal_2986, signal_1528}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1520 ( .a ({signal_2856, signal_1398}), .b ({signal_2993, signal_1535}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1532 ( .a ({signal_2868, signal_1410}), .b ({signal_3005, signal_1547}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1533 ( .a ({signal_2869, signal_1411}), .b ({signal_3006, signal_1548}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1538 ( .a ({signal_2874, signal_1416}), .b ({signal_3011, signal_1553}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1539 ( .a ({signal_2875, signal_1417}), .b ({signal_3012, signal_1554}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1543 ( .a ({signal_2880, signal_1422}), .b ({signal_3016, signal_1558}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1544 ( .a ({signal_2881, signal_1423}), .b ({signal_3017, signal_1559}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1085 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2472, signal_1014}), .clk ( clk ), .r ( Fresh[238] ), .c ({signal_2558, signal_1100}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1124 ( .a ({signal_2399, signal_945}), .b ({signal_2477, signal_1019}), .clk ( clk ), .r ( Fresh[239] ), .c ({signal_2597, signal_1139}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1132 ( .a ({signal_2453, signal_995}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[240] ), .c ({signal_2605, signal_1147}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1140 ( .a ({signal_2468, signal_1010}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[241] ), .c ({signal_2613, signal_1155}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1155 ( .a ({signal_2450, signal_992}), .b ({signal_2478, signal_1020}), .clk ( clk ), .r ( Fresh[242] ), .c ({signal_2628, signal_1170}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1173 ( .a ({signal_2451, signal_993}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[243] ), .c ({signal_2646, signal_1188}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1184 ( .a ({signal_2466, signal_1008}), .b ({signal_2482, signal_1024}), .clk ( clk ), .r ( Fresh[244] ), .c ({signal_2657, signal_1199}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1189 ( .a ({signal_2449, signal_991}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[245] ), .c ({signal_2662, signal_1204}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1190 ( .a ({signal_2417, signal_959}), .b ({signal_2482, signal_1024}), .clk ( clk ), .r ( Fresh[246] ), .c ({signal_2663, signal_1205}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1198 ( .a ({signal_2445, signal_987}), .b ({signal_2482, signal_1024}), .clk ( clk ), .r ( Fresh[247] ), .c ({signal_2671, signal_1213}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1207 ( .a ({signal_2419, signal_961}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[248] ), .c ({signal_2680, signal_1222}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1209 ( .a ({signal_2437, signal_979}), .b ({signal_2484, signal_1026}), .clk ( clk ), .r ( Fresh[249] ), .c ({signal_2682, signal_1224}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1211 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2478, signal_1020}), .clk ( clk ), .r ( Fresh[250] ), .c ({signal_2684, signal_1226}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1212 ( .a ({signal_2418, signal_960}), .b ({signal_2478, signal_1020}), .clk ( clk ), .r ( Fresh[251] ), .c ({signal_2685, signal_1227}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1243 ( .a ({signal_2558, signal_1100}), .b ({signal_2716, signal_1258}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1272 ( .a ({signal_2597, signal_1139}), .b ({signal_2745, signal_1287}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1277 ( .a ({signal_2605, signal_1147}), .b ({signal_2750, signal_1292}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1284 ( .a ({signal_2613, signal_1155}), .b ({signal_2757, signal_1299}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1297 ( .a ({signal_2628, signal_1170}), .b ({signal_2770, signal_1312}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1314 ( .a ({signal_2646, signal_1188}), .b ({signal_2787, signal_1329}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1323 ( .a ({signal_2657, signal_1199}), .b ({signal_2796, signal_1338}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1328 ( .a ({signal_2662, signal_1204}), .b ({signal_2801, signal_1343}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1329 ( .a ({signal_2663, signal_1205}), .b ({signal_2802, signal_1344}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1335 ( .a ({signal_2671, signal_1213}), .b ({signal_2808, signal_1350}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1343 ( .a ({signal_2680, signal_1222}), .b ({signal_2816, signal_1358}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1345 ( .a ({signal_2682, signal_1224}), .b ({signal_2818, signal_1360}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1347 ( .a ({signal_2684, signal_1226}), .b ({signal_2820, signal_1362}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1348 ( .a ({signal_2685, signal_1227}), .b ({signal_2821, signal_1363}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1351 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_2525, signal_1067}), .clk ( clk ), .r ( Fresh[252] ), .c ({signal_2824, signal_1366}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1352 ( .a ({signal_2408, signal_950}), .b ({signal_2526, signal_1068}), .clk ( clk ), .r ( Fresh[253] ), .c ({signal_2825, signal_1367}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1358 ( .a ({signal_2451, signal_993}), .b ({signal_2538, signal_1080}), .clk ( clk ), .r ( Fresh[254] ), .c ({signal_2831, signal_1373}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1359 ( .a ({signal_2419, signal_961}), .b ({signal_2543, signal_1085}), .clk ( clk ), .r ( Fresh[255] ), .c ({signal_2832, signal_1374}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1363 ( .a ({signal_2417, signal_959}), .b ({signal_2547, signal_1089}), .clk ( clk ), .r ( Fresh[256] ), .c ({signal_2836, signal_1378}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1364 ( .a ({signal_2458, signal_1000}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[257] ), .c ({signal_2837, signal_1379}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1370 ( .a ({signal_2407, signal_949}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[258] ), .c ({signal_2843, signal_1385}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1371 ( .a ({signal_2401, signal_946}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[259] ), .c ({signal_2844, signal_1386}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1372 ( .a ({signal_2447, signal_989}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[260] ), .c ({signal_2845, signal_1387}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1373 ( .a ({signal_2531, signal_1073}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[261] ), .c ({signal_2846, signal_1388}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1374 ( .a ({signal_2405, signal_948}), .b ({signal_2555, signal_1097}), .clk ( clk ), .r ( Fresh[262] ), .c ({signal_2847, signal_1389}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1377 ( .a ({signal_2444, signal_986}), .b ({signal_2562, signal_1104}), .clk ( clk ), .r ( Fresh[263] ), .c ({signal_2850, signal_1392}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1378 ( .a ({signal_2490, signal_1032}), .b ({signal_2536, signal_1078}), .clk ( clk ), .r ( Fresh[264] ), .c ({signal_2851, signal_1393}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1379 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[265] ), .c ({signal_2852, signal_1394}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1380 ( .a ({signal_2405, signal_948}), .b ({signal_2547, signal_1089}), .clk ( clk ), .r ( Fresh[266] ), .c ({signal_2853, signal_1395}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1381 ( .a ({signal_2417, signal_959}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[267] ), .c ({signal_2854, signal_1396}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1382 ( .a ({signal_2474, signal_1016}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[268] ), .c ({signal_2855, signal_1397}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1384 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2565, signal_1107}), .clk ( clk ), .r ( Fresh[269] ), .c ({signal_2857, signal_1399}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1385 ( .a ({signal_2466, signal_1008}), .b ({signal_2550, signal_1092}), .clk ( clk ), .r ( Fresh[270] ), .c ({signal_2858, signal_1400}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1386 ( .a ({SI_s1[5], SI_s0[5]}), .b ({signal_2538, signal_1080}), .clk ( clk ), .r ( Fresh[271] ), .c ({signal_2859, signal_1401}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1387 ( .a ({signal_2420, signal_962}), .b ({signal_2544, signal_1086}), .clk ( clk ), .r ( Fresh[272] ), .c ({signal_2860, signal_1402}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1388 ( .a ({signal_2456, signal_998}), .b ({signal_2572, signal_1114}), .clk ( clk ), .r ( Fresh[273] ), .c ({signal_2861, signal_1403}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1389 ( .a ({signal_2459, signal_1001}), .b ({signal_2566, signal_1108}), .clk ( clk ), .r ( Fresh[274] ), .c ({signal_2862, signal_1404}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1390 ( .a ({signal_2407, signal_949}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[275] ), .c ({signal_2863, signal_1405}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1391 ( .a ({signal_2450, signal_992}), .b ({signal_2555, signal_1097}), .clk ( clk ), .r ( Fresh[276] ), .c ({signal_2864, signal_1406}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1392 ( .a ({signal_2456, signal_998}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[277] ), .c ({signal_2865, signal_1407}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1393 ( .a ({signal_2467, signal_1009}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[278] ), .c ({signal_2866, signal_1408}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1394 ( .a ({signal_2407, signal_949}), .b ({signal_2572, signal_1114}), .clk ( clk ), .r ( Fresh[279] ), .c ({signal_2867, signal_1409}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1397 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2560, signal_1102}), .clk ( clk ), .r ( Fresh[280] ), .c ({signal_2870, signal_1412}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1398 ( .a ({signal_2418, signal_960}), .b ({signal_2581, signal_1123}), .clk ( clk ), .r ( Fresh[281] ), .c ({signal_2871, signal_1413}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1399 ( .a ({signal_2411, signal_953}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[282] ), .c ({signal_2872, signal_1414}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1400 ( .a ({signal_2407, signal_949}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[283] ), .c ({signal_2873, signal_1415}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1404 ( .a ({signal_2447, signal_989}), .b ({signal_2536, signal_1078}), .clk ( clk ), .r ( Fresh[284] ), .c ({signal_2877, signal_1419}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1405 ( .a ({signal_2417, signal_959}), .b ({signal_2560, signal_1102}), .clk ( clk ), .r ( Fresh[285] ), .c ({signal_2878, signal_1420}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1406 ( .a ({signal_2446, signal_988}), .b ({signal_2573, signal_1115}), .clk ( clk ), .r ( Fresh[286] ), .c ({signal_2879, signal_1421}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1409 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[287] ), .c ({signal_2882, signal_1424}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1410 ( .a ({signal_2399, signal_945}), .b ({signal_2565, signal_1107}), .clk ( clk ), .r ( Fresh[288] ), .c ({signal_2883, signal_1425}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1411 ( .a ({signal_2447, signal_989}), .b ({signal_2544, signal_1086}), .clk ( clk ), .r ( Fresh[289] ), .c ({signal_2884, signal_1426}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1412 ( .a ({signal_2450, signal_992}), .b ({signal_2586, signal_1128}), .clk ( clk ), .r ( Fresh[290] ), .c ({signal_2885, signal_1427}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1413 ( .a ({signal_2462, signal_1004}), .b ({signal_2530, signal_1072}), .clk ( clk ), .r ( Fresh[291] ), .c ({signal_2886, signal_1428}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1414 ( .a ({signal_2415, signal_957}), .b ({signal_2591, signal_1133}), .clk ( clk ), .r ( Fresh[292] ), .c ({signal_2887, signal_1429}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1415 ( .a ({signal_2401, signal_946}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[293] ), .c ({signal_2888, signal_1430}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1416 ( .a ({signal_2395, signal_943}), .b ({signal_2596, signal_1138}), .clk ( clk ), .r ( Fresh[294] ), .c ({signal_2889, signal_1431}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1417 ( .a ({signal_2418, signal_960}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[295] ), .c ({signal_2890, signal_1432}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1418 ( .a ({signal_2442, signal_984}), .b ({signal_2598, signal_1140}), .clk ( clk ), .r ( Fresh[296] ), .c ({signal_2891, signal_1433}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1419 ( .a ({signal_2455, signal_997}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[297] ), .c ({signal_2892, signal_1434}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1420 ( .a ({signal_2408, signal_950}), .b ({signal_2600, signal_1142}), .clk ( clk ), .r ( Fresh[298] ), .c ({signal_2893, signal_1435}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1421 ( .a ({signal_2411, signal_953}), .b ({signal_2542, signal_1084}), .clk ( clk ), .r ( Fresh[299] ), .c ({signal_2894, signal_1436}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1422 ( .a ({signal_2408, signal_950}), .b ({signal_2533, signal_1075}), .clk ( clk ), .r ( Fresh[300] ), .c ({signal_2895, signal_1437}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1423 ( .a ({signal_2405, signal_948}), .b ({signal_2609, signal_1151}), .clk ( clk ), .r ( Fresh[301] ), .c ({signal_2896, signal_1438}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1424 ( .a ({signal_2465, signal_1007}), .b ({signal_2611, signal_1153}), .clk ( clk ), .r ( Fresh[302] ), .c ({signal_2897, signal_1439}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1425 ( .a ({signal_2407, signal_949}), .b ({signal_2614, signal_1156}), .clk ( clk ), .r ( Fresh[303] ), .c ({signal_2898, signal_1440}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1426 ( .a ({signal_2444, signal_986}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[304] ), .c ({signal_2899, signal_1441}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1427 ( .a ({signal_2408, signal_950}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[305] ), .c ({signal_2900, signal_1442}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1428 ( .a ({signal_2446, signal_988}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[306] ), .c ({signal_2901, signal_1443}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1429 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_2624, signal_1166}), .clk ( clk ), .r ( Fresh[307] ), .c ({signal_2902, signal_1444}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1430 ( .a ({signal_2544, signal_1086}), .b ({signal_2479, signal_1021}), .clk ( clk ), .r ( Fresh[308] ), .c ({signal_2903, signal_1445}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1431 ( .a ({signal_2409, signal_951}), .b ({signal_2626, signal_1168}), .clk ( clk ), .r ( Fresh[309] ), .c ({signal_2904, signal_1446}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1432 ( .a ({signal_2480, signal_1022}), .b ({signal_2600, signal_1142}), .clk ( clk ), .r ( Fresh[310] ), .c ({signal_2905, signal_1447}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1433 ( .a ({signal_2466, signal_1008}), .b ({signal_2594, signal_1136}), .clk ( clk ), .r ( Fresh[311] ), .c ({signal_2906, signal_1448}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1434 ( .a ({signal_2601, signal_1143}), .b ({signal_2603, signal_1145}), .clk ( clk ), .r ( Fresh[312] ), .c ({signal_2907, signal_1449}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1435 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2624, signal_1166}), .clk ( clk ), .r ( Fresh[313] ), .c ({signal_2908, signal_1450}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1436 ( .a ({signal_2439, signal_981}), .b ({signal_2611, signal_1153}), .clk ( clk ), .r ( Fresh[314] ), .c ({signal_2909, signal_1451}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1437 ( .a ({signal_2456, signal_998}), .b ({signal_2634, signal_1176}), .clk ( clk ), .r ( Fresh[315] ), .c ({signal_2910, signal_1452}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1438 ( .a ({signal_2594, signal_1136}), .b ({signal_2611, signal_1153}), .clk ( clk ), .r ( Fresh[316] ), .c ({signal_2911, signal_1453}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1439 ( .a ({signal_2549, signal_1091}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[317] ), .c ({signal_2912, signal_1454}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1440 ( .a ({signal_2437, signal_979}), .b ({signal_2615, signal_1157}), .clk ( clk ), .r ( Fresh[318] ), .c ({signal_2913, signal_1455}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1441 ( .a ({signal_2450, signal_992}), .b ({signal_2636, signal_1178}), .clk ( clk ), .r ( Fresh[319] ), .c ({signal_2914, signal_1456}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1442 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2540, signal_1082}), .clk ( clk ), .r ( Fresh[320] ), .c ({signal_2915, signal_1457}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1443 ( .a ({signal_2415, signal_957}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[321] ), .c ({signal_2916, signal_1458}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1444 ( .a ({signal_2405, signal_948}), .b ({signal_2541, signal_1083}), .clk ( clk ), .r ( Fresh[322] ), .c ({signal_2917, signal_1459}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1445 ( .a ({signal_2401, signal_946}), .b ({signal_2647, signal_1189}), .clk ( clk ), .r ( Fresh[323] ), .c ({signal_2918, signal_1460}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1446 ( .a ({SI_s1[6], SI_s0[6]}), .b ({signal_2648, signal_1190}), .clk ( clk ), .r ( Fresh[324] ), .c ({signal_2919, signal_1461}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1447 ( .a ({signal_2401, signal_946}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[325] ), .c ({signal_2920, signal_1462}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1448 ( .a ({signal_2448, signal_990}), .b ({signal_2615, signal_1157}), .clk ( clk ), .r ( Fresh[326] ), .c ({signal_2921, signal_1463}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1449 ( .a ({signal_2456, signal_998}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[327] ), .c ({signal_2922, signal_1464}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1450 ( .a ({signal_2465, signal_1007}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[328] ), .c ({signal_2923, signal_1465}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1451 ( .a ({signal_2464, signal_1006}), .b ({signal_2656, signal_1198}), .clk ( clk ), .r ( Fresh[329] ), .c ({signal_2924, signal_1466}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1452 ( .a ({signal_2441, signal_983}), .b ({signal_2603, signal_1145}), .clk ( clk ), .r ( Fresh[330] ), .c ({signal_2925, signal_1467}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1453 ( .a ({signal_2438, signal_980}), .b ({signal_2650, signal_1192}), .clk ( clk ), .r ( Fresh[331] ), .c ({signal_2926, signal_1468}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1454 ( .a ({signal_2560, signal_1102}), .b ({signal_2616, signal_1158}), .clk ( clk ), .r ( Fresh[332] ), .c ({signal_2927, signal_1469}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1455 ( .a ({signal_2450, signal_992}), .b ({signal_2635, signal_1177}), .clk ( clk ), .r ( Fresh[333] ), .c ({signal_2928, signal_1470}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1456 ( .a ({signal_2407, signal_949}), .b ({signal_2540, signal_1082}), .clk ( clk ), .r ( Fresh[334] ), .c ({signal_2929, signal_1471}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1457 ( .a ({signal_2446, signal_988}), .b ({signal_2649, signal_1191}), .clk ( clk ), .r ( Fresh[335] ), .c ({signal_2930, signal_1472}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1458 ( .a ({signal_2474, signal_1016}), .b ({signal_2602, signal_1144}), .clk ( clk ), .r ( Fresh[336] ), .c ({signal_2931, signal_1473}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1459 ( .a ({signal_2401, signal_946}), .b ({signal_2635, signal_1177}), .clk ( clk ), .r ( Fresh[337] ), .c ({signal_2932, signal_1474}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1460 ( .a ({signal_2459, signal_1001}), .b ({signal_2644, signal_1186}), .clk ( clk ), .r ( Fresh[338] ), .c ({signal_2933, signal_1475}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1461 ( .a ({signal_2447, signal_989}), .b ({signal_2542, signal_1084}), .clk ( clk ), .r ( Fresh[339] ), .c ({signal_2934, signal_1476}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1462 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2540, signal_1082}), .clk ( clk ), .r ( Fresh[340] ), .c ({signal_2935, signal_1477}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1463 ( .a ({signal_2405, signal_948}), .b ({signal_2664, signal_1206}), .clk ( clk ), .r ( Fresh[341] ), .c ({signal_2936, signal_1478}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1464 ( .a ({signal_2415, signal_957}), .b ({signal_2611, signal_1153}), .clk ( clk ), .r ( Fresh[342] ), .c ({signal_2937, signal_1479}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1465 ( .a ({signal_2451, signal_993}), .b ({signal_2644, signal_1186}), .clk ( clk ), .r ( Fresh[343] ), .c ({signal_2938, signal_1480}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1466 ( .a ({signal_2533, signal_1075}), .b ({signal_2539, signal_1081}), .clk ( clk ), .r ( Fresh[344] ), .c ({signal_2939, signal_1481}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1467 ( .a ({signal_2445, signal_987}), .b ({signal_2626, signal_1168}), .clk ( clk ), .r ( Fresh[345] ), .c ({signal_2940, signal_1482}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1468 ( .a ({signal_2446, signal_988}), .b ({signal_2619, signal_1161}), .clk ( clk ), .r ( Fresh[346] ), .c ({signal_2941, signal_1483}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1469 ( .a ({signal_2479, signal_1021}), .b ({signal_2590, signal_1132}), .clk ( clk ), .r ( Fresh[347] ), .c ({signal_2942, signal_1484}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1470 ( .a ({signal_2420, signal_962}), .b ({signal_2542, signal_1084}), .clk ( clk ), .r ( Fresh[348] ), .c ({signal_2943, signal_1485}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1471 ( .a ({signal_2457, signal_999}), .b ({signal_2666, signal_1208}), .clk ( clk ), .r ( Fresh[349] ), .c ({signal_2944, signal_1486}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1472 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2542, signal_1084}), .clk ( clk ), .r ( Fresh[350] ), .c ({signal_2945, signal_1487}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1473 ( .a ({signal_2474, signal_1016}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[351] ), .c ({signal_2946, signal_1488}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1474 ( .a ({signal_2430, signal_972}), .b ({signal_2659, signal_1201}), .clk ( clk ), .r ( Fresh[352] ), .c ({signal_2947, signal_1489}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1475 ( .a ({signal_2417, signal_959}), .b ({signal_2619, signal_1161}), .clk ( clk ), .r ( Fresh[353] ), .c ({signal_2948, signal_1490}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1476 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[354] ), .c ({signal_2949, signal_1491}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1477 ( .a ({signal_2415, signal_957}), .b ({signal_2675, signal_1217}), .clk ( clk ), .r ( Fresh[355] ), .c ({signal_2950, signal_1492}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1478 ( .a ({signal_2462, signal_1004}), .b ({signal_2553, signal_1095}), .clk ( clk ), .r ( Fresh[356] ), .c ({signal_2951, signal_1493}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1479 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2647, signal_1189}), .clk ( clk ), .r ( Fresh[357] ), .c ({signal_2952, signal_1494}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1480 ( .a ({signal_2434, signal_976}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[358] ), .c ({signal_2953, signal_1495}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1481 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2531, signal_1073}), .clk ( clk ), .r ( Fresh[359] ), .c ({signal_2954, signal_1496}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1482 ( .a ({signal_2405, signal_948}), .b ({signal_2602, signal_1144}), .clk ( clk ), .r ( Fresh[360] ), .c ({signal_2955, signal_1497}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1483 ( .a ({signal_2447, signal_989}), .b ({signal_2602, signal_1144}), .clk ( clk ), .r ( Fresh[361] ), .c ({signal_2956, signal_1498}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1484 ( .a ({signal_2418, signal_960}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[362] ), .c ({signal_2957, signal_1499}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1485 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[363] ), .c ({signal_2958, signal_1500}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1486 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2620, signal_1162}), .clk ( clk ), .r ( Fresh[364] ), .c ({signal_2959, signal_1501}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1487 ( .a ({signal_2407, signal_949}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[365] ), .c ({signal_2960, signal_1502}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1488 ( .a ({signal_2405, signal_948}), .b ({signal_2601, signal_1143}), .clk ( clk ), .r ( Fresh[366] ), .c ({signal_2961, signal_1503}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1489 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_2577, signal_1119}), .clk ( clk ), .r ( Fresh[367] ), .c ({signal_2962, signal_1504}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1490 ( .a ({signal_2824, signal_1366}), .b ({signal_2963, signal_1505}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1491 ( .a ({signal_2825, signal_1367}), .b ({signal_2964, signal_1506}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1497 ( .a ({signal_2831, signal_1373}), .b ({signal_2970, signal_1512}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1498 ( .a ({signal_2832, signal_1374}), .b ({signal_2971, signal_1513}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1502 ( .a ({signal_2836, signal_1378}), .b ({signal_2975, signal_1517}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1503 ( .a ({signal_2837, signal_1379}), .b ({signal_2976, signal_1518}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1508 ( .a ({signal_2843, signal_1385}), .b ({signal_2981, signal_1523}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1509 ( .a ({signal_2844, signal_1386}), .b ({signal_2982, signal_1524}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1510 ( .a ({signal_2845, signal_1387}), .b ({signal_2983, signal_1525}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1511 ( .a ({signal_2846, signal_1388}), .b ({signal_2984, signal_1526}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1512 ( .a ({signal_2847, signal_1389}), .b ({signal_2985, signal_1527}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1514 ( .a ({signal_2850, signal_1392}), .b ({signal_2987, signal_1529}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1515 ( .a ({signal_2851, signal_1393}), .b ({signal_2988, signal_1530}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1516 ( .a ({signal_2852, signal_1394}), .b ({signal_2989, signal_1531}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1517 ( .a ({signal_2853, signal_1395}), .b ({signal_2990, signal_1532}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1518 ( .a ({signal_2854, signal_1396}), .b ({signal_2991, signal_1533}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1519 ( .a ({signal_2855, signal_1397}), .b ({signal_2992, signal_1534}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1521 ( .a ({signal_2857, signal_1399}), .b ({signal_2994, signal_1536}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1522 ( .a ({signal_2858, signal_1400}), .b ({signal_2995, signal_1537}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1523 ( .a ({signal_2859, signal_1401}), .b ({signal_2996, signal_1538}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1524 ( .a ({signal_2860, signal_1402}), .b ({signal_2997, signal_1539}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1525 ( .a ({signal_2861, signal_1403}), .b ({signal_2998, signal_1540}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1526 ( .a ({signal_2862, signal_1404}), .b ({signal_2999, signal_1541}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1527 ( .a ({signal_2863, signal_1405}), .b ({signal_3000, signal_1542}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1528 ( .a ({signal_2864, signal_1406}), .b ({signal_3001, signal_1543}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1529 ( .a ({signal_2865, signal_1407}), .b ({signal_3002, signal_1544}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1530 ( .a ({signal_2866, signal_1408}), .b ({signal_3003, signal_1545}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1531 ( .a ({signal_2867, signal_1409}), .b ({signal_3004, signal_1546}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1534 ( .a ({signal_2870, signal_1412}), .b ({signal_3007, signal_1549}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1535 ( .a ({signal_2871, signal_1413}), .b ({signal_3008, signal_1550}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1536 ( .a ({signal_2872, signal_1414}), .b ({signal_3009, signal_1551}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1537 ( .a ({signal_2873, signal_1415}), .b ({signal_3010, signal_1552}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1540 ( .a ({signal_2877, signal_1419}), .b ({signal_3013, signal_1555}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1541 ( .a ({signal_2878, signal_1420}), .b ({signal_3014, signal_1556}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1542 ( .a ({signal_2879, signal_1421}), .b ({signal_3015, signal_1557}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1545 ( .a ({signal_2882, signal_1424}), .b ({signal_3018, signal_1560}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1546 ( .a ({signal_2883, signal_1425}), .b ({signal_3019, signal_1561}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1547 ( .a ({signal_2884, signal_1426}), .b ({signal_3020, signal_1562}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1548 ( .a ({signal_2885, signal_1427}), .b ({signal_3021, signal_1563}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1549 ( .a ({signal_2886, signal_1428}), .b ({signal_3022, signal_1564}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1550 ( .a ({signal_2887, signal_1429}), .b ({signal_3023, signal_1565}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1551 ( .a ({signal_2888, signal_1430}), .b ({signal_3024, signal_1566}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1552 ( .a ({signal_2889, signal_1431}), .b ({signal_3025, signal_1567}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1553 ( .a ({signal_2890, signal_1432}), .b ({signal_3026, signal_1568}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1554 ( .a ({signal_2891, signal_1433}), .b ({signal_3027, signal_1569}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1555 ( .a ({signal_2892, signal_1434}), .b ({signal_3028, signal_1570}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1556 ( .a ({signal_2893, signal_1435}), .b ({signal_3029, signal_1571}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1557 ( .a ({signal_2894, signal_1436}), .b ({signal_3030, signal_1572}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1558 ( .a ({signal_2895, signal_1437}), .b ({signal_3031, signal_1573}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1559 ( .a ({signal_2896, signal_1438}), .b ({signal_3032, signal_1574}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1560 ( .a ({signal_2897, signal_1439}), .b ({signal_3033, signal_1575}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1561 ( .a ({signal_2898, signal_1440}), .b ({signal_3034, signal_1576}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1562 ( .a ({signal_2899, signal_1441}), .b ({signal_3035, signal_1577}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1563 ( .a ({signal_2900, signal_1442}), .b ({signal_3036, signal_1578}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1564 ( .a ({signal_2901, signal_1443}), .b ({signal_3037, signal_1579}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1565 ( .a ({signal_2902, signal_1444}), .b ({signal_3038, signal_1580}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1566 ( .a ({signal_2903, signal_1445}), .b ({signal_3039, signal_1581}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1567 ( .a ({signal_2905, signal_1447}), .b ({signal_3040, signal_1582}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1568 ( .a ({signal_2906, signal_1448}), .b ({signal_3041, signal_1583}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1569 ( .a ({signal_2907, signal_1449}), .b ({signal_3042, signal_1584}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1570 ( .a ({signal_2908, signal_1450}), .b ({signal_3043, signal_1585}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1571 ( .a ({signal_2909, signal_1451}), .b ({signal_3044, signal_1586}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1572 ( .a ({signal_2910, signal_1452}), .b ({signal_3045, signal_1587}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1573 ( .a ({signal_2911, signal_1453}), .b ({signal_3046, signal_1588}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1574 ( .a ({signal_2912, signal_1454}), .b ({signal_3047, signal_1589}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1575 ( .a ({signal_2913, signal_1455}), .b ({signal_3048, signal_1590}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1576 ( .a ({signal_2914, signal_1456}), .b ({signal_3049, signal_1591}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1577 ( .a ({signal_2915, signal_1457}), .b ({signal_3050, signal_1592}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1578 ( .a ({signal_2916, signal_1458}), .b ({signal_3051, signal_1593}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1579 ( .a ({signal_2917, signal_1459}), .b ({signal_3052, signal_1594}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1580 ( .a ({signal_2918, signal_1460}), .b ({signal_3053, signal_1595}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1581 ( .a ({signal_2920, signal_1462}), .b ({signal_3054, signal_1596}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1582 ( .a ({signal_2921, signal_1463}), .b ({signal_3055, signal_1597}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1583 ( .a ({signal_2922, signal_1464}), .b ({signal_3056, signal_1598}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1584 ( .a ({signal_2923, signal_1465}), .b ({signal_3057, signal_1599}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1585 ( .a ({signal_2924, signal_1466}), .b ({signal_3058, signal_1600}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1586 ( .a ({signal_2925, signal_1467}), .b ({signal_3059, signal_1601}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1587 ( .a ({signal_2926, signal_1468}), .b ({signal_3060, signal_1602}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1588 ( .a ({signal_2927, signal_1469}), .b ({signal_3061, signal_1603}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1589 ( .a ({signal_2928, signal_1470}), .b ({signal_3062, signal_1604}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1590 ( .a ({signal_2929, signal_1471}), .b ({signal_3063, signal_1605}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1591 ( .a ({signal_2930, signal_1472}), .b ({signal_3064, signal_1606}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1592 ( .a ({signal_2931, signal_1473}), .b ({signal_3065, signal_1607}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1593 ( .a ({signal_2932, signal_1474}), .b ({signal_3066, signal_1608}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1594 ( .a ({signal_2933, signal_1475}), .b ({signal_3067, signal_1609}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1595 ( .a ({signal_2934, signal_1476}), .b ({signal_3068, signal_1610}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1596 ( .a ({signal_2935, signal_1477}), .b ({signal_3069, signal_1611}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1597 ( .a ({signal_2937, signal_1479}), .b ({signal_3070, signal_1612}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1598 ( .a ({signal_2938, signal_1480}), .b ({signal_3071, signal_1613}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1599 ( .a ({signal_2939, signal_1481}), .b ({signal_3072, signal_1614}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1600 ( .a ({signal_2940, signal_1482}), .b ({signal_3073, signal_1615}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1601 ( .a ({signal_2941, signal_1483}), .b ({signal_3074, signal_1616}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1602 ( .a ({signal_2942, signal_1484}), .b ({signal_3075, signal_1617}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1603 ( .a ({signal_2943, signal_1485}), .b ({signal_3076, signal_1618}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1604 ( .a ({signal_2944, signal_1486}), .b ({signal_3077, signal_1619}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1605 ( .a ({signal_2945, signal_1487}), .b ({signal_3078, signal_1620}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1606 ( .a ({signal_2946, signal_1488}), .b ({signal_3079, signal_1621}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1607 ( .a ({signal_2947, signal_1489}), .b ({signal_3080, signal_1622}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1608 ( .a ({signal_2948, signal_1490}), .b ({signal_3081, signal_1623}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1609 ( .a ({signal_2949, signal_1491}), .b ({signal_3082, signal_1624}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1610 ( .a ({signal_2950, signal_1492}), .b ({signal_3083, signal_1625}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1611 ( .a ({signal_2951, signal_1493}), .b ({signal_3084, signal_1626}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1612 ( .a ({signal_2952, signal_1494}), .b ({signal_3085, signal_1627}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1613 ( .a ({signal_2953, signal_1495}), .b ({signal_3086, signal_1628}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1614 ( .a ({signal_2954, signal_1496}), .b ({signal_3087, signal_1629}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1615 ( .a ({signal_2955, signal_1497}), .b ({signal_3088, signal_1630}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1616 ( .a ({signal_2956, signal_1498}), .b ({signal_3089, signal_1631}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1617 ( .a ({signal_2957, signal_1499}), .b ({signal_3090, signal_1632}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1618 ( .a ({signal_2958, signal_1500}), .b ({signal_3091, signal_1633}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1619 ( .a ({signal_2959, signal_1501}), .b ({signal_3092, signal_1634}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1620 ( .a ({signal_2960, signal_1502}), .b ({signal_3093, signal_1635}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1621 ( .a ({signal_2961, signal_1503}), .b ({signal_3094, signal_1636}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1622 ( .a ({signal_2962, signal_1504}), .b ({signal_3095, signal_1637}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1623 ( .a ({signal_2438, signal_980}), .b ({signal_2688, signal_1230}), .clk ( clk ), .r ( Fresh[368] ), .c ({signal_3096, signal_1638}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1624 ( .a ({signal_2515, signal_1057}), .b ({signal_2689, signal_1231}), .clk ( clk ), .r ( Fresh[369] ), .c ({signal_3097, signal_1639}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1625 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2694, signal_1236}), .clk ( clk ), .r ( Fresh[370] ), .c ({signal_3098, signal_1640}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1626 ( .a ({signal_2693, signal_1235}), .b ({signal_2714, signal_1256}), .clk ( clk ), .r ( Fresh[371] ), .c ({signal_3099, signal_1641}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1627 ( .a ({signal_2497, signal_1039}), .b ({signal_2715, signal_1257}), .clk ( clk ), .r ( Fresh[372] ), .c ({signal_3100, signal_1642}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1628 ( .a ({signal_2430, signal_972}), .b ({signal_2721, signal_1263}), .clk ( clk ), .r ( Fresh[373] ), .c ({signal_3101, signal_1643}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1629 ( .a ({signal_2708, signal_1250}), .b ({signal_2711, signal_1253}), .clk ( clk ), .r ( Fresh[374] ), .c ({signal_3102, signal_1644}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1630 ( .a ({signal_2725, signal_1267}), .b ({signal_2726, signal_1268}), .clk ( clk ), .r ( Fresh[375] ), .c ({signal_3103, signal_1645}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1631 ( .a ({signal_2504, signal_1046}), .b ({signal_2698, signal_1240}), .clk ( clk ), .r ( Fresh[376] ), .c ({signal_3104, signal_1646}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1632 ( .a ({signal_2727, signal_1269}), .b ({signal_2728, signal_1270}), .clk ( clk ), .r ( Fresh[377] ), .c ({signal_3105, signal_1647}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1633 ( .a ({signal_2693, signal_1235}), .b ({signal_2713, signal_1255}), .clk ( clk ), .r ( Fresh[378] ), .c ({signal_3106, signal_1648}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1634 ( .a ({signal_2731, signal_1273}), .b ({signal_2732, signal_1274}), .clk ( clk ), .r ( Fresh[379] ), .c ({signal_3107, signal_1649}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1635 ( .a ({signal_2513, signal_1055}), .b ({signal_2712, signal_1254}), .clk ( clk ), .r ( Fresh[380] ), .c ({signal_3108, signal_1650}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1636 ( .a ({signal_2434, signal_976}), .b ({signal_2699, signal_1241}), .clk ( clk ), .r ( Fresh[381] ), .c ({signal_3109, signal_1651}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1637 ( .a ({signal_2694, signal_1236}), .b ({signal_2517, signal_1059}), .clk ( clk ), .r ( Fresh[382] ), .c ({signal_3110, signal_1652}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1638 ( .a ({signal_2738, signal_1280}), .b ({signal_2739, signal_1281}), .clk ( clk ), .r ( Fresh[383] ), .c ({signal_3111, signal_1653}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1639 ( .a ({signal_2741, signal_1283}), .b ({signal_2742, signal_1284}), .clk ( clk ), .r ( Fresh[384] ), .c ({signal_3112, signal_1654}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1640 ( .a ({signal_2691, signal_1233}), .b ({signal_2744, signal_1286}), .clk ( clk ), .r ( Fresh[385] ), .c ({signal_3113, signal_1655}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1641 ( .a ({signal_2695, signal_1237}), .b ({signal_2746, signal_1288}), .clk ( clk ), .r ( Fresh[386] ), .c ({signal_3114, signal_1656}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1642 ( .a ({signal_2517, signal_1059}), .b ({signal_2696, signal_1238}), .clk ( clk ), .r ( Fresh[387] ), .c ({signal_3115, signal_1657}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1643 ( .a ({signal_2700, signal_1242}), .b ({signal_2701, signal_1243}), .clk ( clk ), .r ( Fresh[388] ), .c ({signal_3116, signal_1658}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1645 ( .a ({signal_2752, signal_1294}), .b ({signal_2753, signal_1295}), .clk ( clk ), .r ( Fresh[389] ), .c ({signal_3118, signal_1660}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1646 ( .a ({signal_2696, signal_1238}), .b ({signal_2760, signal_1302}), .clk ( clk ), .r ( Fresh[390] ), .c ({signal_3119, signal_1661}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1647 ( .a ({signal_2463, signal_1005}), .b ({signal_2764, signal_1306}), .clk ( clk ), .r ( Fresh[391] ), .c ({signal_3120, signal_1662}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1648 ( .a ({signal_2710, signal_1252}), .b ({signal_2768, signal_1310}), .clk ( clk ), .r ( Fresh[392] ), .c ({signal_3121, signal_1663}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1649 ( .a ({signal_2499, signal_1041}), .b ({signal_2841, signal_1383}), .clk ( clk ), .r ( Fresh[393] ), .c ({signal_3122, signal_1664}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1650 ( .a ({SI_s1[3], SI_s0[3]}), .b ({signal_2755, signal_1297}), .clk ( clk ), .r ( Fresh[394] ), .c ({signal_3123, signal_1665}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1651 ( .a ({signal_2702, signal_1244}), .b ({signal_2769, signal_1311}), .clk ( clk ), .r ( Fresh[395] ), .c ({signal_3124, signal_1666}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1653 ( .a ({signal_2834, signal_1376}), .b ({signal_2775, signal_1317}), .clk ( clk ), .r ( Fresh[396] ), .c ({signal_3126, signal_1668}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1654 ( .a ({signal_2693, signal_1235}), .b ({signal_2777, signal_1319}), .clk ( clk ), .r ( Fresh[397] ), .c ({signal_3127, signal_1669}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1655 ( .a ({signal_2848, signal_1390}), .b ({signal_2523, signal_1065}), .clk ( clk ), .r ( Fresh[398] ), .c ({signal_3128, signal_1670}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1656 ( .a ({signal_2456, signal_998}), .b ({signal_2778, signal_1320}), .clk ( clk ), .r ( Fresh[399] ), .c ({signal_3129, signal_1671}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1657 ( .a ({signal_2718, signal_1260}), .b ({signal_2758, signal_1300}), .clk ( clk ), .r ( Fresh[400] ), .c ({signal_3130, signal_1672}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1658 ( .a ({signal_2456, signal_998}), .b ({signal_2779, signal_1321}), .clk ( clk ), .r ( Fresh[401] ), .c ({signal_3131, signal_1673}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1659 ( .a ({signal_2774, signal_1316}), .b ({signal_2780, signal_1322}), .clk ( clk ), .r ( Fresh[402] ), .c ({signal_3132, signal_1674}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1660 ( .a ({signal_2521, signal_1063}), .b ({signal_2781, signal_1323}), .clk ( clk ), .r ( Fresh[403] ), .c ({signal_3133, signal_1675}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1661 ( .a ({signal_2782, signal_1324}), .b ({signal_2783, signal_1325}), .clk ( clk ), .r ( Fresh[404] ), .c ({signal_3134, signal_1676}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1663 ( .a ({signal_2698, signal_1240}), .b ({signal_2755, signal_1297}), .clk ( clk ), .r ( Fresh[405] ), .c ({signal_3136, signal_1678}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1664 ( .a ({signal_2722, signal_1264}), .b ({signal_2789, signal_1331}), .clk ( clk ), .r ( Fresh[406] ), .c ({signal_3137, signal_1679}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1665 ( .a ({signal_2700, signal_1242}), .b ({signal_2790, signal_1332}), .clk ( clk ), .r ( Fresh[407] ), .c ({signal_3138, signal_1680}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1666 ( .a ({signal_2724, signal_1266}), .b ({signal_2792, signal_1334}), .clk ( clk ), .r ( Fresh[408] ), .c ({signal_3139, signal_1681}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1667 ( .a ({signal_2755, signal_1297}), .b ({signal_2795, signal_1337}), .clk ( clk ), .r ( Fresh[409] ), .c ({signal_3140, signal_1682}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1668 ( .a ({signal_2729, signal_1271}), .b ({signal_2789, signal_1331}), .clk ( clk ), .r ( Fresh[410] ), .c ({signal_3141, signal_1683}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1669 ( .a ({signal_2437, signal_979}), .b ({signal_2778, signal_1320}), .clk ( clk ), .r ( Fresh[411] ), .c ({signal_3142, signal_1684}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1670 ( .a ({signal_2747, signal_1289}), .b ({signal_2798, signal_1340}), .clk ( clk ), .r ( Fresh[412] ), .c ({signal_3143, signal_1685}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1671 ( .a ({signal_2492, signal_1034}), .b ({signal_2799, signal_1341}), .clk ( clk ), .r ( Fresh[413] ), .c ({signal_3144, signal_1686}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1673 ( .a ({signal_2734, signal_1276}), .b ({signal_2788, signal_1330}), .clk ( clk ), .r ( Fresh[414] ), .c ({signal_3146, signal_1688}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1674 ( .a ({signal_2776, signal_1318}), .b ({signal_2876, signal_1418}), .clk ( clk ), .r ( Fresh[415] ), .c ({signal_3147, signal_1689}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1675 ( .a ({signal_2717, signal_1259}), .b ({signal_2782, signal_1324}), .clk ( clk ), .r ( Fresh[416] ), .c ({signal_3148, signal_1690}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1676 ( .a ({signal_2735, signal_1277}), .b ({signal_2804, signal_1346}), .clk ( clk ), .r ( Fresh[417] ), .c ({signal_3149, signal_1691}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1677 ( .a ({signal_2805, signal_1347}), .b ({signal_2806, signal_1348}), .clk ( clk ), .r ( Fresh[418] ), .c ({signal_3150, signal_1692}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1678 ( .a ({signal_2708, signal_1250}), .b ({signal_2807, signal_1349}), .clk ( clk ), .r ( Fresh[419] ), .c ({signal_3151, signal_1693}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1679 ( .a ({signal_2809, signal_1351}), .b ({signal_2810, signal_1352}), .clk ( clk ), .r ( Fresh[420] ), .c ({signal_3152, signal_1694}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1680 ( .a ({signal_2693, signal_1235}), .b ({signal_2767, signal_1309}), .clk ( clk ), .r ( Fresh[421] ), .c ({signal_3153, signal_1695}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1681 ( .a ({signal_2813, signal_1355}), .b ({signal_2814, signal_1356}), .clk ( clk ), .r ( Fresh[422] ), .c ({signal_3154, signal_1696}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1682 ( .a ({signal_2773, signal_1315}), .b ({signal_2815, signal_1357}), .clk ( clk ), .r ( Fresh[423] ), .c ({signal_3155, signal_1697}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1684 ( .a ({signal_2747, signal_1289}), .b ({signal_2748, signal_1290}), .clk ( clk ), .r ( Fresh[424] ), .c ({signal_3157, signal_1699}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1687 ( .a ({signal_2701, signal_1243}), .b ({signal_2748, signal_1290}), .clk ( clk ), .r ( Fresh[425] ), .c ({signal_3160, signal_1702}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1693 ( .a ({signal_2748, signal_1290}), .b ({signal_2763, signal_1305}), .clk ( clk ), .r ( Fresh[426] ), .c ({signal_3166, signal_1708}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1698 ( .a ({signal_2751, signal_1293}), .b ({signal_2822, signal_1364}), .clk ( clk ), .r ( Fresh[427] ), .c ({signal_3171, signal_1713}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1700 ( .a ({signal_3096, signal_1638}), .b ({signal_3173, signal_1715}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1701 ( .a ({signal_3097, signal_1639}), .b ({signal_3174, signal_1716}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1702 ( .a ({signal_3099, signal_1641}), .b ({signal_3175, signal_1717}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1703 ( .a ({signal_3100, signal_1642}), .b ({signal_3176, signal_1718}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1704 ( .a ({signal_3101, signal_1643}), .b ({signal_3177, signal_1719}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1705 ( .a ({signal_3102, signal_1644}), .b ({signal_3178, signal_1720}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1706 ( .a ({signal_3104, signal_1646}), .b ({signal_3179, signal_1721}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1707 ( .a ({signal_3105, signal_1647}), .b ({signal_3180, signal_1722}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1708 ( .a ({signal_3106, signal_1648}), .b ({signal_3181, signal_1723}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1709 ( .a ({signal_3108, signal_1650}), .b ({signal_3182, signal_1724}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1710 ( .a ({signal_3109, signal_1651}), .b ({signal_3183, signal_1725}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1711 ( .a ({signal_3110, signal_1652}), .b ({signal_3184, signal_1726}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1712 ( .a ({signal_3114, signal_1656}), .b ({signal_3185, signal_1727}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1713 ( .a ({signal_3115, signal_1657}), .b ({signal_3186, signal_1728}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1714 ( .a ({signal_3116, signal_1658}), .b ({signal_3187, signal_1729}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1716 ( .a ({signal_3120, signal_1662}), .b ({signal_3189, signal_1731}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1717 ( .a ({signal_3121, signal_1663}), .b ({signal_3190, signal_1732}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1718 ( .a ({signal_3122, signal_1664}), .b ({signal_3191, signal_1733}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1719 ( .a ({signal_3123, signal_1665}), .b ({signal_3192, signal_1734}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1720 ( .a ({signal_3124, signal_1666}), .b ({signal_3193, signal_1735}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1722 ( .a ({signal_3127, signal_1669}), .b ({signal_3195, signal_1737}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1723 ( .a ({signal_3131, signal_1673}), .b ({signal_3196, signal_1738}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1724 ( .a ({signal_3134, signal_1676}), .b ({signal_3197, signal_1739}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1726 ( .a ({signal_3136, signal_1678}), .b ({signal_3199, signal_1741}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1727 ( .a ({signal_3137, signal_1679}), .b ({signal_3200, signal_1742}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1728 ( .a ({signal_3138, signal_1680}), .b ({signal_3201, signal_1743}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1729 ( .a ({signal_3139, signal_1681}), .b ({signal_3202, signal_1744}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1730 ( .a ({signal_3140, signal_1682}), .b ({signal_3203, signal_1745}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1731 ( .a ({signal_3144, signal_1686}), .b ({signal_3204, signal_1746}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1732 ( .a ({signal_3147, signal_1689}), .b ({signal_3205, signal_1747}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1733 ( .a ({signal_3151, signal_1693}), .b ({signal_3206, signal_1748}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1734 ( .a ({signal_3154, signal_1696}), .b ({signal_3207, signal_1749}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1735 ( .a ({signal_3155, signal_1697}), .b ({signal_3208, signal_1750}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1736 ( .a ({signal_3157, signal_1699}), .b ({signal_3209, signal_1751}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1739 ( .a ({signal_3160, signal_1702}), .b ({signal_3212, signal_1754}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1745 ( .a ({signal_3166, signal_1708}), .b ({signal_3218, signal_1760}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1749 ( .a ({signal_3171, signal_1713}), .b ({signal_3222, signal_1764}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1751 ( .a ({signal_2560, signal_1102}), .b ({signal_2965, signal_1507}), .clk ( clk ), .r ( Fresh[428] ), .c ({signal_3224, signal_1766}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1753 ( .a ({signal_2395, signal_943}), .b ({signal_2966, signal_1508}), .clk ( clk ), .r ( Fresh[429] ), .c ({signal_3226, signal_1768}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1754 ( .a ({SI_s1[4], SI_s0[4]}), .b ({signal_2967, signal_1509}), .clk ( clk ), .r ( Fresh[430] ), .c ({signal_3227, signal_1769}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1755 ( .a ({signal_2541, signal_1083}), .b ({signal_2968, signal_1510}), .clk ( clk ), .r ( Fresh[431] ), .c ({signal_3228, signal_1770}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1756 ( .a ({signal_2415, signal_957}), .b ({signal_2965, signal_1507}), .clk ( clk ), .r ( Fresh[432] ), .c ({signal_3229, signal_1771}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1757 ( .a ({signal_2590, signal_1132}), .b ({signal_2969, signal_1511}), .clk ( clk ), .r ( Fresh[433] ), .c ({signal_3230, signal_1772}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1758 ( .a ({signal_2457, signal_999}), .b ({signal_2969, signal_1511}), .clk ( clk ), .r ( Fresh[434] ), .c ({signal_3231, signal_1773}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1760 ( .a ({signal_2454, signal_996}), .b ({signal_2972, signal_1514}), .clk ( clk ), .r ( Fresh[435] ), .c ({signal_3233, signal_1775}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1761 ( .a ({signal_2452, signal_994}), .b ({signal_2973, signal_1515}), .clk ( clk ), .r ( Fresh[436] ), .c ({signal_3234, signal_1776}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1762 ( .a ({signal_2450, signal_992}), .b ({signal_2974, signal_1516}), .clk ( clk ), .r ( Fresh[437] ), .c ({signal_3235, signal_1777}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1764 ( .a ({signal_2467, signal_1009}), .b ({signal_2977, signal_1519}), .clk ( clk ), .r ( Fresh[438] ), .c ({signal_3237, signal_1779}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1765 ( .a ({signal_2463, signal_1005}), .b ({signal_2978, signal_1520}), .clk ( clk ), .r ( Fresh[439] ), .c ({signal_3238, signal_1780}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1766 ( .a ({signal_2449, signal_991}), .b ({signal_2979, signal_1521}), .clk ( clk ), .r ( Fresh[440] ), .c ({signal_3239, signal_1781}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1767 ( .a ({signal_2407, signal_949}), .b ({signal_2980, signal_1522}), .clk ( clk ), .r ( Fresh[441] ), .c ({signal_3240, signal_1782}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1769 ( .a ({signal_2536, signal_1078}), .b ({signal_2980, signal_1522}), .clk ( clk ), .r ( Fresh[442] ), .c ({signal_3242, signal_1784}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1770 ( .a ({signal_2543, signal_1085}), .b ({signal_2986, signal_1528}), .clk ( clk ), .r ( Fresh[443] ), .c ({signal_3243, signal_1785}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1772 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2979, signal_1521}), .clk ( clk ), .r ( Fresh[444] ), .c ({signal_3245, signal_1787}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1773 ( .a ({signal_2611, signal_1153}), .b ({signal_2993, signal_1535}), .clk ( clk ), .r ( Fresh[445] ), .c ({signal_3246, signal_1788}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1776 ( .a ({signal_2439, signal_981}), .b ({signal_2978, signal_1520}), .clk ( clk ), .r ( Fresh[446] ), .c ({signal_3249, signal_1791}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1778 ( .a ({signal_2443, signal_985}), .b ({signal_3005, signal_1547}), .clk ( clk ), .r ( Fresh[447] ), .c ({signal_3251, signal_1793}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1779 ( .a ({signal_2544, signal_1086}), .b ({signal_3006, signal_1548}), .clk ( clk ), .r ( Fresh[448] ), .c ({signal_3252, signal_1794}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1782 ( .a ({signal_2456, signal_998}), .b ({signal_3011, signal_1553}), .clk ( clk ), .r ( Fresh[449] ), .c ({signal_3255, signal_1797}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1783 ( .a ({signal_2466, signal_1008}), .b ({signal_3012, signal_1554}), .clk ( clk ), .r ( Fresh[450] ), .c ({signal_3256, signal_1798}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1784 ( .a ({signal_2540, signal_1082}), .b ({signal_2973, signal_1515}), .clk ( clk ), .r ( Fresh[451] ), .c ({signal_3257, signal_1799}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1785 ( .a ({signal_2465, signal_1007}), .b ({signal_3016, signal_1558}), .clk ( clk ), .r ( Fresh[452] ), .c ({signal_3258, signal_1800}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1786 ( .a ({signal_2456, signal_998}), .b ({signal_3017, signal_1559}), .clk ( clk ), .r ( Fresh[453] ), .c ({signal_3259, signal_1801}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1835 ( .a ({signal_3224, signal_1766}), .b ({signal_3308, signal_1850}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1836 ( .a ({signal_3228, signal_1770}), .b ({signal_3309, signal_1851}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1837 ( .a ({signal_3230, signal_1772}), .b ({signal_3310, signal_1852}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1838 ( .a ({signal_3231, signal_1773}), .b ({signal_3311, signal_1853}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1839 ( .a ({signal_3233, signal_1775}), .b ({signal_3312, signal_1854}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1840 ( .a ({signal_3234, signal_1776}), .b ({signal_3313, signal_1855}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1841 ( .a ({signal_3235, signal_1777}), .b ({signal_3314, signal_1856}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1843 ( .a ({signal_3237, signal_1779}), .b ({signal_3316, signal_1858}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1844 ( .a ({signal_3238, signal_1780}), .b ({signal_3317, signal_1859}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1845 ( .a ({signal_3239, signal_1781}), .b ({signal_3318, signal_1860}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1846 ( .a ({signal_3242, signal_1784}), .b ({signal_3319, signal_1861}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1847 ( .a ({signal_3243, signal_1785}), .b ({signal_3320, signal_1862}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1848 ( .a ({signal_3245, signal_1787}), .b ({signal_3321, signal_1863}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1849 ( .a ({signal_3246, signal_1788}), .b ({signal_3322, signal_1864}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1850 ( .a ({signal_3249, signal_1791}), .b ({signal_3323, signal_1865}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1851 ( .a ({signal_3251, signal_1793}), .b ({signal_3324, signal_1866}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1852 ( .a ({signal_3252, signal_1794}), .b ({signal_3325, signal_1867}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1854 ( .a ({signal_3255, signal_1797}), .b ({signal_3327, signal_1869}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1855 ( .a ({signal_3256, signal_1798}), .b ({signal_3328, signal_1870}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1856 ( .a ({signal_3257, signal_1799}), .b ({signal_3329, signal_1871}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1857 ( .a ({signal_3258, signal_1800}), .b ({signal_3330, signal_1872}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1858 ( .a ({signal_3259, signal_1801}), .b ({signal_3331, signal_1873}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1644 ( .a ({signal_2750, signal_1292}), .b ({signal_2751, signal_1293}), .clk ( clk ), .r ( Fresh[454] ), .c ({signal_3117, signal_1659}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1652 ( .a ({signal_2462, signal_1004}), .b ({signal_2843, signal_1385}), .clk ( clk ), .r ( Fresh[455] ), .c ({signal_3125, signal_1667}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1662 ( .a ({signal_2786, signal_1328}), .b ({signal_2787, signal_1329}), .clk ( clk ), .r ( Fresh[456] ), .c ({signal_3135, signal_1677}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1672 ( .a ({signal_2800, signal_1342}), .b ({signal_2801, signal_1343}), .clk ( clk ), .r ( Fresh[457] ), .c ({signal_3145, signal_1687}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1683 ( .a ({signal_2740, signal_1282}), .b ({signal_2816, signal_1358}), .clk ( clk ), .r ( Fresh[458] ), .c ({signal_3156, signal_1698}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1685 ( .a ({signal_2749, signal_1291}), .b ({signal_2818, signal_1360}), .clk ( clk ), .r ( Fresh[459] ), .c ({signal_3158, signal_1700}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1686 ( .a ({signal_2417, signal_959}), .b ({signal_2904, signal_1446}), .clk ( clk ), .r ( Fresh[460] ), .c ({signal_3159, signal_1701}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1688 ( .a ({signal_2458, signal_1000}), .b ({signal_2904, signal_1446}), .clk ( clk ), .r ( Fresh[461] ), .c ({signal_3161, signal_1703}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1689 ( .a ({signal_2458, signal_1000}), .b ({signal_2918, signal_1460}), .clk ( clk ), .r ( Fresh[462] ), .c ({signal_3162, signal_1704}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1690 ( .a ({signal_2407, signal_949}), .b ({signal_2919, signal_1461}), .clk ( clk ), .r ( Fresh[463] ), .c ({signal_3163, signal_1705}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1691 ( .a ({signal_2434, signal_976}), .b ({signal_2920, signal_1462}), .clk ( clk ), .r ( Fresh[464] ), .c ({signal_3164, signal_1706}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1692 ( .a ({signal_2420, signal_962}), .b ({signal_2908, signal_1450}), .clk ( clk ), .r ( Fresh[465] ), .c ({signal_3165, signal_1707}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1694 ( .a ({SI_s1[7], SI_s0[7]}), .b ({signal_2936, signal_1478}), .clk ( clk ), .r ( Fresh[466] ), .c ({signal_3167, signal_1709}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1695 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_2821, signal_1363}), .clk ( clk ), .r ( Fresh[467] ), .c ({signal_3168, signal_1710}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1696 ( .a ({signal_2504, signal_1046}), .b ({signal_2893, signal_1435}), .clk ( clk ), .r ( Fresh[468] ), .c ({signal_3169, signal_1711}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1697 ( .a ({signal_2450, signal_992}), .b ({signal_2932, signal_1474}), .clk ( clk ), .r ( Fresh[469] ), .c ({signal_3170, signal_1712}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1699 ( .a ({signal_2408, signal_950}), .b ({signal_2955, signal_1497}), .clk ( clk ), .r ( Fresh[470] ), .c ({signal_3172, signal_1714}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1715 ( .a ({signal_3117, signal_1659}), .b ({signal_3188, signal_1730}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1721 ( .a ({signal_3125, signal_1667}), .b ({signal_3194, signal_1736}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1725 ( .a ({signal_3135, signal_1677}), .b ({signal_3198, signal_1740}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1737 ( .a ({signal_3158, signal_1700}), .b ({signal_3210, signal_1752}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1738 ( .a ({signal_3159, signal_1701}), .b ({signal_3211, signal_1753}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1740 ( .a ({signal_3161, signal_1703}), .b ({signal_3213, signal_1755}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1741 ( .a ({signal_3162, signal_1704}), .b ({signal_3214, signal_1756}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1742 ( .a ({signal_3163, signal_1705}), .b ({signal_3215, signal_1757}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1743 ( .a ({signal_3164, signal_1706}), .b ({signal_3216, signal_1758}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1744 ( .a ({signal_3165, signal_1707}), .b ({signal_3217, signal_1759}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1746 ( .a ({signal_3167, signal_1709}), .b ({signal_3219, signal_1761}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1747 ( .a ({signal_3169, signal_1711}), .b ({signal_3220, signal_1762}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1748 ( .a ({signal_3170, signal_1712}), .b ({signal_3221, signal_1763}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1750 ( .a ({signal_3172, signal_1714}), .b ({signal_3223, signal_1765}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1752 ( .a ({signal_2989, signal_1531}), .b ({signal_2990, signal_1532}), .clk ( clk ), .r ( Fresh[471] ), .c ({signal_3225, signal_1767}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1759 ( .a ({signal_2506, signal_1048}), .b ({signal_2970, signal_1512}), .clk ( clk ), .r ( Fresh[472] ), .c ({signal_3232, signal_1774}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1763 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_2975, signal_1517}), .clk ( clk ), .r ( Fresh[473] ), .c ({signal_3236, signal_1778}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1768 ( .a ({signal_2983, signal_1525}), .b ({signal_2984, signal_1526}), .clk ( clk ), .r ( Fresh[474] ), .c ({signal_3241, signal_1783}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1771 ( .a ({signal_2981, signal_1523}), .b ({signal_2988, signal_1530}), .clk ( clk ), .r ( Fresh[475] ), .c ({signal_3244, signal_1786}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1774 ( .a ({signal_2720, signal_1262}), .b ({signal_2994, signal_1536}), .clk ( clk ), .r ( Fresh[476] ), .c ({signal_3247, signal_1789}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1775 ( .a ({signal_2999, signal_1541}), .b ({signal_3000, signal_1542}), .clk ( clk ), .r ( Fresh[477] ), .c ({signal_3248, signal_1790}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1777 ( .a ({signal_2702, signal_1244}), .b ({signal_3004, signal_1546}), .clk ( clk ), .r ( Fresh[478] ), .c ({signal_3250, signal_1792}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1780 ( .a ({signal_2733, signal_1275}), .b ({signal_3107, signal_1649}), .clk ( clk ), .r ( Fresh[479] ), .c ({signal_3253, signal_1795}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1781 ( .a ({signal_3052, signal_1594}), .b ({signal_3069, signal_1611}), .clk ( clk ), .r ( Fresh[480] ), .c ({signal_3254, signal_1796}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1787 ( .a ({signal_2713, signal_1255}), .b ({signal_3019, signal_1561}), .clk ( clk ), .r ( Fresh[481] ), .c ({signal_3260, signal_1802}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1788 ( .a ({signal_3021, signal_1563}), .b ({signal_2811, signal_1353}), .clk ( clk ), .r ( Fresh[482] ), .c ({signal_3261, signal_1803}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1789 ( .a ({signal_2807, signal_1349}), .b ({signal_3111, signal_1653}), .clk ( clk ), .r ( Fresh[483] ), .c ({signal_3262, signal_1804}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1790 ( .a ({signal_2690, signal_1232}), .b ({signal_3112, signal_1654}), .clk ( clk ), .r ( Fresh[484] ), .c ({signal_3263, signal_1805}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1791 ( .a ({signal_2743, signal_1285}), .b ({signal_3113, signal_1655}), .clk ( clk ), .r ( Fresh[485] ), .c ({signal_3264, signal_1806}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1792 ( .a ({signal_3024, signal_1566}), .b ({signal_3025, signal_1567}), .clk ( clk ), .r ( Fresh[486] ), .c ({signal_3265, signal_1807}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1793 ( .a ({signal_2745, signal_1287}), .b ({signal_3026, signal_1568}), .clk ( clk ), .r ( Fresh[487] ), .c ({signal_3266, signal_1808}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1794 ( .a ({signal_3098, signal_1640}), .b ({signal_3027, signal_1569}), .clk ( clk ), .r ( Fresh[488] ), .c ({signal_3267, signal_1809}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1795 ( .a ({signal_2407, signal_949}), .b ({signal_3029, signal_1571}), .clk ( clk ), .r ( Fresh[489] ), .c ({signal_3268, signal_1810}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1796 ( .a ({signal_2971, signal_1513}), .b ({signal_3030, signal_1572}), .clk ( clk ), .r ( Fresh[490] ), .c ({signal_3269, signal_1811}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1797 ( .a ({signal_2703, signal_1245}), .b ({signal_3031, signal_1573}), .clk ( clk ), .r ( Fresh[491] ), .c ({signal_3270, signal_1812}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1798 ( .a ({signal_2704, signal_1246}), .b ({signal_3118, signal_1660}), .clk ( clk ), .r ( Fresh[492] ), .c ({signal_3271, signal_1813}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1799 ( .a ({signal_2521, signal_1063}), .b ({signal_3032, signal_1574}), .clk ( clk ), .r ( Fresh[493] ), .c ({signal_3272, signal_1814}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1800 ( .a ({signal_2759, signal_1301}), .b ({signal_3035, signal_1577}), .clk ( clk ), .r ( Fresh[494] ), .c ({signal_3273, signal_1815}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1801 ( .a ({signal_2707, signal_1249}), .b ({signal_3119, signal_1661}), .clk ( clk ), .r ( Fresh[495] ), .c ({signal_3274, signal_1816}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1802 ( .a ({signal_2761, signal_1303}), .b ({signal_3024, signal_1566}), .clk ( clk ), .r ( Fresh[496] ), .c ({signal_3275, signal_1817}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1803 ( .a ({signal_3037, signal_1579}), .b ({signal_3038, signal_1580}), .clk ( clk ), .r ( Fresh[497] ), .c ({signal_3276, signal_1818}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1804 ( .a ({signal_2982, signal_1524}), .b ({signal_3043, signal_1585}), .clk ( clk ), .r ( Fresh[498] ), .c ({signal_3277, signal_1819}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1805 ( .a ({signal_3032, signal_1574}), .b ({signal_3044, signal_1586}), .clk ( clk ), .r ( Fresh[499] ), .c ({signal_3278, signal_1820}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1806 ( .a ({signal_2512, signal_1054}), .b ({signal_3126, signal_1668}), .clk ( clk ), .r ( Fresh[500] ), .c ({signal_3279, signal_1821}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1807 ( .a ({signal_2711, signal_1253}), .b ({signal_3124, signal_1666}), .clk ( clk ), .r ( Fresh[501] ), .c ({signal_3280, signal_1822}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1808 ( .a ({signal_2717, signal_1259}), .b ({signal_3128, signal_1670}), .clk ( clk ), .r ( Fresh[502] ), .c ({signal_3281, signal_1823}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1809 ( .a ({signal_2410, signal_952}), .b ({signal_3129, signal_1671}), .clk ( clk ), .r ( Fresh[503] ), .c ({signal_3282, signal_1824}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1810 ( .a ({signal_3087, signal_1629}), .b ({signal_3088, signal_1630}), .clk ( clk ), .r ( Fresh[504] ), .c ({signal_3283, signal_1825}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1811 ( .a ({signal_2987, signal_1529}), .b ({signal_3130, signal_1672}), .clk ( clk ), .r ( Fresh[505] ), .c ({signal_3284, signal_1826}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1812 ( .a ({signal_2996, signal_1538}), .b ({signal_3057, signal_1599}), .clk ( clk ), .r ( Fresh[506] ), .c ({signal_3285, signal_1827}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1813 ( .a ({signal_3002, signal_1544}), .b ({signal_3063, signal_1605}), .clk ( clk ), .r ( Fresh[507] ), .c ({signal_3286, signal_1828}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1814 ( .a ({signal_3003, signal_1545}), .b ({signal_3065, signal_1607}), .clk ( clk ), .r ( Fresh[508] ), .c ({signal_3287, signal_1829}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1815 ( .a ({signal_2797, signal_1339}), .b ({signal_3066, signal_1608}), .clk ( clk ), .r ( Fresh[509] ), .c ({signal_3288, signal_1830}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1816 ( .a ({signal_2405, signal_948}), .b ({signal_3142, signal_1684}), .clk ( clk ), .r ( Fresh[510] ), .c ({signal_3289, signal_1831}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1817 ( .a ({signal_2730, signal_1272}), .b ({signal_3143, signal_1685}), .clk ( clk ), .r ( Fresh[511] ), .c ({signal_3290, signal_1832}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1818 ( .a ({signal_3029, signal_1571}), .b ({signal_3054, signal_1596}), .clk ( clk ), .r ( Fresh[512] ), .c ({signal_3291, signal_1833}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1820 ( .a ({signal_2802, signal_1344}), .b ({signal_3068, signal_1610}), .clk ( clk ), .r ( Fresh[513] ), .c ({signal_3293, signal_1835}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1821 ( .a ({signal_2520, signal_1062}), .b ({signal_3070, signal_1612}), .clk ( clk ), .r ( Fresh[514] ), .c ({signal_3294, signal_1836}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1822 ( .a ({signal_2803, signal_1345}), .b ({signal_3073, signal_1615}), .clk ( clk ), .r ( Fresh[515] ), .c ({signal_3295, signal_1837}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1823 ( .a ({signal_3014, signal_1556}), .b ({signal_3075, signal_1617}), .clk ( clk ), .r ( Fresh[516] ), .c ({signal_3296, signal_1838}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1824 ( .a ({signal_2736, signal_1278}), .b ({signal_3150, signal_1692}), .clk ( clk ), .r ( Fresh[517] ), .c ({signal_3297, signal_1839}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1825 ( .a ({signal_2696, signal_1238}), .b ({signal_3078, signal_1620}), .clk ( clk ), .r ( Fresh[518] ), .c ({signal_3298, signal_1840}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1826 ( .a ({signal_2737, signal_1279}), .b ({signal_3073, signal_1615}), .clk ( clk ), .r ( Fresh[519] ), .c ({signal_3299, signal_1841}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1827 ( .a ({signal_2691, signal_1233}), .b ({signal_3153, signal_1695}), .clk ( clk ), .r ( Fresh[520] ), .c ({signal_3300, signal_1842}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1828 ( .a ({signal_3022, signal_1564}), .b ({signal_3081, signal_1623}), .clk ( clk ), .r ( Fresh[521] ), .c ({signal_3301, signal_1843}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1829 ( .a ({signal_2744, signal_1286}), .b ({signal_3082, signal_1624}), .clk ( clk ), .r ( Fresh[522] ), .c ({signal_3302, signal_1844}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1830 ( .a ({signal_3084, signal_1626}), .b ({signal_3085, signal_1627}), .clk ( clk ), .r ( Fresh[523] ), .c ({signal_3303, signal_1845}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1831 ( .a ({signal_3050, signal_1592}), .b ({signal_3086, signal_1628}), .clk ( clk ), .r ( Fresh[524] ), .c ({signal_3304, signal_1846}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1832 ( .a ({signal_2981, signal_1523}), .b ({signal_3092, signal_1634}), .clk ( clk ), .r ( Fresh[525] ), .c ({signal_3305, signal_1847}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1833 ( .a ({signal_2820, signal_1362}), .b ({signal_3093, signal_1635}), .clk ( clk ), .r ( Fresh[526] ), .c ({signal_3306, signal_1848}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1842 ( .a ({signal_3236, signal_1778}), .b ({signal_3315, signal_1857}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1853 ( .a ({signal_3253, signal_1795}), .b ({signal_3326, signal_1868}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1859 ( .a ({signal_3263, signal_1805}), .b ({signal_3332, signal_1874}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1860 ( .a ({signal_3265, signal_1807}), .b ({signal_3333, signal_1875}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1861 ( .a ({signal_3270, signal_1812}), .b ({signal_3334, signal_1876}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1862 ( .a ({signal_3274, signal_1816}), .b ({signal_3335, signal_1877}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1863 ( .a ({signal_3275, signal_1817}), .b ({signal_3336, signal_1878}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1864 ( .a ({signal_3279, signal_1821}), .b ({signal_3337, signal_1879}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1865 ( .a ({signal_3280, signal_1822}), .b ({signal_3338, signal_1880}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1866 ( .a ({signal_3281, signal_1823}), .b ({signal_3339, signal_1881}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1867 ( .a ({signal_3282, signal_1824}), .b ({signal_3340, signal_1882}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1868 ( .a ({signal_3286, signal_1828}), .b ({signal_3341, signal_1883}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1869 ( .a ({signal_3287, signal_1829}), .b ({signal_3342, signal_1884}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1870 ( .a ({signal_3289, signal_1831}), .b ({signal_3343, signal_1885}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1871 ( .a ({signal_3290, signal_1832}), .b ({signal_3344, signal_1886}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1873 ( .a ({signal_3300, signal_1842}), .b ({signal_3346, signal_1888}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1874 ( .a ({signal_3302, signal_1844}), .b ({signal_3347, signal_1889}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1876 ( .a ({signal_3173, signal_1715}), .b ({signal_2723, signal_1265}), .clk ( clk ), .r ( Fresh[527] ), .c ({signal_3349, signal_1891}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1877 ( .a ({signal_2416, signal_958}), .b ({signal_3174, signal_1716}), .clk ( clk ), .r ( Fresh[528] ), .c ({signal_3350, signal_1892}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1878 ( .a ({signal_2446, signal_988}), .b ({signal_3175, signal_1717}), .clk ( clk ), .r ( Fresh[529] ), .c ({signal_3351, signal_1893}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1879 ( .a ({signal_2458, signal_1000}), .b ({signal_3176, signal_1718}), .clk ( clk ), .r ( Fresh[530] ), .c ({signal_3352, signal_1894}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1880 ( .a ({signal_2408, signal_950}), .b ({signal_3226, signal_1768}), .clk ( clk ), .r ( Fresh[531] ), .c ({signal_3353, signal_1895}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1881 ( .a ({signal_2412, signal_954}), .b ({signal_3177, signal_1719}), .clk ( clk ), .r ( Fresh[532] ), .c ({signal_3354, signal_1896}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1882 ( .a ({signal_3178, signal_1720}), .b ({signal_2791, signal_1333}), .clk ( clk ), .r ( Fresh[533] ), .c ({signal_3355, signal_1897}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1883 ( .a ({signal_2465, signal_1007}), .b ({signal_3179, signal_1721}), .clk ( clk ), .r ( Fresh[534] ), .c ({signal_3356, signal_1898}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1884 ( .a ({signal_2395, signal_943}), .b ({signal_3180, signal_1722}), .clk ( clk ), .r ( Fresh[535] ), .c ({signal_3357, signal_1899}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1885 ( .a ({signal_2403, signal_947}), .b ({signal_3181, signal_1723}), .clk ( clk ), .r ( Fresh[536] ), .c ({signal_3358, signal_1900}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1886 ( .a ({signal_2420, signal_962}), .b ({signal_3227, signal_1769}), .clk ( clk ), .r ( Fresh[537] ), .c ({signal_3359, signal_1901}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1887 ( .a ({signal_2456, signal_998}), .b ({signal_3182, signal_1724}), .clk ( clk ), .r ( Fresh[538] ), .c ({signal_3360, signal_1902}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1888 ( .a ({signal_2466, signal_1008}), .b ({signal_3184, signal_1726}), .clk ( clk ), .r ( Fresh[539] ), .c ({signal_3361, signal_1903}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1889 ( .a ({signal_2409, signal_951}), .b ({signal_3229, signal_1771}), .clk ( clk ), .r ( Fresh[540] ), .c ({signal_3362, signal_1904}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1890 ( .a ({signal_2458, signal_1000}), .b ({signal_3185, signal_1727}), .clk ( clk ), .r ( Fresh[541] ), .c ({signal_3363, signal_1905}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1891 ( .a ({signal_2408, signal_950}), .b ({signal_3186, signal_1728}), .clk ( clk ), .r ( Fresh[542] ), .c ({signal_3364, signal_1906}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1892 ( .a ({signal_2603, signal_1145}), .b ({signal_3187, signal_1729}), .clk ( clk ), .r ( Fresh[543] ), .c ({signal_3365, signal_1907}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1894 ( .a ({SI_s1[1], SI_s0[1]}), .b ({signal_3189, signal_1731}), .clk ( clk ), .r ( Fresh[544] ), .c ({signal_3367, signal_1909}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1895 ( .a ({signal_2421, signal_963}), .b ({signal_3190, signal_1732}), .clk ( clk ), .r ( Fresh[545] ), .c ({signal_3368, signal_1910}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1896 ( .a ({signal_2553, signal_1095}), .b ({signal_3191, signal_1733}), .clk ( clk ), .r ( Fresh[546] ), .c ({signal_3369, signal_1911}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1897 ( .a ({signal_2536, signal_1078}), .b ({signal_3192, signal_1734}), .clk ( clk ), .r ( Fresh[547] ), .c ({signal_3370, signal_1912}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1898 ( .a ({signal_2531, signal_1073}), .b ({signal_3240, signal_1782}), .clk ( clk ), .r ( Fresh[548] ), .c ({signal_3371, signal_1913}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1899 ( .a ({signal_2616, signal_1158}), .b ({signal_3193, signal_1735}), .clk ( clk ), .r ( Fresh[549] ), .c ({signal_3372, signal_1914}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1900 ( .a ({signal_2466, signal_1008}), .b ({signal_3195, signal_1737}), .clk ( clk ), .r ( Fresh[550] ), .c ({signal_3373, signal_1915}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1901 ( .a ({signal_3196, signal_1738}), .b ({signal_3132, signal_1674}), .clk ( clk ), .r ( Fresh[551] ), .c ({signal_3374, signal_1916}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1903 ( .a ({signal_2407, signal_949}), .b ({signal_3197, signal_1739}), .clk ( clk ), .r ( Fresh[552] ), .c ({signal_3376, signal_1918}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1905 ( .a ({signal_2553, signal_1095}), .b ({signal_3199, signal_1741}), .clk ( clk ), .r ( Fresh[553] ), .c ({signal_3378, signal_1920}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1906 ( .a ({signal_2450, signal_992}), .b ({signal_3200, signal_1742}), .clk ( clk ), .r ( Fresh[554] ), .c ({signal_3379, signal_1921}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1907 ( .a ({signal_2405, signal_948}), .b ({signal_3201, signal_1743}), .clk ( clk ), .r ( Fresh[555] ), .c ({signal_3380, signal_1922}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1908 ( .a ({signal_2412, signal_954}), .b ({signal_3202, signal_1744}), .clk ( clk ), .r ( Fresh[556] ), .c ({signal_3381, signal_1923}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1909 ( .a ({signal_2478, signal_1020}), .b ({signal_3240, signal_1782}), .clk ( clk ), .r ( Fresh[557] ), .c ({signal_3382, signal_1924}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1910 ( .a ({signal_2463, signal_1005}), .b ({signal_3203, signal_1745}), .clk ( clk ), .r ( Fresh[558] ), .c ({signal_3383, signal_1925}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1913 ( .a ({signal_2415, signal_957}), .b ({signal_3204, signal_1746}), .clk ( clk ), .r ( Fresh[559] ), .c ({signal_3386, signal_1928}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1914 ( .a ({signal_2450, signal_992}), .b ({signal_3205, signal_1747}), .clk ( clk ), .r ( Fresh[560] ), .c ({signal_3387, signal_1929}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1915 ( .a ({signal_2458, signal_1000}), .b ({signal_3206, signal_1748}), .clk ( clk ), .r ( Fresh[561] ), .c ({signal_3388, signal_1930}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1916 ( .a ({signal_2620, signal_1162}), .b ({signal_3183, signal_1725}), .clk ( clk ), .r ( Fresh[562] ), .c ({signal_3389, signal_1931}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1917 ( .a ({signal_2529, signal_1071}), .b ({signal_3187, signal_1729}), .clk ( clk ), .r ( Fresh[563] ), .c ({signal_3390, signal_1932}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1919 ( .a ({signal_2393, signal_942}), .b ({signal_3207, signal_1749}), .clk ( clk ), .r ( Fresh[564] ), .c ({signal_3392, signal_1934}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1920 ( .a ({signal_2405, signal_948}), .b ({signal_3208, signal_1750}), .clk ( clk ), .r ( Fresh[565] ), .c ({signal_3393, signal_1935}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1923 ( .a ({signal_2539, signal_1081}), .b ({signal_3209, signal_1751}), .clk ( clk ), .r ( Fresh[566] ), .c ({signal_3396, signal_1938}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1927 ( .a ({signal_2438, signal_980}), .b ({signal_3212, signal_1754}), .clk ( clk ), .r ( Fresh[567] ), .c ({signal_3400, signal_1942}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1932 ( .a ({signal_2417, signal_959}), .b ({signal_3218, signal_1760}), .clk ( clk ), .r ( Fresh[568] ), .c ({signal_3405, signal_1947}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1944 ( .a ({signal_2439, signal_981}), .b ({signal_3222, signal_1764}), .clk ( clk ), .r ( Fresh[569] ), .c ({signal_3417, signal_1959}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1948 ( .a ({signal_3350, signal_1892}), .b ({signal_3421, signal_1963}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1949 ( .a ({signal_3351, signal_1893}), .b ({signal_3422, signal_1964}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1950 ( .a ({signal_3353, signal_1895}), .b ({signal_3423, signal_1965}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1951 ( .a ({signal_3355, signal_1897}), .b ({signal_3424, signal_1966}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1952 ( .a ({signal_3356, signal_1898}), .b ({signal_3425, signal_1967}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1953 ( .a ({signal_3358, signal_1900}), .b ({signal_3426, signal_1968}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1954 ( .a ({signal_3359, signal_1901}), .b ({signal_3427, signal_1969}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1955 ( .a ({signal_3360, signal_1902}), .b ({signal_3428, signal_1970}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1956 ( .a ({signal_3361, signal_1903}), .b ({signal_3429, signal_1971}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1957 ( .a ({signal_3362, signal_1904}), .b ({signal_3430, signal_1972}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1958 ( .a ({signal_3363, signal_1905}), .b ({signal_3431, signal_1973}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1959 ( .a ({signal_3364, signal_1906}), .b ({signal_3432, signal_1974}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1960 ( .a ({signal_3365, signal_1907}), .b ({signal_3433, signal_1975}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1962 ( .a ({signal_3367, signal_1909}), .b ({signal_3435, signal_1977}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1963 ( .a ({signal_3368, signal_1910}), .b ({signal_3436, signal_1978}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1964 ( .a ({signal_3369, signal_1911}), .b ({signal_3437, signal_1979}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1965 ( .a ({signal_3370, signal_1912}), .b ({signal_3438, signal_1980}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1966 ( .a ({signal_3371, signal_1913}), .b ({signal_3439, signal_1981}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1967 ( .a ({signal_3372, signal_1914}), .b ({signal_3440, signal_1982}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1968 ( .a ({signal_3373, signal_1915}), .b ({signal_3441, signal_1983}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1970 ( .a ({signal_3376, signal_1918}), .b ({signal_3443, signal_1985}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1972 ( .a ({signal_3378, signal_1920}), .b ({signal_3445, signal_1987}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1973 ( .a ({signal_3379, signal_1921}), .b ({signal_3446, signal_1988}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1974 ( .a ({signal_3380, signal_1922}), .b ({signal_3447, signal_1989}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1975 ( .a ({signal_3381, signal_1923}), .b ({signal_3448, signal_1990}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1976 ( .a ({signal_3382, signal_1924}), .b ({signal_3449, signal_1991}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1977 ( .a ({signal_3383, signal_1925}), .b ({signal_3450, signal_1992}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1979 ( .a ({signal_3386, signal_1928}), .b ({signal_3452, signal_1994}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1980 ( .a ({signal_3387, signal_1929}), .b ({signal_3453, signal_1995}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1981 ( .a ({signal_3388, signal_1930}), .b ({signal_3454, signal_1996}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1982 ( .a ({signal_3389, signal_1931}), .b ({signal_3455, signal_1997}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1983 ( .a ({signal_3390, signal_1932}), .b ({signal_3456, signal_1998}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1984 ( .a ({signal_3392, signal_1934}), .b ({signal_3457, signal_1999}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1985 ( .a ({signal_3393, signal_1935}), .b ({signal_3458, signal_2000}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1988 ( .a ({signal_3396, signal_1938}), .b ({signal_3461, signal_2003}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1990 ( .a ({signal_3400, signal_1942}), .b ({signal_3463, signal_2005}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1991 ( .a ({signal_3405, signal_1947}), .b ({signal_3464, signal_2006}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1996 ( .a ({signal_3417, signal_1959}), .b ({signal_3469, signal_2011}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2000 ( .a ({signal_3321, signal_1863}), .b ({signal_3052, signal_1594}), .clk ( clk ), .r ( Fresh[570] ), .c ({signal_3473, signal_2015}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2001 ( .a ({signal_3310, signal_1852}), .b ({signal_3023, signal_1565}), .clk ( clk ), .r ( Fresh[571] ), .c ({signal_3474, signal_2016}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2003 ( .a ({signal_3313, signal_1855}), .b ({signal_3314, signal_1856}), .clk ( clk ), .r ( Fresh[572] ), .c ({signal_3476, signal_2018}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2004 ( .a ({signal_2762, signal_1304}), .b ({signal_3316, signal_1858}), .clk ( clk ), .r ( Fresh[573] ), .c ({signal_3477, signal_2019}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2005 ( .a ({signal_2520, signal_1062}), .b ({signal_3317, signal_1859}), .clk ( clk ), .r ( Fresh[574] ), .c ({signal_3478, signal_2020}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2006 ( .a ({signal_2708, signal_1250}), .b ({signal_3318, signal_1860}), .clk ( clk ), .r ( Fresh[575] ), .c ({signal_3479, signal_2021}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2008 ( .a ({signal_2785, signal_1327}), .b ({signal_3322, signal_1864}), .clk ( clk ), .r ( Fresh[576] ), .c ({signal_3481, signal_2023}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2011 ( .a ({signal_2520, signal_1062}), .b ({signal_3323, signal_1865}), .clk ( clk ), .r ( Fresh[577] ), .c ({signal_3484, signal_2026}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2012 ( .a ({signal_3067, signal_1609}), .b ({signal_3325, signal_1867}), .clk ( clk ), .r ( Fresh[578] ), .c ({signal_3485, signal_2027}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2014 ( .a ({signal_3327, signal_1869}), .b ({signal_3146, signal_1688}), .clk ( clk ), .r ( Fresh[579] ), .c ({signal_3487, signal_2029}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2015 ( .a ({signal_3065, signal_1607}), .b ({signal_3329, signal_1871}), .clk ( clk ), .r ( Fresh[580] ), .c ({signal_3488, signal_2030}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2048 ( .a ({signal_3477, signal_2019}), .b ({signal_3521, signal_2063}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2052 ( .a ({signal_3484, signal_2026}), .b ({signal_3525, signal_2067}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1819 ( .a ({signal_3008, signal_1550}), .b ({signal_3145, signal_1687}), .clk ( clk ), .r ( Fresh[581] ), .c ({signal_3292, signal_1834}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1834 ( .a ({signal_3024, signal_1566}), .b ({signal_3168, signal_1710}), .clk ( clk ), .r ( Fresh[582] ), .c ({signal_3307, signal_1849}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1872 ( .a ({signal_3292, signal_1834}), .b ({signal_3345, signal_1887}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1875 ( .a ({signal_3307, signal_1849}), .b ({signal_3348, signal_1890}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1893 ( .a ({signal_2452, signal_994}), .b ({signal_3188, signal_1730}), .clk ( clk ), .r ( Fresh[583] ), .c ({signal_3366, signal_1908}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1902 ( .a ({signal_3225, signal_1767}), .b ({signal_3244, signal_1786}), .clk ( clk ), .r ( Fresh[584] ), .c ({signal_3375, signal_1917}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1904 ( .a ({signal_2452, signal_994}), .b ({signal_3198, signal_1740}), .clk ( clk ), .r ( Fresh[585] ), .c ({signal_3377, signal_1919}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1911 ( .a ({signal_3248, signal_1790}), .b ({signal_3062, signal_1604}), .clk ( clk ), .r ( Fresh[586] ), .c ({signal_3384, signal_1926}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1912 ( .a ({signal_2748, signal_1290}), .b ({signal_3250, signal_1792}), .clk ( clk ), .r ( Fresh[587] ), .c ({signal_3385, signal_1927}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1918 ( .a ({signal_2812, signal_1354}), .b ({signal_3262, signal_1804}), .clk ( clk ), .r ( Fresh[588] ), .c ({signal_3391, signal_1933}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1921 ( .a ({signal_2692, signal_1234}), .b ({signal_3264, signal_1806}), .clk ( clk ), .r ( Fresh[589] ), .c ({signal_3394, signal_1936}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1922 ( .a ({signal_3266, signal_1808}), .b ({signal_3267, signal_1809}), .clk ( clk ), .r ( Fresh[590] ), .c ({signal_3395, signal_1937}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1924 ( .a ({signal_2435, signal_977}), .b ({signal_3210, signal_1752}), .clk ( clk ), .r ( Fresh[591] ), .c ({signal_3397, signal_1939}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1925 ( .a ({signal_3034, signal_1576}), .b ({signal_3273, signal_1815}), .clk ( clk ), .r ( Fresh[592] ), .c ({signal_3398, signal_1940}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1926 ( .a ({signal_3040, signal_1582}), .b ({signal_3211, signal_1753}), .clk ( clk ), .r ( Fresh[593] ), .c ({signal_3399, signal_1941}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1928 ( .a ({signal_2771, signal_1313}), .b ({signal_3277, signal_1819}), .clk ( clk ), .r ( Fresh[594] ), .c ({signal_3401, signal_1943}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1929 ( .a ({signal_3247, signal_1789}), .b ({signal_3090, signal_1632}), .clk ( clk ), .r ( Fresh[595] ), .c ({signal_3402, signal_1944}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1930 ( .a ({signal_3214, signal_1756}), .b ({signal_3215, signal_1757}), .clk ( clk ), .r ( Fresh[596] ), .c ({signal_3403, signal_1945}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1931 ( .a ({signal_3055, signal_1597}), .b ({signal_3217, signal_1759}), .clk ( clk ), .r ( Fresh[597] ), .c ({signal_3404, signal_1946}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1933 ( .a ({signal_2793, signal_1335}), .b ({signal_3285, signal_1827}), .clk ( clk ), .r ( Fresh[598] ), .c ({signal_3406, signal_1948}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1934 ( .a ({signal_3053, signal_1595}), .b ({signal_3291, signal_1833}), .clk ( clk ), .r ( Fresh[599] ), .c ({signal_3407, signal_1949}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1935 ( .a ({signal_3009, signal_1551}), .b ({signal_3293, signal_1835}), .clk ( clk ), .r ( Fresh[600] ), .c ({signal_3408, signal_1950}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1936 ( .a ({signal_3219, signal_1761}), .b ({signal_3294, signal_1836}), .clk ( clk ), .r ( Fresh[601] ), .c ({signal_3409, signal_1951}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1937 ( .a ({signal_3071, signal_1613}), .b ({signal_3213, signal_1755}), .clk ( clk ), .r ( Fresh[602] ), .c ({signal_3410, signal_1952}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1938 ( .a ({signal_3148, signal_1690}), .b ({signal_3295, signal_1837}), .clk ( clk ), .r ( Fresh[603] ), .c ({signal_3411, signal_1953}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1939 ( .a ({signal_3013, signal_1555}), .b ({signal_3296, signal_1838}), .clk ( clk ), .r ( Fresh[604] ), .c ({signal_3412, signal_1954}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1940 ( .a ({signal_2519, signal_1061}), .b ({signal_3298, signal_1840}), .clk ( clk ), .r ( Fresh[605] ), .c ({signal_3413, signal_1955}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1941 ( .a ({signal_3020, signal_1562}), .b ({signal_3221, signal_1763}), .clk ( clk ), .r ( Fresh[606] ), .c ({signal_3414, signal_1956}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1942 ( .a ({signal_3152, signal_1694}), .b ({signal_3299, signal_1841}), .clk ( clk ), .r ( Fresh[607] ), .c ({signal_3415, signal_1957}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1943 ( .a ({signal_3261, signal_1803}), .b ({signal_3094, signal_1636}), .clk ( clk ), .r ( Fresh[608] ), .c ({signal_3416, signal_1958}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1945 ( .a ({signal_3283, signal_1825}), .b ({signal_3304, signal_1846}), .clk ( clk ), .r ( Fresh[609] ), .c ({signal_3418, signal_1960}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1946 ( .a ({signal_3026, signal_1568}), .b ({signal_3223, signal_1765}), .clk ( clk ), .r ( Fresh[610] ), .c ({signal_3419, signal_1961}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1947 ( .a ({signal_3254, signal_1796}), .b ({signal_3305, signal_1847}), .clk ( clk ), .r ( Fresh[611] ), .c ({signal_3420, signal_1962}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1961 ( .a ({signal_3366, signal_1908}), .b ({signal_3434, signal_1976}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1969 ( .a ({signal_3375, signal_1917}), .b ({signal_3442, signal_1984}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1971 ( .a ({signal_3377, signal_1919}), .b ({signal_3444, signal_1986}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1978 ( .a ({signal_3385, signal_1927}), .b ({signal_3451, signal_1993}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1986 ( .a ({signal_3394, signal_1936}), .b ({signal_3459, signal_2001}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1987 ( .a ({signal_3395, signal_1937}), .b ({signal_3460, signal_2002}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1989 ( .a ({signal_3397, signal_1939}), .b ({signal_3462, signal_2004}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1992 ( .a ({signal_3407, signal_1949}), .b ({signal_3465, signal_2007}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1993 ( .a ({signal_3409, signal_1951}), .b ({signal_3466, signal_2008}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1994 ( .a ({signal_3415, signal_1957}), .b ({signal_3467, signal_2009}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1995 ( .a ({signal_3416, signal_1958}), .b ({signal_3468, signal_2010}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1997 ( .a ({signal_3418, signal_1960}), .b ({signal_3470, signal_2012}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_1998 ( .a ({signal_3420, signal_1962}), .b ({signal_3471, signal_2013}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_1999 ( .a ({signal_3315, signal_1857}), .b ({signal_2819, signal_1361}), .clk ( clk ), .r ( Fresh[612] ), .c ({signal_3472, signal_2014}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2002 ( .a ({signal_3311, signal_1853}), .b ({signal_3232, signal_1774}), .clk ( clk ), .r ( Fresh[613] ), .c ({signal_3475, signal_2017}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2007 ( .a ({signal_2415, signal_957}), .b ({signal_3352, signal_1894}), .clk ( clk ), .r ( Fresh[614] ), .c ({signal_3480, signal_2022}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2009 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_3354, signal_1896}), .clk ( clk ), .r ( Fresh[615] ), .c ({signal_3482, signal_2024}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2010 ( .a ({signal_2447, signal_989}), .b ({signal_3357, signal_1899}), .clk ( clk ), .r ( Fresh[616] ), .c ({signal_3483, signal_2025}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2013 ( .a ({signal_2442, signal_984}), .b ({signal_3326, signal_1868}), .clk ( clk ), .r ( Fresh[617] ), .c ({signal_3486, signal_2028}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2016 ( .a ({signal_2449, signal_991}), .b ({signal_3332, signal_1874}), .clk ( clk ), .r ( Fresh[618] ), .c ({signal_3489, signal_2031}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2017 ( .a ({signal_2456, signal_998}), .b ({signal_3333, signal_1875}), .clk ( clk ), .r ( Fresh[619] ), .c ({signal_3490, signal_2032}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2018 ( .a ({signal_2405, signal_948}), .b ({signal_3334, signal_1876}), .clk ( clk ), .r ( Fresh[620] ), .c ({signal_3491, signal_2033}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2019 ( .a ({signal_3312, signal_1854}), .b ({signal_3271, signal_1813}), .clk ( clk ), .r ( Fresh[621] ), .c ({signal_3492, signal_2034}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2020 ( .a ({signal_2417, signal_959}), .b ({signal_3335, signal_1877}), .clk ( clk ), .r ( Fresh[622] ), .c ({signal_3493, signal_2035}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2021 ( .a ({signal_2438, signal_980}), .b ({signal_3336, signal_1878}), .clk ( clk ), .r ( Fresh[623] ), .c ({signal_3494, signal_2036}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2022 ( .a ({signal_2419, signal_961}), .b ({signal_3337, signal_1879}), .clk ( clk ), .r ( Fresh[624] ), .c ({signal_3495, signal_2037}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2023 ( .a ({signal_2445, signal_987}), .b ({signal_3338, signal_1880}), .clk ( clk ), .r ( Fresh[625] ), .c ({signal_3496, signal_2038}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2024 ( .a ({signal_2459, signal_1001}), .b ({signal_3339, signal_1881}), .clk ( clk ), .r ( Fresh[626] ), .c ({signal_3497, signal_2039}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2025 ( .a ({signal_3320, signal_1862}), .b ({signal_3340, signal_1882}), .clk ( clk ), .r ( Fresh[627] ), .c ({signal_3498, signal_2040}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2026 ( .a ({signal_3284, signal_1826}), .b ({signal_3374, signal_1916}), .clk ( clk ), .r ( Fresh[628] ), .c ({signal_3499, signal_2041}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2028 ( .a ({signal_2401, signal_946}), .b ({signal_3341, signal_1883}), .clk ( clk ), .r ( Fresh[629] ), .c ({signal_3501, signal_2043}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2029 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_3342, signal_1884}), .clk ( clk ), .r ( Fresh[630] ), .c ({signal_3502, signal_2044}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2030 ( .a ({signal_3324, signal_1866}), .b ({signal_3288, signal_1830}), .clk ( clk ), .r ( Fresh[631] ), .c ({signal_3503, signal_2045}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2031 ( .a ({signal_2462, signal_1004}), .b ({signal_3344, signal_1886}), .clk ( clk ), .r ( Fresh[632] ), .c ({signal_3504, signal_2046}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2033 ( .a ({signal_3331, signal_1873}), .b ({signal_3297, signal_1839}), .clk ( clk ), .r ( Fresh[633] ), .c ({signal_3506, signal_2048}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2034 ( .a ({signal_3309, signal_1851}), .b ({signal_3276, signal_1818}), .clk ( clk ), .r ( Fresh[634] ), .c ({signal_3507, signal_2049}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2035 ( .a ({signal_2538, signal_1080}), .b ({signal_3346, signal_1888}), .clk ( clk ), .r ( Fresh[635] ), .c ({signal_3508, signal_2050}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2036 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_3347, signal_1889}), .clk ( clk ), .r ( Fresh[636] ), .c ({signal_3509, signal_2051}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2046 ( .a ({signal_3472, signal_2014}), .b ({signal_3519, signal_2061}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2047 ( .a ({signal_3475, signal_2017}), .b ({signal_3520, signal_2062}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2049 ( .a ({signal_3480, signal_2022}), .b ({signal_3522, signal_2064}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2050 ( .a ({signal_3482, signal_2024}), .b ({signal_3523, signal_2065}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2051 ( .a ({signal_3483, signal_2025}), .b ({signal_3524, signal_2066}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2053 ( .a ({signal_3486, signal_2028}), .b ({signal_3526, signal_2068}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2054 ( .a ({signal_3489, signal_2031}), .b ({signal_3527, signal_2069}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2055 ( .a ({signal_3490, signal_2032}), .b ({signal_3528, signal_2070}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2056 ( .a ({signal_3491, signal_2033}), .b ({signal_3529, signal_2071}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2057 ( .a ({signal_3492, signal_2034}), .b ({signal_3530, signal_2072}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2058 ( .a ({signal_3493, signal_2035}), .b ({signal_3531, signal_2073}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2059 ( .a ({signal_3494, signal_2036}), .b ({signal_3532, signal_2074}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2060 ( .a ({signal_3495, signal_2037}), .b ({signal_3533, signal_2075}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2061 ( .a ({signal_3496, signal_2038}), .b ({signal_3534, signal_2076}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2062 ( .a ({signal_3497, signal_2039}), .b ({signal_3535, signal_2077}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2063 ( .a ({signal_3499, signal_2041}), .b ({signal_3536, signal_2078}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2065 ( .a ({signal_3501, signal_2043}), .b ({signal_3538, signal_2080}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2066 ( .a ({signal_3502, signal_2044}), .b ({signal_3539, signal_2081}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2067 ( .a ({signal_3504, signal_2046}), .b ({signal_3540, signal_2082}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2069 ( .a ({signal_3506, signal_2048}), .b ({signal_3542, signal_2084}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2070 ( .a ({signal_3508, signal_2050}), .b ({signal_3543, signal_2085}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2071 ( .a ({signal_3509, signal_2051}), .b ({signal_3544, signal_2086}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2074 ( .a ({signal_3435, signal_1977}), .b ({signal_2823, signal_1365}), .clk ( clk ), .r ( Fresh[637] ), .c ({signal_3547, signal_2089}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2075 ( .a ({signal_3029, signal_1571}), .b ({signal_3422, signal_1964}), .clk ( clk ), .r ( Fresh[638] ), .c ({signal_3548, signal_2090}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2076 ( .a ({signal_2700, signal_1242}), .b ({signal_3473, signal_2015}), .clk ( clk ), .r ( Fresh[639] ), .c ({signal_3549, signal_2091}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2077 ( .a ({signal_2998, signal_1540}), .b ({signal_3427, signal_1969}), .clk ( clk ), .r ( Fresh[640] ), .c ({signal_3550, signal_2092}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2078 ( .a ({signal_3421, signal_1963}), .b ({signal_3330, signal_1872}), .clk ( clk ), .r ( Fresh[641] ), .c ({signal_3551, signal_2093}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2079 ( .a ({signal_3431, signal_1973}), .b ({signal_3432, signal_1974}), .clk ( clk ), .r ( Fresh[642] ), .c ({signal_3552, signal_2094}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2080 ( .a ({signal_2754, signal_1296}), .b ({signal_3476, signal_2018}), .clk ( clk ), .r ( Fresh[643] ), .c ({signal_3553, signal_2095}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2081 ( .a ({signal_2766, signal_1308}), .b ({signal_3478, signal_2020}), .clk ( clk ), .r ( Fresh[644] ), .c ({signal_3554, signal_2096}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2082 ( .a ({signal_2709, signal_1251}), .b ({signal_3479, signal_2021}), .clk ( clk ), .r ( Fresh[645] ), .c ({signal_3555, signal_2097}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2083 ( .a ({signal_3041, signal_1583}), .b ({signal_3439, signal_1981}), .clk ( clk ), .r ( Fresh[646] ), .c ({signal_3556, signal_2098}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2085 ( .a ({signal_2784, signal_1326}), .b ({signal_3443, signal_1985}), .clk ( clk ), .r ( Fresh[647] ), .c ({signal_3558, signal_2100}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2086 ( .a ({signal_2719, signal_1261}), .b ({signal_3481, signal_2023}), .clk ( clk ), .r ( Fresh[648] ), .c ({signal_3559, signal_2101}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2087 ( .a ({signal_3349, signal_1891}), .b ({signal_3447, signal_1989}), .clk ( clk ), .r ( Fresh[649] ), .c ({signal_3560, signal_2102}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2088 ( .a ({signal_3448, signal_1990}), .b ({signal_3449, signal_1991}), .clk ( clk ), .r ( Fresh[650] ), .c ({signal_3561, signal_2103}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2089 ( .a ({signal_3058, signal_1600}), .b ({signal_3450, signal_1992}), .clk ( clk ), .r ( Fresh[651] ), .c ({signal_3562, signal_2104}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2091 ( .a ({signal_3485, signal_2027}), .b ({signal_3343, signal_1885}), .clk ( clk ), .r ( Fresh[652] ), .c ({signal_3564, signal_2106}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2092 ( .a ({signal_2729, signal_1271}), .b ({signal_3452, signal_1994}), .clk ( clk ), .r ( Fresh[653] ), .c ({signal_3565, signal_2107}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2093 ( .a ({signal_3328, signal_1870}), .b ({signal_3453, signal_1995}), .clk ( clk ), .r ( Fresh[654] ), .c ({signal_3566, signal_2108}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2094 ( .a ({signal_3260, signal_1802}), .b ({signal_3454, signal_1996}), .clk ( clk ), .r ( Fresh[655] ), .c ({signal_3567, signal_2109}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2095 ( .a ({signal_3429, signal_1971}), .b ({signal_3455, signal_1997}), .clk ( clk ), .r ( Fresh[656] ), .c ({signal_3568, signal_2110}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2096 ( .a ({signal_3214, signal_1756}), .b ({signal_3456, signal_1998}), .clk ( clk ), .r ( Fresh[657] ), .c ({signal_3569, signal_2111}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2097 ( .a ({signal_3430, signal_1972}), .b ({signal_3090, signal_1632}), .clk ( clk ), .r ( Fresh[658] ), .c ({signal_3570, signal_2112}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2099 ( .a ({signal_3156, signal_1698}), .b ({signal_3458, signal_2000}), .clk ( clk ), .r ( Fresh[659] ), .c ({signal_3572, signal_2114}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2101 ( .a ({signal_3433, signal_1975}), .b ({signal_3461, signal_2003}), .clk ( clk ), .r ( Fresh[660] ), .c ({signal_3574, signal_2116}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2104 ( .a ({signal_2770, signal_1312}), .b ({signal_3463, signal_2005}), .clk ( clk ), .r ( Fresh[661] ), .c ({signal_3577, signal_2119}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2110 ( .a ({signal_3487, signal_2029}), .b ({signal_3306, signal_1848}), .clk ( clk ), .r ( Fresh[662] ), .c ({signal_3583, signal_2125}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2124 ( .a ({signal_3547, signal_2089}), .b ({signal_3597, signal_2139}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2125 ( .a ({signal_3549, signal_2091}), .b ({signal_3598, signal_2140}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2126 ( .a ({signal_3550, signal_2092}), .b ({signal_3599, signal_2141}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2127 ( .a ({signal_3554, signal_2096}), .b ({signal_3600, signal_2142}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2128 ( .a ({signal_3555, signal_2097}), .b ({signal_3601, signal_2143}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2130 ( .a ({signal_3559, signal_2101}), .b ({signal_3603, signal_2145}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2133 ( .a ({signal_3577, signal_2119}), .b ({signal_3606, signal_2148}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2135 ( .a ({signal_3583, signal_2125}), .b ({signal_3608, signal_2150}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2144 ( .a ({signal_2420, signal_962}), .b ({signal_3521, signal_2063}), .clk ( clk ), .r ( Fresh[663] ), .c ({signal_3617, signal_2159}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2148 ( .a ({signal_2451, signal_993}), .b ({signal_3525, signal_2067}), .clk ( clk ), .r ( Fresh[664] ), .c ({signal_3621, signal_2163}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2185 ( .a ({signal_3617, signal_2159}), .b ({signal_3658, signal_2200}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2186 ( .a ({signal_3621, signal_2163}), .b ({signal_3659, signal_2201}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2027 ( .a ({signal_2998, signal_1540}), .b ({signal_3384, signal_1926}), .clk ( clk ), .r ( Fresh[665] ), .c ({signal_3500, signal_2042}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2032 ( .a ({signal_2443, signal_985}), .b ({signal_3345, signal_1887}), .clk ( clk ), .r ( Fresh[666] ), .c ({signal_3505, signal_2047}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2037 ( .a ({signal_2706, signal_1248}), .b ({signal_3398, signal_1940}), .clk ( clk ), .r ( Fresh[667] ), .c ({signal_3510, signal_2052}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2038 ( .a ({signal_2772, signal_1314}), .b ({signal_3401, signal_1943}), .clk ( clk ), .r ( Fresh[668] ), .c ({signal_3511, signal_2053}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2039 ( .a ({signal_2995, signal_1537}), .b ({signal_3404, signal_1946}), .clk ( clk ), .r ( Fresh[669] ), .c ({signal_3512, signal_2054}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2040 ( .a ({signal_2794, signal_1336}), .b ({signal_3406, signal_1948}), .clk ( clk ), .r ( Fresh[670] ), .c ({signal_3513, signal_2055}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2041 ( .a ({signal_3010, signal_1552}), .b ({signal_3408, signal_1950}), .clk ( clk ), .r ( Fresh[671] ), .c ({signal_3514, signal_2056}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2042 ( .a ({signal_3076, signal_1618}), .b ({signal_3412, signal_1954}), .clk ( clk ), .r ( Fresh[672] ), .c ({signal_3515, signal_2057}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2043 ( .a ({signal_3018, signal_1560}), .b ({signal_3413, signal_1955}), .clk ( clk ), .r ( Fresh[673] ), .c ({signal_3516, signal_2058}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2044 ( .a ({signal_3080, signal_1622}), .b ({signal_3414, signal_1956}), .clk ( clk ), .r ( Fresh[674] ), .c ({signal_3517, signal_2059}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2045 ( .a ({signal_2991, signal_1533}), .b ({signal_3419, signal_1961}), .clk ( clk ), .r ( Fresh[675] ), .c ({signal_3518, signal_2060}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2064 ( .a ({signal_3500, signal_2042}), .b ({signal_3537, signal_2079}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2068 ( .a ({signal_3505, signal_2047}), .b ({signal_3541, signal_2083}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2072 ( .a ({signal_3510, signal_2052}), .b ({signal_3545, signal_2087}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2073 ( .a ({signal_3516, signal_2058}), .b ({signal_3546, signal_2088}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2084 ( .a ({signal_2467, signal_1009}), .b ({signal_3442, signal_1984}), .clk ( clk ), .r ( Fresh[676] ), .c ({signal_3557, signal_2099}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2090 ( .a ({signal_2408, signal_950}), .b ({signal_3451, signal_1993}), .clk ( clk ), .r ( Fresh[677] ), .c ({signal_3563, signal_2105}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2098 ( .a ({signal_3391, signal_1933}), .b ({signal_3457, signal_1999}), .clk ( clk ), .r ( Fresh[678] ), .c ({signal_3571, signal_2113}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2100 ( .a ({signal_2417, signal_959}), .b ({signal_3459, signal_2001}), .clk ( clk ), .r ( Fresh[679] ), .c ({signal_3573, signal_2115}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2102 ( .a ({signal_3269, signal_1811}), .b ({signal_3462, signal_2004}), .clk ( clk ), .r ( Fresh[680] ), .c ({signal_3575, signal_2117}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2103 ( .a ({signal_3438, signal_1980}), .b ({signal_3399, signal_1941}), .clk ( clk ), .r ( Fresh[681] ), .c ({signal_3576, signal_2118}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2105 ( .a ({signal_3441, signal_1983}), .b ({signal_3399, signal_1941}), .clk ( clk ), .r ( Fresh[682] ), .c ({signal_3578, signal_2120}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2106 ( .a ({signal_3049, signal_1591}), .b ({signal_3498, signal_2040}), .clk ( clk ), .r ( Fresh[683] ), .c ({signal_3579, signal_2121}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2107 ( .a ({signal_3423, signal_1965}), .b ({signal_3402, signal_1944}), .clk ( clk ), .r ( Fresh[684] ), .c ({signal_3580, signal_2122}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2108 ( .a ({signal_3426, signal_1968}), .b ({signal_3503, signal_2045}), .clk ( clk ), .r ( Fresh[685] ), .c ({signal_3581, signal_2123}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2109 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_3465, signal_2007}), .clk ( clk ), .r ( Fresh[686] ), .c ({signal_3582, signal_2124}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2111 ( .a ({signal_2453, signal_995}), .b ({signal_3466, signal_2008}), .clk ( clk ), .r ( Fresh[687] ), .c ({signal_3584, signal_2126}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2112 ( .a ({signal_3428, signal_1970}), .b ({signal_3410, signal_1952}), .clk ( clk ), .r ( Fresh[688] ), .c ({signal_3585, signal_2127}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2113 ( .a ({signal_3079, signal_1621}), .b ({signal_3507, signal_2049}), .clk ( clk ), .r ( Fresh[689] ), .c ({signal_3586, signal_2128}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2114 ( .a ({signal_2442, signal_984}), .b ({signal_3467, signal_2009}), .clk ( clk ), .r ( Fresh[690] ), .c ({signal_3587, signal_2129}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2115 ( .a ({signal_2467, signal_1009}), .b ({signal_3468, signal_2010}), .clk ( clk ), .r ( Fresh[691] ), .c ({signal_3588, signal_2130}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2117 ( .a ({signal_2462, signal_1004}), .b ({signal_3470, signal_2012}), .clk ( clk ), .r ( Fresh[692] ), .c ({signal_3590, signal_2132}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2120 ( .a ({signal_2408, signal_950}), .b ({signal_3471, signal_2013}), .clk ( clk ), .r ( Fresh[693] ), .c ({signal_3593, signal_2135}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2129 ( .a ({signal_3557, signal_2099}), .b ({signal_3602, signal_2144}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2131 ( .a ({signal_3563, signal_2105}), .b ({signal_3604, signal_2146}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2132 ( .a ({signal_3573, signal_2115}), .b ({signal_3605, signal_2147}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2134 ( .a ({signal_3582, signal_2124}), .b ({signal_3607, signal_2149}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2136 ( .a ({signal_3584, signal_2126}), .b ({signal_3609, signal_2151}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2137 ( .a ({signal_3587, signal_2129}), .b ({signal_3610, signal_2152}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2138 ( .a ({signal_3588, signal_2130}), .b ({signal_3611, signal_2153}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2139 ( .a ({signal_3590, signal_2132}), .b ({signal_3612, signal_2154}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2141 ( .a ({signal_3593, signal_2135}), .b ({signal_3614, signal_2156}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2142 ( .a ({signal_2756, signal_1298}), .b ({signal_3519, signal_2061}), .clk ( clk ), .r ( Fresh[694] ), .c ({signal_3615, signal_2157}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2143 ( .a ({signal_2439, signal_981}), .b ({signal_3520, signal_2062}), .clk ( clk ), .r ( Fresh[695] ), .c ({signal_3616, signal_2158}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2145 ( .a ({signal_3213, signal_1755}), .b ({signal_3548, signal_2090}), .clk ( clk ), .r ( Fresh[696] ), .c ({signal_3618, signal_2160}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2146 ( .a ({signal_3523, signal_2065}), .b ({signal_3445, signal_1987}), .clk ( clk ), .r ( Fresh[697] ), .c ({signal_3619, signal_2161}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2147 ( .a ({signal_3064, signal_1606}), .b ({signal_3524, signal_2066}), .clk ( clk ), .r ( Fresh[698] ), .c ({signal_3620, signal_2162}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2149 ( .a ({signal_3149, signal_1691}), .b ({signal_3551, signal_2093}), .clk ( clk ), .r ( Fresh[699] ), .c ({signal_3622, signal_2164}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2150 ( .a ({signal_3028, signal_1570}), .b ({signal_3552, signal_2094}), .clk ( clk ), .r ( Fresh[700] ), .c ({signal_3623, signal_2165}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2151 ( .a ({signal_2459, signal_1001}), .b ({signal_3530, signal_2072}), .clk ( clk ), .r ( Fresh[701] ), .c ({signal_3624, signal_2166}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2152 ( .a ({signal_2522, signal_1064}), .b ({signal_3553, signal_2095}), .clk ( clk ), .r ( Fresh[702] ), .c ({signal_3625, signal_2167}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2153 ( .a ({signal_3042, signal_1584}), .b ({signal_3556, signal_2098}), .clk ( clk ), .r ( Fresh[703] ), .c ({signal_3626, signal_2168}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2154 ( .a ({signal_2774, signal_1316}), .b ({signal_3533, signal_2075}), .clk ( clk ), .r ( Fresh[704] ), .c ({signal_3627, signal_2169}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2155 ( .a ({signal_3522, signal_2064}), .b ({signal_3534, signal_2076}), .clk ( clk ), .r ( Fresh[705] ), .c ({signal_3628, signal_2170}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2156 ( .a ({signal_3048, signal_1590}), .b ({signal_3535, signal_2077}), .clk ( clk ), .r ( Fresh[706] ), .c ({signal_3629, signal_2171}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2157 ( .a ({signal_2443, signal_985}), .b ({signal_3536, signal_2078}), .clk ( clk ), .r ( Fresh[707] ), .c ({signal_3630, signal_2172}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2158 ( .a ({signal_3133, signal_1675}), .b ({signal_3558, signal_2100}), .clk ( clk ), .r ( Fresh[708] ), .c ({signal_3631, signal_2173}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2159 ( .a ({signal_3056, signal_1598}), .b ({signal_3560, signal_2102}), .clk ( clk ), .r ( Fresh[709] ), .c ({signal_3632, signal_2174}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2160 ( .a ({signal_3424, signal_1966}), .b ({signal_3561, signal_2103}), .clk ( clk ), .r ( Fresh[710] ), .c ({signal_3633, signal_2175}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2161 ( .a ({signal_3059, signal_1601}), .b ({signal_3562, signal_2104}), .clk ( clk ), .r ( Fresh[711] ), .c ({signal_3634, signal_2176}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2163 ( .a ({signal_3001, signal_1543}), .b ({signal_3538, signal_2080}), .clk ( clk ), .r ( Fresh[712] ), .c ({signal_3636, signal_2178}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2164 ( .a ({signal_2747, signal_1289}), .b ({signal_3565, signal_2107}), .clk ( clk ), .r ( Fresh[713] ), .c ({signal_3637, signal_2179}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2165 ( .a ({signal_3566, signal_2108}), .b ({signal_3411, signal_1953}), .clk ( clk ), .r ( Fresh[714] ), .c ({signal_3638, signal_2180}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2166 ( .a ({signal_2443, signal_985}), .b ({signal_3542, signal_2084}), .clk ( clk ), .r ( Fresh[715] ), .c ({signal_3639, signal_2181}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2167 ( .a ({signal_3543, signal_2085}), .b ({signal_3469, signal_2011}), .clk ( clk ), .r ( Fresh[716] ), .c ({signal_3640, signal_2182}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2168 ( .a ({signal_3301, signal_1843}), .b ({signal_3570, signal_2112}), .clk ( clk ), .r ( Fresh[717] ), .c ({signal_3641, signal_2183}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2169 ( .a ({signal_3083, signal_1625}), .b ({signal_3544, signal_2086}), .clk ( clk ), .r ( Fresh[718] ), .c ({signal_3642, signal_2184}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2171 ( .a ({signal_2817, signal_1359}), .b ({signal_3572, signal_2114}), .clk ( clk ), .r ( Fresh[719] ), .c ({signal_3644, signal_2186}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2184 ( .a ({signal_3616, signal_2158}), .b ({signal_3657, signal_2199}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2187 ( .a ({signal_3624, signal_2166}), .b ({signal_3660, signal_2202}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2188 ( .a ({signal_3630, signal_2172}), .b ({signal_3661, signal_2203}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2189 ( .a ({signal_3632, signal_2174}), .b ({signal_3662, signal_2204}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2191 ( .a ({signal_3637, signal_2179}), .b ({signal_3664, signal_2206}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2192 ( .a ({signal_3638, signal_2180}), .b ({signal_3665, signal_2207}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2193 ( .a ({signal_3639, signal_2181}), .b ({signal_3666, signal_2208}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2194 ( .a ({signal_3644, signal_2186}), .b ({signal_3667, signal_2209}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2201 ( .a ({signal_2765, signal_1307}), .b ({signal_3597, signal_2139}), .clk ( clk ), .r ( Fresh[720] ), .c ({signal_3674, signal_2216}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2202 ( .a ({signal_2455, signal_997}), .b ({signal_3598, signal_2140}), .clk ( clk ), .r ( Fresh[721] ), .c ({signal_3675, signal_2217}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2203 ( .a ({signal_2403, signal_947}), .b ({signal_3599, signal_2141}), .clk ( clk ), .r ( Fresh[722] ), .c ({signal_3676, signal_2218}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2204 ( .a ({signal_2443, signal_985}), .b ({signal_3600, signal_2142}), .clk ( clk ), .r ( Fresh[723] ), .c ({signal_3677, signal_2219}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2205 ( .a ({signal_2445, signal_987}), .b ({signal_3601, signal_2143}), .clk ( clk ), .r ( Fresh[724] ), .c ({signal_3678, signal_2220}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2206 ( .a ({signal_2442, signal_984}), .b ({signal_3603, signal_2145}), .clk ( clk ), .r ( Fresh[725] ), .c ({signal_3679, signal_2221}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2213 ( .a ({signal_2401, signal_946}), .b ({signal_3606, signal_2148}), .clk ( clk ), .r ( Fresh[726] ), .c ({signal_3686, signal_2228}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2221 ( .a ({signal_2455, signal_997}), .b ({signal_3608, signal_2150}), .clk ( clk ), .r ( Fresh[727] ), .c ({signal_3694, signal_2236}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2233 ( .a ({signal_3674, signal_2216}), .b ({signal_3706, signal_2248}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2234 ( .a ({signal_3675, signal_2217}), .b ({signal_3707, signal_2249}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2235 ( .a ({signal_3676, signal_2218}), .b ({signal_3708, signal_2250}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2236 ( .a ({signal_3677, signal_2219}), .b ({signal_3709, signal_2251}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2237 ( .a ({signal_3678, signal_2220}), .b ({signal_3710, signal_2252}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2238 ( .a ({signal_3679, signal_2221}), .b ({signal_3711, signal_2253}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2240 ( .a ({signal_3686, signal_2228}), .b ({signal_3713, signal_2255}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2242 ( .a ({signal_3694, signal_2236}), .b ({signal_3715, signal_2257}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2248 ( .a ({signal_3532, signal_2074}), .b ({signal_3658, signal_2200}), .clk ( clk ), .r ( Fresh[728] ), .c ({signal_3721, signal_2263}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2116 ( .a ({signal_2773, signal_1315}), .b ({signal_3511, signal_2053}), .clk ( clk ), .r ( Fresh[729] ), .c ({signal_3589, signal_2131}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2118 ( .a ({signal_3216, signal_1758}), .b ({signal_3512, signal_2054}), .clk ( clk ), .r ( Fresh[730] ), .c ({signal_3591, signal_2133}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2119 ( .a ({signal_3103, signal_1645}), .b ({signal_3513, signal_2055}), .clk ( clk ), .r ( Fresh[731] ), .c ({signal_3592, signal_2134}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2121 ( .a ({signal_3074, signal_1616}), .b ({signal_3515, signal_2057}), .clk ( clk ), .r ( Fresh[732] ), .c ({signal_3594, signal_2136}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2122 ( .a ({signal_3220, signal_1762}), .b ({signal_3517, signal_2059}), .clk ( clk ), .r ( Fresh[733] ), .c ({signal_3595, signal_2137}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2123 ( .a ({signal_2992, signal_1534}), .b ({signal_3518, signal_2060}), .clk ( clk ), .r ( Fresh[734] ), .c ({signal_3596, signal_2138}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2140 ( .a ({signal_3592, signal_2134}), .b ({signal_3613, signal_2155}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2162 ( .a ({SI_s1[2], SI_s0[2]}), .b ({signal_3537, signal_2079}), .clk ( clk ), .r ( Fresh[735] ), .c ({signal_3635, signal_2177}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2170 ( .a ({signal_3303, signal_1845}), .b ({signal_3571, signal_2113}), .clk ( clk ), .r ( Fresh[736] ), .c ({signal_3643, signal_2185}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2172 ( .a ({signal_3529, signal_2071}), .b ({signal_3575, signal_2117}), .clk ( clk ), .r ( Fresh[737] ), .c ({signal_3645, signal_2187}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2173 ( .a ({signal_2459, signal_1001}), .b ({signal_3545, signal_2087}), .clk ( clk ), .r ( Fresh[738] ), .c ({signal_3646, signal_2188}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2174 ( .a ({signal_3308, signal_1850}), .b ({signal_3579, signal_2121}), .clk ( clk ), .r ( Fresh[739] ), .c ({signal_3647, signal_2189}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2175 ( .a ({signal_3089, signal_1631}), .b ({signal_3580, signal_2122}), .clk ( clk ), .r ( Fresh[740] ), .c ({signal_3648, signal_2190}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2176 ( .a ({signal_3141, signal_1683}), .b ({signal_3581, signal_2123}), .clk ( clk ), .r ( Fresh[741] ), .c ({signal_3649, signal_2191}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2177 ( .a ({signal_3541, signal_2083}), .b ({signal_3514, signal_2056}), .clk ( clk ), .r ( Fresh[742] ), .c ({signal_3650, signal_2192}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2178 ( .a ({signal_2408, signal_950}), .b ({signal_3546, signal_2088}), .clk ( clk ), .r ( Fresh[743] ), .c ({signal_3651, signal_2193}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2179 ( .a ({signal_3268, signal_1810}), .b ({signal_3586, signal_2128}), .clk ( clk ), .r ( Fresh[744] ), .c ({signal_3652, signal_2194}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2190 ( .a ({signal_3635, signal_2177}), .b ({signal_3663, signal_2205}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2195 ( .a ({signal_3646, signal_2188}), .b ({signal_3668, signal_2210}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2196 ( .a ({signal_3648, signal_2190}), .b ({signal_3669, signal_2211}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2197 ( .a ({signal_3649, signal_2191}), .b ({signal_3670, signal_2212}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2198 ( .a ({signal_3651, signal_2193}), .b ({signal_3671, signal_2213}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2200 ( .a ({signal_2757, signal_1299}), .b ({signal_3615, signal_2157}), .clk ( clk ), .r ( Fresh[745] ), .c ({signal_3673, signal_2215}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2207 ( .a ({signal_3539, signal_2081}), .b ({signal_3604, signal_2146}), .clk ( clk ), .r ( Fresh[746] ), .c ({signal_3680, signal_2222}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2208 ( .a ({signal_3015, signal_1557}), .b ({signal_3622, signal_2164}), .clk ( clk ), .r ( Fresh[747] ), .c ({signal_3681, signal_2223}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2209 ( .a ({signal_3527, signal_2069}), .b ({signal_3605, signal_2147}), .clk ( clk ), .r ( Fresh[748] ), .c ({signal_3682, signal_2224}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2210 ( .a ({signal_2697, signal_1239}), .b ({signal_3623, signal_2165}), .clk ( clk ), .r ( Fresh[749] ), .c ({signal_3683, signal_2225}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2211 ( .a ({signal_3272, signal_1814}), .b ({signal_3625, signal_2167}), .clk ( clk ), .r ( Fresh[750] ), .c ({signal_3684, signal_2226}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2212 ( .a ({signal_3576, signal_2118}), .b ({signal_3626, signal_2168}), .clk ( clk ), .r ( Fresh[751] ), .c ({signal_3685, signal_2227}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2214 ( .a ({signal_3278, signal_1820}), .b ({signal_3627, signal_2169}), .clk ( clk ), .r ( Fresh[752] ), .c ({signal_3687, signal_2229}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2215 ( .a ({signal_3578, signal_2120}), .b ({signal_3628, signal_2170}), .clk ( clk ), .r ( Fresh[753] ), .c ({signal_3688, signal_2230}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2216 ( .a ({signal_2964, signal_1506}), .b ({signal_3629, signal_2171}), .clk ( clk ), .r ( Fresh[754] ), .c ({signal_3689, signal_2231}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2217 ( .a ({signal_3051, signal_1593}), .b ({signal_3631, signal_2173}), .clk ( clk ), .r ( Fresh[755] ), .c ({signal_3690, signal_2232}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2218 ( .a ({signal_3464, signal_2006}), .b ({signal_3633, signal_2175}), .clk ( clk ), .r ( Fresh[756] ), .c ({signal_3691, signal_2233}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2219 ( .a ({signal_2518, signal_1060}), .b ({signal_3634, signal_2176}), .clk ( clk ), .r ( Fresh[757] ), .c ({signal_3692, signal_2234}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2220 ( .a ({signal_2796, signal_1338}), .b ({signal_3636, signal_2178}), .clk ( clk ), .r ( Fresh[758] ), .c ({signal_3693, signal_2235}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2222 ( .a ({signal_3609, signal_2151}), .b ({signal_3585, signal_2127}), .clk ( clk ), .r ( Fresh[759] ), .c ({signal_3695, signal_2237}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2223 ( .a ({signal_3611, signal_2153}), .b ({signal_3640, signal_2182}), .clk ( clk ), .r ( Fresh[760] ), .c ({signal_3696, signal_2238}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2224 ( .a ({signal_2407, signal_949}), .b ({signal_3642, signal_2184}), .clk ( clk ), .r ( Fresh[761] ), .c ({signal_3697, signal_2239}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2239 ( .a ({signal_3681, signal_2223}), .b ({signal_3712, signal_2254}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2241 ( .a ({signal_3690, signal_2232}), .b ({signal_3714, signal_2256}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2243 ( .a ({signal_3697, signal_2239}), .b ({signal_3716, signal_2258}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2249 ( .a ({signal_3620, signal_2162}), .b ({signal_3659, signal_2201}), .clk ( clk ), .r ( Fresh[762] ), .c ({signal_3722, signal_2264}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2250 ( .a ({signal_3602, signal_2144}), .b ({signal_3661, signal_2203}), .clk ( clk ), .r ( Fresh[763] ), .c ({signal_3723, signal_2265}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2251 ( .a ({signal_2462, signal_1004}), .b ({signal_3662, signal_2204}), .clk ( clk ), .r ( Fresh[764] ), .c ({signal_3724, signal_2266}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2252 ( .a ({signal_2446, signal_988}), .b ({signal_3664, signal_2206}), .clk ( clk ), .r ( Fresh[765] ), .c ({signal_3725, signal_2267}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2253 ( .a ({signal_2442, signal_984}), .b ({signal_3665, signal_2207}), .clk ( clk ), .r ( Fresh[766] ), .c ({signal_3726, signal_2268}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2254 ( .a ({signal_2443, signal_985}), .b ({signal_3667, signal_2209}), .clk ( clk ), .r ( Fresh[767] ), .c ({signal_3727, signal_2269}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2271 ( .a ({signal_3724, signal_2266}), .b ({signal_3744, signal_2286}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2272 ( .a ({signal_3725, signal_2267}), .b ({signal_3745, signal_2287}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2273 ( .a ({signal_3726, signal_2268}), .b ({signal_3746, signal_2288}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2274 ( .a ({signal_3727, signal_2269}), .b ({signal_3747, signal_2289}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2282 ( .a ({signal_3708, signal_2250}), .b ({signal_3095, signal_1637}), .clk ( clk ), .r ( Fresh[768] ), .c ({signal_3755, signal_2297}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2283 ( .a ({signal_2442, signal_984}), .b ({signal_3706, signal_2248}), .clk ( clk ), .r ( Fresh[769] ), .c ({signal_3756, signal_2298}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2285 ( .a ({signal_2976, signal_1518}), .b ({signal_3721, signal_2263}), .clk ( clk ), .r ( Fresh[770] ), .c ({signal_3758, signal_2300}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2286 ( .a ({signal_3276, signal_1818}), .b ({signal_3709, signal_2251}), .clk ( clk ), .r ( Fresh[771] ), .c ({signal_3759, signal_2301}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2297 ( .a ({signal_3756, signal_2298}), .b ({signal_3770, signal_2312}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2180 ( .a ({signal_2712, signal_1254}), .b ({signal_3589, signal_2131}), .clk ( clk ), .r ( Fresh[772] ), .c ({signal_3653, signal_2195}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2181 ( .a ({signal_3446, signal_1988}), .b ({signal_3591, signal_2133}), .clk ( clk ), .r ( Fresh[773] ), .c ({signal_3654, signal_2196}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2182 ( .a ({signal_3077, signal_1619}), .b ({signal_3594, signal_2136}), .clk ( clk ), .r ( Fresh[774] ), .c ({signal_3655, signal_2197}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2183 ( .a ({signal_2808, signal_1350}), .b ({signal_3595, signal_2137}), .clk ( clk ), .r ( Fresh[775] ), .c ({signal_3656, signal_2198}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2199 ( .a ({signal_3653, signal_2195}), .b ({signal_3672, signal_2214}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2225 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_3643, signal_2185}), .clk ( clk ), .r ( Fresh[776] ), .c ({signal_3698, signal_2240}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2226 ( .a ({signal_3574, signal_2116}), .b ({signal_3645, signal_2187}), .clk ( clk ), .r ( Fresh[777] ), .c ({signal_3699, signal_2241}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2227 ( .a ({signal_2443, signal_985}), .b ({signal_3613, signal_2155}), .clk ( clk ), .r ( Fresh[778] ), .c ({signal_3700, signal_2242}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2228 ( .a ({signal_3650, signal_2192}), .b ({signal_3614, signal_2156}), .clk ( clk ), .r ( Fresh[779] ), .c ({signal_3701, signal_2243}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2229 ( .a ({signal_3567, signal_2109}), .b ({signal_3652, signal_2194}), .clk ( clk ), .r ( Fresh[780] ), .c ({signal_3702, signal_2244}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2244 ( .a ({signal_3698, signal_2240}), .b ({signal_3717, signal_2259}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2245 ( .a ({signal_3700, signal_2242}), .b ({signal_3718, signal_2260}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2246 ( .a ({signal_3702, signal_2244}), .b ({signal_3719, signal_2261}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2247 ( .a ({signal_2705, signal_1247}), .b ({signal_3673, signal_2215}), .clk ( clk ), .r ( Fresh[781] ), .c ({signal_3720, signal_2262}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2255 ( .a ({signal_3474, signal_2016}), .b ({signal_3682, signal_2224}), .clk ( clk ), .r ( Fresh[782] ), .c ({signal_3728, signal_2270}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2256 ( .a ({signal_3268, signal_1810}), .b ({signal_3683, signal_2225}), .clk ( clk ), .r ( Fresh[783] ), .c ({signal_3729, signal_2271}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2257 ( .a ({signal_3033, signal_1575}), .b ({signal_3684, signal_2226}), .clk ( clk ), .r ( Fresh[784] ), .c ({signal_3730, signal_2272}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2258 ( .a ({signal_3437, signal_1979}), .b ({signal_3685, signal_2227}), .clk ( clk ), .r ( Fresh[785] ), .c ({signal_3731, signal_2273}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2259 ( .a ({signal_3045, signal_1587}), .b ({signal_3687, signal_2229}), .clk ( clk ), .r ( Fresh[786] ), .c ({signal_3732, signal_2274}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2260 ( .a ({signal_3319, signal_1861}), .b ({signal_3688, signal_2230}), .clk ( clk ), .r ( Fresh[787] ), .c ({signal_3733, signal_2275}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2261 ( .a ({signal_2716, signal_1258}), .b ({signal_3689, signal_2231}), .clk ( clk ), .r ( Fresh[788] ), .c ({signal_3734, signal_2276}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2262 ( .a ({SI_s1[0], SI_s0[0]}), .b ({signal_3669, signal_2211}), .clk ( clk ), .r ( Fresh[789] ), .c ({signal_3735, signal_2277}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2263 ( .a ({signal_2524, signal_1066}), .b ({signal_3692, signal_2234}), .clk ( clk ), .r ( Fresh[790] ), .c ({signal_3736, signal_2278}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2264 ( .a ({signal_3663, signal_2205}), .b ({signal_3693, signal_2235}), .clk ( clk ), .r ( Fresh[791] ), .c ({signal_3737, signal_2279}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2265 ( .a ({signal_2450, signal_992}), .b ({signal_3670, signal_2212}), .clk ( clk ), .r ( Fresh[792] ), .c ({signal_3738, signal_2280}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2266 ( .a ({signal_3072, signal_1614}), .b ({signal_3695, signal_2237}), .clk ( clk ), .r ( Fresh[793] ), .c ({signal_3739, signal_2281}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2275 ( .a ({signal_3729, signal_2271}), .b ({signal_3748, signal_2290}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2276 ( .a ({signal_3730, signal_2272}), .b ({signal_3749, signal_2291}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2277 ( .a ({signal_3732, signal_2274}), .b ({signal_3750, signal_2292}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2278 ( .a ({signal_3734, signal_2276}), .b ({signal_3751, signal_2293}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2279 ( .a ({signal_3735, signal_2277}), .b ({signal_3752, signal_2294}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2280 ( .a ({signal_3738, signal_2280}), .b ({signal_3753, signal_2295}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2287 ( .a ({signal_3722, signal_2264}), .b ({signal_3680, signal_2222}), .clk ( clk ), .r ( Fresh[794] ), .c ({signal_3760, signal_2302}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2288 ( .a ({signal_2459, signal_1001}), .b ({signal_3712, signal_2254}), .clk ( clk ), .r ( Fresh[795] ), .c ({signal_3761, signal_2303}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2290 ( .a ({signal_2459, signal_1001}), .b ({signal_3714, signal_2256}), .clk ( clk ), .r ( Fresh[796] ), .c ({signal_3763, signal_2305}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2299 ( .a ({signal_3761, signal_2303}), .b ({signal_3772, signal_2314}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2301 ( .a ({signal_3763, signal_2305}), .b ({signal_3774, signal_2316}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2304 ( .a ({signal_3007, signal_1549}), .b ({signal_3755, signal_2297}), .clk ( clk ), .r ( Fresh[797] ), .c ({signal_3777, signal_2319}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2305 ( .a ({signal_3036, signal_1578}), .b ({signal_3758, signal_2300}), .clk ( clk ), .r ( Fresh[798] ), .c ({signal_3778, signal_2320}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2306 ( .a ({signal_3039, signal_1581}), .b ({signal_3759, signal_2301}), .clk ( clk ), .r ( Fresh[799] ), .c ({signal_3779, signal_2321}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2307 ( .a ({signal_3744, signal_2286}), .b ({signal_3691, signal_2233}), .clk ( clk ), .r ( Fresh[800] ), .c ({signal_3780, signal_2322}) ) ;

    /* cells in depth 17 */

    /* cells in depth 18 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2230 ( .a ({signal_3403, signal_1945}), .b ({signal_3654, signal_2196}), .clk ( clk ), .r ( Fresh[801] ), .c ({signal_3703, signal_2245}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2231 ( .a ({signal_3488, signal_2030}), .b ({signal_3655, signal_2197}), .clk ( clk ), .r ( Fresh[802] ), .c ({signal_3704, signal_2246}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2232 ( .a ({signal_3569, signal_2111}), .b ({signal_3656, signal_2198}), .clk ( clk ), .r ( Fresh[803] ), .c ({signal_3705, signal_2247}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2267 ( .a ({signal_3434, signal_1976}), .b ({signal_3699, signal_2241}), .clk ( clk ), .r ( Fresh[804] ), .c ({signal_3740, signal_2282}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2268 ( .a ({signal_2420, signal_962}), .b ({signal_3672, signal_2214}), .clk ( clk ), .r ( Fresh[805] ), .c ({signal_3741, signal_2283}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2281 ( .a ({signal_3741, signal_2283}), .b ({signal_3754, signal_2296}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2284 ( .a ({signal_2963, signal_1505}), .b ({signal_3720, signal_2262}), .clk ( clk ), .r ( Fresh[806] ), .c ({signal_3757, signal_2299}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2289 ( .a ({signal_3716, signal_2258}), .b ({signal_3717, signal_2259}), .clk ( clk ), .r ( Fresh[807] ), .c ({signal_3762, signal_2304}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2291 ( .a ({signal_3528, signal_2070}), .b ({signal_3728, signal_2270}), .clk ( clk ), .r ( Fresh[808] ), .c ({signal_3764, signal_2306}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2292 ( .a ({signal_3440, signal_1982}), .b ({signal_3731, signal_2273}), .clk ( clk ), .r ( Fresh[809] ), .c ({signal_3765, signal_2307}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2293 ( .a ({signal_3047, signal_1589}), .b ({signal_3733, signal_2275}), .clk ( clk ), .r ( Fresh[810] ), .c ({signal_3766, signal_2308}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2294 ( .a ({signal_3425, signal_1967}), .b ({signal_3736, signal_2278}), .clk ( clk ), .r ( Fresh[811] ), .c ({signal_3767, signal_2309}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2295 ( .a ({signal_3348, signal_1890}), .b ({signal_3719, signal_2261}), .clk ( clk ), .r ( Fresh[812] ), .c ({signal_3768, signal_2310}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2298 ( .a ({signal_3757, signal_2299}), .b ({signal_3771, signal_2313}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2300 ( .a ({signal_3762, signal_2304}), .b ({signal_3773, signal_2315}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2302 ( .a ({signal_3767, signal_2309}), .b ({signal_3775, signal_2317}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2303 ( .a ({signal_3768, signal_2310}), .b ({signal_3776, signal_2318}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2308 ( .a ({signal_3460, signal_2002}), .b ({signal_3748, signal_2290}), .clk ( clk ), .r ( Fresh[813] ), .c ({signal_3781, signal_2323}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2309 ( .a ({signal_2443, signal_985}), .b ({signal_3749, signal_2291}), .clk ( clk ), .r ( Fresh[814] ), .c ({signal_3782, signal_2324}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2310 ( .a ({signal_2443, signal_985}), .b ({signal_3750, signal_2292}), .clk ( clk ), .r ( Fresh[815] ), .c ({signal_3783, signal_2325}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2311 ( .a ({signal_2407, signal_949}), .b ({signal_3751, signal_2293}), .clk ( clk ), .r ( Fresh[816] ), .c ({signal_3784, signal_2326}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2312 ( .a ({signal_3711, signal_2253}), .b ({signal_3752, signal_2294}), .clk ( clk ), .r ( Fresh[817] ), .c ({signal_3785, signal_2327}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2313 ( .a ({signal_3760, signal_2302}), .b ({signal_3737, signal_2279}), .clk ( clk ), .r ( Fresh[818] ), .c ({signal_3786, signal_2328}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2314 ( .a ({signal_3564, signal_2106}), .b ({signal_3753, signal_2295}), .clk ( clk ), .r ( Fresh[819] ), .c ({signal_3787, signal_2329}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2315 ( .a ({signal_3745, signal_2287}), .b ({signal_3701, signal_2243}), .clk ( clk ), .r ( Fresh[820] ), .c ({signal_3788, signal_2330}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2320 ( .a ({signal_3781, signal_2323}), .b ({signal_3793, signal_2335}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2321 ( .a ({signal_3782, signal_2324}), .b ({signal_3794, signal_2336}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2322 ( .a ({signal_3783, signal_2325}), .b ({signal_3795, signal_2337}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2323 ( .a ({signal_3784, signal_2326}), .b ({signal_3796, signal_2338}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2324 ( .a ({signal_3526, signal_2068}), .b ({signal_3777, signal_2319}), .clk ( clk ), .r ( Fresh[821] ), .c ({signal_3797, signal_2339}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2326 ( .a ({signal_3666, signal_2208}), .b ({signal_3772, signal_2314}), .clk ( clk ), .r ( Fresh[822] ), .c ({signal_3799, signal_2341}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2328 ( .a ({signal_3531, signal_2073}), .b ({signal_3778, signal_2320}), .clk ( clk ), .r ( Fresh[823] ), .c ({signal_3801, signal_2343}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2329 ( .a ({signal_3770, signal_2312}), .b ({signal_3779, signal_2321}), .clk ( clk ), .r ( Fresh[824] ), .c ({signal_3802, signal_2344}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2330 ( .a ({signal_3707, signal_2249}), .b ({signal_3774, signal_2316}), .clk ( clk ), .r ( Fresh[825] ), .c ({signal_3803, signal_2345}) ) ;

    /* cells in depth 19 */

    /* cells in depth 20 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2269 ( .a ({signal_3619, signal_2161}), .b ({signal_3703, signal_2245}), .clk ( clk ), .r ( Fresh[826] ), .c ({signal_3742, signal_2284}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2270 ( .a ({signal_3568, signal_2110}), .b ({signal_3705, signal_2247}), .clk ( clk ), .r ( Fresh[827] ), .c ({signal_3743, signal_2285}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2296 ( .a ({signal_3657, signal_2199}), .b ({signal_3740, signal_2282}), .clk ( clk ), .r ( Fresh[828] ), .c ({signal_3769, signal_2311}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2316 ( .a ({signal_3436, signal_1978}), .b ({signal_3765, signal_2307}), .clk ( clk ), .r ( Fresh[829] ), .c ({signal_3789, signal_2331}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2317 ( .a ({signal_3713, signal_2255}), .b ({signal_3754, signal_2296}), .clk ( clk ), .r ( Fresh[830] ), .c ({signal_3790, signal_2332}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2318 ( .a ({signal_3746, signal_2288}), .b ({signal_3704, signal_2246}), .clk ( clk ), .r ( Fresh[831] ), .c ({signal_3791, signal_2333}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2325 ( .a ({signal_2439, signal_981}), .b ({signal_3771, signal_2313}), .clk ( clk ), .r ( Fresh[832] ), .c ({signal_3798, signal_2340}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2327 ( .a ({signal_3641, signal_2183}), .b ({signal_3773, signal_2315}), .clk ( clk ), .r ( Fresh[833] ), .c ({signal_3800, signal_2342}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2331 ( .a ({signal_3444, signal_1986}), .b ({signal_3785, signal_2327}), .clk ( clk ), .r ( Fresh[834] ), .c ({signal_3804, signal_2346}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2332 ( .a ({signal_2442, signal_984}), .b ({signal_3775, signal_2317}), .clk ( clk ), .r ( Fresh[835] ), .c ({signal_3805, signal_2347}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2333 ( .a ({signal_3540, signal_2082}), .b ({signal_3787, signal_2329}), .clk ( clk ), .r ( Fresh[836] ), .c ({signal_3806, signal_2348}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2335 ( .a ({signal_3798, signal_2340}), .b ({signal_3808, signal_2350}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2336 ( .a ({signal_3805, signal_2347}), .b ({signal_3809, signal_2351}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2337 ( .a ({signal_3671, signal_2213}), .b ({signal_3799, signal_2341}), .clk ( clk ), .r ( Fresh[837] ), .c ({signal_3810, signal_2352}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2339 ( .a ({signal_3710, signal_2252}), .b ({signal_3802, signal_2344}), .clk ( clk ), .r ( Fresh[838] ), .c ({signal_3812, signal_2354}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2340 ( .a ({signal_3618, signal_2160}), .b ({signal_3795, signal_2337}), .clk ( clk ), .r ( Fresh[839] ), .c ({signal_3813, signal_2355}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2341 ( .a ({signal_3647, signal_2189}), .b ({signal_3796, signal_2338}), .clk ( clk ), .r ( Fresh[840] ), .c ({signal_3814, signal_2356}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2342 ( .a ({signal_3596, signal_2138}), .b ({signal_3803, signal_2345}), .clk ( clk ), .r ( Fresh[841] ), .c ({signal_3815, signal_2357}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2343 ( .a ({signal_3797, signal_2339}), .b ({signal_3788, signal_2330}), .clk ( clk ), .r ( Fresh[842] ), .c ({signal_3816, signal_2358}) ) ;

    /* cells in depth 21 */

    /* cells in depth 22 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2319 ( .a ({signal_3660, signal_2202}), .b ({signal_3769, signal_2311}), .clk ( clk ), .r ( Fresh[843] ), .c ({signal_3792, signal_2334}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2334 ( .a ({signal_3194, signal_1736}), .b ({signal_3789, signal_2331}), .clk ( clk ), .r ( Fresh[844] ), .c ({signal_3807, signal_2349}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2338 ( .a ({signal_3696, signal_2238}), .b ({signal_3800, signal_2342}), .clk ( clk ), .r ( Fresh[845] ), .c ({signal_3811, signal_2353}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2344 ( .a ({signal_3804, signal_2346}), .b ({signal_3742, signal_2284}), .clk ( clk ), .r ( Fresh[846] ), .c ({signal_3817, signal_2359}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2346 ( .a ({signal_3668, signal_2210}), .b ({signal_3808, signal_2350}), .clk ( clk ), .r ( Fresh[847] ), .c ({signal_3819, signal_2361}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2348 ( .a ({signal_2985, signal_1527}), .b ({signal_3813, signal_2355}), .clk ( clk ), .r ( Fresh[848] ), .c ({signal_3821, signal_2363}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2349 ( .a ({signal_3612, signal_2154}), .b ({signal_3814, signal_2356}), .clk ( clk ), .r ( Fresh[849] ), .c ({signal_3822, signal_2364}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2350 ( .a ({signal_3091, signal_1633}), .b ({signal_3809, signal_2351}), .clk ( clk ), .r ( Fresh[850] ), .c ({signal_3823, signal_2365}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2351 ( .a ({signal_3607, signal_2149}), .b ({signal_3816, signal_2358}), .clk ( clk ), .r ( Fresh[851] ), .c ({signal_3824, signal_2366}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2352 ( .a ({signal_3810, signal_2352}), .b ({signal_3791, signal_2333}), .clk ( clk ), .r ( Fresh[852] ), .c ({signal_3825, signal_2367}) ) ;

    /* cells in depth 23 */

    /* cells in depth 24 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2345 ( .a ({signal_3793, signal_2335}), .b ({signal_3792, signal_2334}), .clk ( clk ), .r ( Fresh[853] ), .c ({signal_3818, signal_2360}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2347 ( .a ({signal_3610, signal_2152}), .b ({signal_3811, signal_2353}), .clk ( clk ), .r ( Fresh[854] ), .c ({signal_3820, signal_2362}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2353 ( .a ({signal_3812, signal_2354}), .b ({signal_3807, signal_2349}), .clk ( clk ), .r ( Fresh[855] ), .c ({signal_3826, signal_2368}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2354 ( .a ({signal_3815, signal_2357}), .b ({signal_3817, signal_2359}), .clk ( clk ), .r ( Fresh[856] ), .c ({signal_3827, signal_2369}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2357 ( .a ({signal_3046, signal_1588}), .b ({signal_3821, signal_2363}), .clk ( clk ), .r ( Fresh[857] ), .c ({signal_3830, signal_2372}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2358 ( .a ({signal_3766, signal_2308}), .b ({signal_3822, signal_2364}), .clk ( clk ), .r ( Fresh[858] ), .c ({signal_3831, signal_2373}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2359 ( .a ({signal_3060, signal_1602}), .b ({signal_3823, signal_2365}), .clk ( clk ), .r ( Fresh[859] ), .c ({signal_3832, signal_2374}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2360 ( .a ({signal_3715, signal_2257}), .b ({signal_3824, signal_2366}), .clk ( clk ), .r ( Fresh[860] ), .c ({signal_3833, signal_2375}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2361 ( .a ({signal_3776, signal_2318}), .b ({signal_3825, signal_2367}), .clk ( clk ), .r ( Fresh[861] ), .c ({signal_3834, signal_2376}) ) ;

    /* cells in depth 25 */

    /* cells in depth 26 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2355 ( .a ({signal_3794, signal_2336}), .b ({signal_3818, signal_2360}), .clk ( clk ), .r ( Fresh[862] ), .c ({signal_3828, signal_2370}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2356 ( .a ({signal_3747, signal_2289}), .b ({signal_3820, signal_2362}), .clk ( clk ), .r ( Fresh[863] ), .c ({signal_3829, signal_2371}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2362 ( .a ({signal_3801, signal_2343}), .b ({signal_3826, signal_2368}), .clk ( clk ), .r ( Fresh[864] ), .c ({signal_3835, signal_2377}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2363 ( .a ({signal_3723, signal_2265}), .b ({signal_3827, signal_2369}), .clk ( clk ), .r ( Fresh[865] ), .c ({signal_3836, signal_2378}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2365 ( .a ({signal_3836, signal_2378}), .b ({signal_3838, signal_26}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2368 ( .a ({signal_3241, signal_1783}), .b ({signal_3830, signal_2372}), .clk ( clk ), .r ( Fresh[866] ), .c ({signal_3841, signal_2381}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2369 ( .a ({signal_2997, signal_1539}), .b ({signal_3832, signal_2374}), .clk ( clk ), .r ( Fresh[867] ), .c ({signal_3842, signal_2382}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2370 ( .a ({signal_3806, signal_2348}), .b ({signal_3833, signal_2375}), .clk ( clk ), .r ( Fresh[868] ), .c ({signal_3843, signal_2383}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2371 ( .a ({signal_3739, signal_2281}), .b ({signal_3834, signal_2376}), .clk ( clk ), .r ( Fresh[869] ), .c ({signal_3844, signal_2384}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2374 ( .a ({signal_3843, signal_2383}), .b ({signal_3847, signal_28}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2375 ( .a ({signal_3844, signal_2384}), .b ({signal_3848, signal_29}) ) ;

    /* cells in depth 27 */

    /* cells in depth 28 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2364 ( .a ({signal_3764, signal_2306}), .b ({signal_3828, signal_2370}), .clk ( clk ), .r ( Fresh[870] ), .c ({signal_3837, signal_2379}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2366 ( .a ({signal_3837, signal_2379}), .b ({signal_3839, signal_23}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2367 ( .a ({signal_3743, signal_2285}), .b ({signal_3829, signal_2371}), .clk ( clk ), .r ( Fresh[871] ), .c ({signal_3840, signal_2380}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2372 ( .a ({signal_3819, signal_2361}), .b ({signal_3835, signal_2377}), .clk ( clk ), .r ( Fresh[872] ), .c ({signal_3845, signal_2385}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2373 ( .a ({signal_3840, signal_2380}), .b ({signal_3846, signal_30}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2376 ( .a ({signal_3845, signal_2385}), .b ({signal_3849, signal_24}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2377 ( .a ({signal_3831, signal_2373}), .b ({signal_3841, signal_2381}), .clk ( clk ), .r ( Fresh[873] ), .c ({signal_3850, signal_2386}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2378 ( .a ({signal_3061, signal_1603}), .b ({signal_3842, signal_2382}), .clk ( clk ), .r ( Fresh[874] ), .c ({signal_3851, signal_2387}) ) ;

    /* cells in depth 29 */

    /* cells in depth 30 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2379 ( .a ({signal_3790, signal_2332}), .b ({signal_3850, signal_2386}), .clk ( clk ), .r ( Fresh[875] ), .c ({signal_3852, signal_2388}) ) ;
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2380 ( .a ({signal_3718, signal_2260}), .b ({signal_3851, signal_2387}), .clk ( clk ), .r ( Fresh[876] ), .c ({signal_3853, signal_2389}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2381 ( .a ({signal_3852, signal_2388}), .b ({signal_3854, signal_25}) ) ;

    /* cells in depth 31 */

    /* cells in depth 32 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2382 ( .a ({signal_3780, signal_2322}), .b ({signal_3853, signal_2389}), .clk ( clk ), .r ( Fresh[877] ), .c ({signal_3855, signal_2390}) ) ;

    /* cells in depth 33 */

    /* cells in depth 34 */
    and_HPC2 #(.security_order(1), .pipeline(0)) cell_2383 ( .a ({signal_3786, signal_2328}), .b ({signal_3855, signal_2390}), .clk ( clk ), .r ( Fresh[878] ), .c ({signal_3856, signal_2391}) ) ;
    not_masked #(.security_order(1), .pipeline(0)) cell_2384 ( .a ({signal_3856, signal_2391}), .b ({signal_3857, signal_27}) ) ;

    /* register cells */
    reg_masked #(.security_order(1), .pipeline(0)) cell_0 ( .clk ( signal_4746 ), .D ({signal_3839, signal_23}), .Q ({SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_1 ( .clk ( signal_4746 ), .D ({signal_3849, signal_24}), .Q ({SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_2 ( .clk ( signal_4746 ), .D ({signal_3854, signal_25}), .Q ({SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_3 ( .clk ( signal_4746 ), .D ({signal_3838, signal_26}), .Q ({SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_4 ( .clk ( signal_4746 ), .D ({signal_3857, signal_27}), .Q ({SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_5 ( .clk ( signal_4746 ), .D ({signal_3847, signal_28}), .Q ({SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_6 ( .clk ( signal_4746 ), .D ({signal_3848, signal_29}), .Q ({SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.security_order(1), .pipeline(0)) cell_7 ( .clk ( signal_4746 ), .D ({signal_3846, signal_30}), .Q ({SO_s1[0], SO_s0[0]}) ) ;
endmodule
