/* modified netlist. Source: module AES in file ../CaseStudies/07_AES128_byte_serial_encryption/netlists/AES.v */
/* 0 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 1 register stage(s) in total */

module AES_LMDPL_Pipeline_d1 (plaintext_s0, key_s0, clk, start, Po_rst, Fresh, plaintext_s1, key_s1, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input start ;
    input Po_rst ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [33:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire nReset ;
    wire selMC ;
    wire selSR ;
    wire selXOR ;
    wire enRCon ;
    wire finalStep ;
    wire intFinal ;
    wire intselXOR ;
    wire notFirst ;
    wire n10 ;
    wire n9 ;
    wire n12 ;
    wire n13 ;
    wire ctrl_n16 ;
    wire ctrl_n15 ;
    wire ctrl_n14 ;
    wire ctrl_n11 ;
    wire ctrl_n10 ;
    wire ctrl_n9 ;
    wire ctrl_n8 ;
    wire ctrl_n7 ;
    wire ctrl_n5 ;
    wire ctrl_n4 ;
    wire ctrl_n2 ;
    wire ctrl_n12 ;
    wire ctrl_n6 ;
    wire ctrl_N14 ;
    wire ctrl_seq4Out_1_ ;
    wire ctrl_seq4In_1_ ;
    wire ctrl_nRstSeq4 ;
    wire ctrl_n13 ;
    wire ctrl_seq6Out_4_ ;
    wire ctrl_seq6In_1_ ;
    wire ctrl_seq6In_2_ ;
    wire ctrl_seq6In_3_ ;
    wire ctrl_seq6In_4_ ;
    wire ctrl_seq6_SFF_0_QD ;
    wire ctrl_seq6_SFF_1_QD ;
    wire ctrl_seq6_SFF_2_QD ;
    wire ctrl_seq6_SFF_3_QD ;
    wire ctrl_seq6_SFF_4_QD ;
    wire ctrl_seq4_SFF_0_QD ;
    wire ctrl_seq4_SFF_1_QD ;
    wire stateArray_n33 ;
    wire stateArray_n32 ;
    wire stateArray_n31 ;
    wire stateArray_n30 ;
    wire stateArray_n29 ;
    wire stateArray_n28 ;
    wire stateArray_n27 ;
    wire stateArray_n26 ;
    wire stateArray_n25 ;
    wire stateArray_n24 ;
    wire stateArray_n23 ;
    wire stateArray_n22 ;
    wire stateArray_n21 ;
    wire stateArray_n20 ;
    wire stateArray_n19 ;
    wire stateArray_n18 ;
    wire stateArray_n17 ;
    wire stateArray_n16 ;
    wire stateArray_n15 ;
    wire stateArray_n14 ;
    wire stateArray_n13 ;
    wire stateArray_S00reg_gff_1_SFF_0_QD ;
    wire stateArray_S00reg_gff_1_SFF_1_QD ;
    wire stateArray_S00reg_gff_1_SFF_2_QD ;
    wire stateArray_S00reg_gff_1_SFF_3_QD ;
    wire stateArray_S00reg_gff_1_SFF_4_QD ;
    wire stateArray_S00reg_gff_1_SFF_5_QD ;
    wire stateArray_S00reg_gff_1_SFF_6_QD ;
    wire stateArray_S00reg_gff_1_SFF_7_QD ;
    wire stateArray_S01reg_gff_1_SFF_0_QD ;
    wire stateArray_S01reg_gff_1_SFF_1_QD ;
    wire stateArray_S01reg_gff_1_SFF_2_QD ;
    wire stateArray_S01reg_gff_1_SFF_3_QD ;
    wire stateArray_S01reg_gff_1_SFF_4_QD ;
    wire stateArray_S01reg_gff_1_SFF_5_QD ;
    wire stateArray_S01reg_gff_1_SFF_6_QD ;
    wire stateArray_S01reg_gff_1_SFF_7_QD ;
    wire stateArray_S02reg_gff_1_SFF_0_QD ;
    wire stateArray_S02reg_gff_1_SFF_1_QD ;
    wire stateArray_S02reg_gff_1_SFF_2_QD ;
    wire stateArray_S02reg_gff_1_SFF_3_QD ;
    wire stateArray_S02reg_gff_1_SFF_4_QD ;
    wire stateArray_S02reg_gff_1_SFF_5_QD ;
    wire stateArray_S02reg_gff_1_SFF_6_QD ;
    wire stateArray_S02reg_gff_1_SFF_7_QD ;
    wire stateArray_S03reg_gff_1_SFF_0_QD ;
    wire stateArray_S03reg_gff_1_SFF_1_QD ;
    wire stateArray_S03reg_gff_1_SFF_2_QD ;
    wire stateArray_S03reg_gff_1_SFF_3_QD ;
    wire stateArray_S03reg_gff_1_SFF_4_QD ;
    wire stateArray_S03reg_gff_1_SFF_5_QD ;
    wire stateArray_S03reg_gff_1_SFF_6_QD ;
    wire stateArray_S03reg_gff_1_SFF_7_QD ;
    wire stateArray_S10reg_gff_1_SFF_0_QD ;
    wire stateArray_S10reg_gff_1_SFF_1_QD ;
    wire stateArray_S10reg_gff_1_SFF_2_QD ;
    wire stateArray_S10reg_gff_1_SFF_3_QD ;
    wire stateArray_S10reg_gff_1_SFF_4_QD ;
    wire stateArray_S10reg_gff_1_SFF_5_QD ;
    wire stateArray_S10reg_gff_1_SFF_6_QD ;
    wire stateArray_S10reg_gff_1_SFF_7_QD ;
    wire stateArray_S11reg_gff_1_SFF_0_QD ;
    wire stateArray_S11reg_gff_1_SFF_1_QD ;
    wire stateArray_S11reg_gff_1_SFF_2_QD ;
    wire stateArray_S11reg_gff_1_SFF_3_QD ;
    wire stateArray_S11reg_gff_1_SFF_4_QD ;
    wire stateArray_S11reg_gff_1_SFF_5_QD ;
    wire stateArray_S11reg_gff_1_SFF_6_QD ;
    wire stateArray_S11reg_gff_1_SFF_7_QD ;
    wire stateArray_S12reg_gff_1_SFF_0_QD ;
    wire stateArray_S12reg_gff_1_SFF_1_QD ;
    wire stateArray_S12reg_gff_1_SFF_2_QD ;
    wire stateArray_S12reg_gff_1_SFF_3_QD ;
    wire stateArray_S12reg_gff_1_SFF_4_QD ;
    wire stateArray_S12reg_gff_1_SFF_5_QD ;
    wire stateArray_S12reg_gff_1_SFF_6_QD ;
    wire stateArray_S12reg_gff_1_SFF_7_QD ;
    wire stateArray_S13reg_gff_1_SFF_0_QD ;
    wire stateArray_S13reg_gff_1_SFF_1_QD ;
    wire stateArray_S13reg_gff_1_SFF_2_QD ;
    wire stateArray_S13reg_gff_1_SFF_3_QD ;
    wire stateArray_S13reg_gff_1_SFF_4_QD ;
    wire stateArray_S13reg_gff_1_SFF_5_QD ;
    wire stateArray_S13reg_gff_1_SFF_6_QD ;
    wire stateArray_S13reg_gff_1_SFF_7_QD ;
    wire stateArray_S20reg_gff_1_SFF_0_QD ;
    wire stateArray_S20reg_gff_1_SFF_1_QD ;
    wire stateArray_S20reg_gff_1_SFF_2_QD ;
    wire stateArray_S20reg_gff_1_SFF_3_QD ;
    wire stateArray_S20reg_gff_1_SFF_4_QD ;
    wire stateArray_S20reg_gff_1_SFF_5_QD ;
    wire stateArray_S20reg_gff_1_SFF_6_QD ;
    wire stateArray_S20reg_gff_1_SFF_7_QD ;
    wire stateArray_S21reg_gff_1_SFF_0_QD ;
    wire stateArray_S21reg_gff_1_SFF_1_QD ;
    wire stateArray_S21reg_gff_1_SFF_2_QD ;
    wire stateArray_S21reg_gff_1_SFF_3_QD ;
    wire stateArray_S21reg_gff_1_SFF_4_QD ;
    wire stateArray_S21reg_gff_1_SFF_5_QD ;
    wire stateArray_S21reg_gff_1_SFF_6_QD ;
    wire stateArray_S21reg_gff_1_SFF_7_QD ;
    wire stateArray_S22reg_gff_1_SFF_0_QD ;
    wire stateArray_S22reg_gff_1_SFF_1_QD ;
    wire stateArray_S22reg_gff_1_SFF_2_QD ;
    wire stateArray_S22reg_gff_1_SFF_3_QD ;
    wire stateArray_S22reg_gff_1_SFF_4_QD ;
    wire stateArray_S22reg_gff_1_SFF_5_QD ;
    wire stateArray_S22reg_gff_1_SFF_6_QD ;
    wire stateArray_S22reg_gff_1_SFF_7_QD ;
    wire stateArray_S23reg_gff_1_SFF_0_QD ;
    wire stateArray_S23reg_gff_1_SFF_1_QD ;
    wire stateArray_S23reg_gff_1_SFF_2_QD ;
    wire stateArray_S23reg_gff_1_SFF_3_QD ;
    wire stateArray_S23reg_gff_1_SFF_4_QD ;
    wire stateArray_S23reg_gff_1_SFF_5_QD ;
    wire stateArray_S23reg_gff_1_SFF_6_QD ;
    wire stateArray_S23reg_gff_1_SFF_7_QD ;
    wire stateArray_S30reg_gff_1_SFF_0_QD ;
    wire stateArray_S30reg_gff_1_SFF_1_QD ;
    wire stateArray_S30reg_gff_1_SFF_2_QD ;
    wire stateArray_S30reg_gff_1_SFF_3_QD ;
    wire stateArray_S30reg_gff_1_SFF_4_QD ;
    wire stateArray_S30reg_gff_1_SFF_5_QD ;
    wire stateArray_S30reg_gff_1_SFF_6_QD ;
    wire stateArray_S30reg_gff_1_SFF_7_QD ;
    wire stateArray_S31reg_gff_1_SFF_0_QD ;
    wire stateArray_S31reg_gff_1_SFF_1_QD ;
    wire stateArray_S31reg_gff_1_SFF_2_QD ;
    wire stateArray_S31reg_gff_1_SFF_3_QD ;
    wire stateArray_S31reg_gff_1_SFF_4_QD ;
    wire stateArray_S31reg_gff_1_SFF_5_QD ;
    wire stateArray_S31reg_gff_1_SFF_6_QD ;
    wire stateArray_S31reg_gff_1_SFF_7_QD ;
    wire stateArray_S32reg_gff_1_SFF_0_QD ;
    wire stateArray_S32reg_gff_1_SFF_1_QD ;
    wire stateArray_S32reg_gff_1_SFF_2_QD ;
    wire stateArray_S32reg_gff_1_SFF_3_QD ;
    wire stateArray_S32reg_gff_1_SFF_4_QD ;
    wire stateArray_S32reg_gff_1_SFF_5_QD ;
    wire stateArray_S32reg_gff_1_SFF_6_QD ;
    wire stateArray_S32reg_gff_1_SFF_7_QD ;
    wire stateArray_S33reg_gff_1_SFF_0_QD ;
    wire stateArray_S33reg_gff_1_SFF_1_QD ;
    wire stateArray_S33reg_gff_1_SFF_2_QD ;
    wire stateArray_S33reg_gff_1_SFF_3_QD ;
    wire stateArray_S33reg_gff_1_SFF_4_QD ;
    wire stateArray_S33reg_gff_1_SFF_5_QD ;
    wire stateArray_S33reg_gff_1_SFF_6_QD ;
    wire stateArray_S33reg_gff_1_SFF_7_QD ;
    wire MUX_StateInMC_n7 ;
    wire MUX_StateInMC_n6 ;
    wire MUX_StateInMC_n5 ;
    wire KeyArray_n55 ;
    wire KeyArray_n54 ;
    wire KeyArray_n53 ;
    wire KeyArray_n52 ;
    wire KeyArray_n51 ;
    wire KeyArray_n50 ;
    wire KeyArray_n49 ;
    wire KeyArray_n48 ;
    wire KeyArray_n47 ;
    wire KeyArray_n46 ;
    wire KeyArray_n45 ;
    wire KeyArray_n44 ;
    wire KeyArray_n43 ;
    wire KeyArray_n42 ;
    wire KeyArray_n41 ;
    wire KeyArray_n40 ;
    wire KeyArray_n39 ;
    wire KeyArray_n38 ;
    wire KeyArray_n37 ;
    wire KeyArray_n36 ;
    wire KeyArray_n35 ;
    wire KeyArray_n34 ;
    wire KeyArray_n33 ;
    wire KeyArray_n32 ;
    wire KeyArray_n31 ;
    wire KeyArray_n30 ;
    wire KeyArray_n29 ;
    wire KeyArray_n28 ;
    wire KeyArray_n27 ;
    wire KeyArray_n26 ;
    wire KeyArray_n25 ;
    wire KeyArray_n24 ;
    wire KeyArray_n23 ;
    wire KeyArray_n22 ;
    wire KeyArray_outS01ser_0_ ;
    wire KeyArray_outS01ser_1_ ;
    wire KeyArray_outS01ser_2_ ;
    wire KeyArray_outS01ser_3_ ;
    wire KeyArray_outS01ser_4_ ;
    wire KeyArray_outS01ser_5_ ;
    wire KeyArray_outS01ser_6_ ;
    wire KeyArray_outS01ser_7_ ;
    wire KeyArray_S00reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S00reg_gff_1_SFF_0_QD ;
    wire KeyArray_S00reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_1_QD ;
    wire KeyArray_S00reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_2_QD ;
    wire KeyArray_S00reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_3_QD ;
    wire KeyArray_S00reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_4_QD ;
    wire KeyArray_S00reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_5_QD ;
    wire KeyArray_S00reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_6_QD ;
    wire KeyArray_S00reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S00reg_gff_1_SFF_7_QD ;
    wire KeyArray_S01reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_0_QD ;
    wire KeyArray_S01reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_1_QD ;
    wire KeyArray_S01reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_2_QD ;
    wire KeyArray_S01reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_3_QD ;
    wire KeyArray_S01reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_4_QD ;
    wire KeyArray_S01reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_5_QD ;
    wire KeyArray_S01reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_6_QD ;
    wire KeyArray_S01reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S01reg_gff_1_SFF_7_QD ;
    wire KeyArray_S02reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_0_QD ;
    wire KeyArray_S02reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_1_QD ;
    wire KeyArray_S02reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_2_QD ;
    wire KeyArray_S02reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_3_QD ;
    wire KeyArray_S02reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_4_QD ;
    wire KeyArray_S02reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_5_QD ;
    wire KeyArray_S02reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_6_QD ;
    wire KeyArray_S02reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S02reg_gff_1_SFF_7_QD ;
    wire KeyArray_S03reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_0_QD ;
    wire KeyArray_S03reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_1_QD ;
    wire KeyArray_S03reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_2_QD ;
    wire KeyArray_S03reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_3_QD ;
    wire KeyArray_S03reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S03reg_gff_1_SFF_4_QD ;
    wire KeyArray_S03reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_5_QD ;
    wire KeyArray_S03reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_6_QD ;
    wire KeyArray_S03reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S03reg_gff_1_SFF_7_QD ;
    wire KeyArray_S10reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_0_QD ;
    wire KeyArray_S10reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_1_QD ;
    wire KeyArray_S10reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_2_QD ;
    wire KeyArray_S10reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_3_QD ;
    wire KeyArray_S10reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_4_QD ;
    wire KeyArray_S10reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_5_QD ;
    wire KeyArray_S10reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_6_QD ;
    wire KeyArray_S10reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S10reg_gff_1_SFF_7_QD ;
    wire KeyArray_S11reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_0_QD ;
    wire KeyArray_S11reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_1_QD ;
    wire KeyArray_S11reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_2_QD ;
    wire KeyArray_S11reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_3_QD ;
    wire KeyArray_S11reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_4_QD ;
    wire KeyArray_S11reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_5_QD ;
    wire KeyArray_S11reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_6_QD ;
    wire KeyArray_S11reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S11reg_gff_1_SFF_7_QD ;
    wire KeyArray_S12reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_0_QD ;
    wire KeyArray_S12reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_1_QD ;
    wire KeyArray_S12reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_2_QD ;
    wire KeyArray_S12reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_3_QD ;
    wire KeyArray_S12reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_4_QD ;
    wire KeyArray_S12reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_5_QD ;
    wire KeyArray_S12reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_6_QD ;
    wire KeyArray_S12reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S12reg_gff_1_SFF_7_QD ;
    wire KeyArray_S13reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_0_QD ;
    wire KeyArray_S13reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_1_QD ;
    wire KeyArray_S13reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_2_QD ;
    wire KeyArray_S13reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_3_QD ;
    wire KeyArray_S13reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S13reg_gff_1_SFF_4_QD ;
    wire KeyArray_S13reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_5_QD ;
    wire KeyArray_S13reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_6_QD ;
    wire KeyArray_S13reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S13reg_gff_1_SFF_7_QD ;
    wire KeyArray_S20reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_0_QD ;
    wire KeyArray_S20reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_1_QD ;
    wire KeyArray_S20reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_2_QD ;
    wire KeyArray_S20reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_3_QD ;
    wire KeyArray_S20reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_4_QD ;
    wire KeyArray_S20reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_5_QD ;
    wire KeyArray_S20reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_6_QD ;
    wire KeyArray_S20reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S20reg_gff_1_SFF_7_QD ;
    wire KeyArray_S21reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_0_QD ;
    wire KeyArray_S21reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_1_QD ;
    wire KeyArray_S21reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_2_QD ;
    wire KeyArray_S21reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_3_QD ;
    wire KeyArray_S21reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_4_QD ;
    wire KeyArray_S21reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_5_QD ;
    wire KeyArray_S21reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_6_QD ;
    wire KeyArray_S21reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S21reg_gff_1_SFF_7_QD ;
    wire KeyArray_S22reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_0_QD ;
    wire KeyArray_S22reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_1_QD ;
    wire KeyArray_S22reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_2_QD ;
    wire KeyArray_S22reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_3_QD ;
    wire KeyArray_S22reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_4_QD ;
    wire KeyArray_S22reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_5_QD ;
    wire KeyArray_S22reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_6_QD ;
    wire KeyArray_S22reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S22reg_gff_1_SFF_7_QD ;
    wire KeyArray_S23reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_0_QD ;
    wire KeyArray_S23reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_1_QD ;
    wire KeyArray_S23reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_2_QD ;
    wire KeyArray_S23reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_3_QD ;
    wire KeyArray_S23reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S23reg_gff_1_SFF_4_QD ;
    wire KeyArray_S23reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_5_QD ;
    wire KeyArray_S23reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_6_QD ;
    wire KeyArray_S23reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S23reg_gff_1_SFF_7_QD ;
    wire KeyArray_S30reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_0_QD ;
    wire KeyArray_S30reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_1_QD ;
    wire KeyArray_S30reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_2_QD ;
    wire KeyArray_S30reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_3_QD ;
    wire KeyArray_S30reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_4_QD ;
    wire KeyArray_S30reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_5_QD ;
    wire KeyArray_S30reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_6_QD ;
    wire KeyArray_S30reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S30reg_gff_1_SFF_7_QD ;
    wire KeyArray_S31reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_0_QD ;
    wire KeyArray_S31reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_1_QD ;
    wire KeyArray_S31reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_2_QD ;
    wire KeyArray_S31reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_3_QD ;
    wire KeyArray_S31reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_4_QD ;
    wire KeyArray_S31reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_5_QD ;
    wire KeyArray_S31reg_gff_1_SFF_6_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_6_QD ;
    wire KeyArray_S31reg_gff_1_SFF_7_n6 ;
    wire KeyArray_S31reg_gff_1_SFF_7_QD ;
    wire KeyArray_S32reg_gff_1_SFF_0_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_0_QD ;
    wire KeyArray_S32reg_gff_1_SFF_1_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_1_QD ;
    wire KeyArray_S32reg_gff_1_SFF_2_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_2_QD ;
    wire KeyArray_S32reg_gff_1_SFF_3_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_3_QD ;
    wire KeyArray_S32reg_gff_1_SFF_4_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_4_QD ;
    wire KeyArray_S32reg_gff_1_SFF_5_n6 ;
    wire KeyArray_S32reg_gff_1_SFF_5_QD ;
    wire KeyArray_S32reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S32reg_gff_1_SFF_6_QD ;
    wire KeyArray_S32reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S32reg_gff_1_SFF_7_QD ;
    wire KeyArray_S33reg_gff_1_SFF_0_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_0_QD ;
    wire KeyArray_S33reg_gff_1_SFF_1_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_1_QD ;
    wire KeyArray_S33reg_gff_1_SFF_2_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_2_QD ;
    wire KeyArray_S33reg_gff_1_SFF_3_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_3_QD ;
    wire KeyArray_S33reg_gff_1_SFF_4_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_4_QD ;
    wire KeyArray_S33reg_gff_1_SFF_5_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_5_QD ;
    wire KeyArray_S33reg_gff_1_SFF_6_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_6_QD ;
    wire KeyArray_S33reg_gff_1_SFF_7_n5 ;
    wire KeyArray_S33reg_gff_1_SFF_7_QD ;
    wire MixColumns_line0_n16 ;
    wire MixColumns_line0_n15 ;
    wire MixColumns_line0_n14 ;
    wire MixColumns_line0_n13 ;
    wire MixColumns_line0_n12 ;
    wire MixColumns_line0_n11 ;
    wire MixColumns_line0_n10 ;
    wire MixColumns_line0_n9 ;
    wire MixColumns_line0_n8 ;
    wire MixColumns_line0_n7 ;
    wire MixColumns_line0_n6 ;
    wire MixColumns_line0_n5 ;
    wire MixColumns_line0_n4 ;
    wire MixColumns_line0_n3 ;
    wire MixColumns_line0_n2 ;
    wire MixColumns_line0_n1 ;
    wire MixColumns_line1_n16 ;
    wire MixColumns_line1_n15 ;
    wire MixColumns_line1_n14 ;
    wire MixColumns_line1_n13 ;
    wire MixColumns_line1_n12 ;
    wire MixColumns_line1_n11 ;
    wire MixColumns_line1_n10 ;
    wire MixColumns_line1_n9 ;
    wire MixColumns_line1_n8 ;
    wire MixColumns_line1_n7 ;
    wire MixColumns_line1_n6 ;
    wire MixColumns_line1_n5 ;
    wire MixColumns_line1_n4 ;
    wire MixColumns_line1_n3 ;
    wire MixColumns_line1_n2 ;
    wire MixColumns_line1_n1 ;
    wire MixColumns_line1_S02_1_ ;
    wire MixColumns_line1_S02_3_ ;
    wire MixColumns_line1_S02_4_ ;
    wire MixColumns_line2_n16 ;
    wire MixColumns_line2_n15 ;
    wire MixColumns_line2_n14 ;
    wire MixColumns_line2_n13 ;
    wire MixColumns_line2_n12 ;
    wire MixColumns_line2_n11 ;
    wire MixColumns_line2_n10 ;
    wire MixColumns_line2_n9 ;
    wire MixColumns_line2_n8 ;
    wire MixColumns_line2_n7 ;
    wire MixColumns_line2_n6 ;
    wire MixColumns_line2_n5 ;
    wire MixColumns_line2_n4 ;
    wire MixColumns_line2_n3 ;
    wire MixColumns_line2_n2 ;
    wire MixColumns_line2_n1 ;
    wire MixColumns_line2_S02_1_ ;
    wire MixColumns_line2_S02_3_ ;
    wire MixColumns_line2_S02_4_ ;
    wire MixColumns_line3_n16 ;
    wire MixColumns_line3_n15 ;
    wire MixColumns_line3_n14 ;
    wire MixColumns_line3_n13 ;
    wire MixColumns_line3_n12 ;
    wire MixColumns_line3_n11 ;
    wire MixColumns_line3_n10 ;
    wire MixColumns_line3_n9 ;
    wire MixColumns_line3_n8 ;
    wire MixColumns_line3_n7 ;
    wire MixColumns_line3_n6 ;
    wire MixColumns_line3_n5 ;
    wire MixColumns_line3_n4 ;
    wire MixColumns_line3_n3 ;
    wire MixColumns_line3_n2 ;
    wire MixColumns_line3_n1 ;
    wire MixColumns_line3_S02_1_ ;
    wire MixColumns_line3_S02_3_ ;
    wire MixColumns_line3_S02_4_ ;
    wire MixColumns_line3_timesTHREE_input2_1_ ;
    wire MixColumns_line3_timesTHREE_input2_3_ ;
    wire MixColumns_line3_timesTHREE_input2_4_ ;
    wire calcRCon_n38 ;
    wire calcRCon_n37 ;
    wire calcRCon_n36 ;
    wire calcRCon_n35 ;
    wire calcRCon_n34 ;
    wire calcRCon_n33 ;
    wire calcRCon_n32 ;
    wire calcRCon_n31 ;
    wire calcRCon_n30 ;
    wire calcRCon_n29 ;
    wire calcRCon_n28 ;
    wire calcRCon_n27 ;
    wire calcRCon_n26 ;
    wire calcRCon_n25 ;
    wire calcRCon_n24 ;
    wire calcRCon_n23 ;
    wire calcRCon_n22 ;
    wire calcRCon_n21 ;
    wire calcRCon_n20 ;
    wire calcRCon_n19 ;
    wire calcRCon_n18 ;
    wire calcRCon_n17 ;
    wire calcRCon_n10 ;
    wire calcRCon_n9 ;
    wire calcRCon_n8 ;
    wire calcRCon_n7 ;
    wire calcRCon_n6 ;
    wire calcRCon_n5 ;
    wire calcRCon_n3 ;
    wire calcRCon_n11 ;
    wire calcRCon_n44 ;
    wire calcRCon_n16 ;
    wire calcRCon_n45 ;
    wire calcRCon_n46 ;
    wire calcRCon_n47 ;
    wire calcRCon_n15 ;
    wire calcRCon_n48 ;
    wire calcRCon_n12 ;
    wire calcRCon_n49 ;
    wire calcRCon_n14 ;
    wire calcRCon_n50 ;
    wire calcRCon_n13 ;
    wire calcRCon_s_current_state_0_ ;
    wire calcRCon_s_current_state_1_ ;
    wire calcRCon_s_current_state_2_ ;
    wire calcRCon_s_current_state_3_ ;
    wire calcRCon_s_current_state_4_ ;
    wire calcRCon_s_current_state_5_ ;
    wire calcRCon_s_current_state_6_ ;
    wire calcRCon_n51 ;
    wire Inst_bSbox_L29 ;
    wire Inst_bSbox_L28 ;
    wire Inst_bSbox_L27 ;
    wire Inst_bSbox_L26 ;
    wire Inst_bSbox_L25 ;
    wire Inst_bSbox_L24 ;
    wire Inst_bSbox_L23 ;
    wire Inst_bSbox_L22 ;
    wire Inst_bSbox_L21 ;
    wire Inst_bSbox_L20 ;
    wire Inst_bSbox_L19 ;
    wire Inst_bSbox_L18 ;
    wire Inst_bSbox_L17 ;
    wire Inst_bSbox_L16 ;
    wire Inst_bSbox_L15 ;
    wire Inst_bSbox_L14 ;
    wire Inst_bSbox_L13 ;
    wire Inst_bSbox_L12 ;
    wire Inst_bSbox_L11 ;
    wire Inst_bSbox_L10 ;
    wire Inst_bSbox_L9 ;
    wire Inst_bSbox_L8 ;
    wire Inst_bSbox_L7 ;
    wire Inst_bSbox_L6 ;
    wire Inst_bSbox_L5 ;
    wire Inst_bSbox_L4 ;
    wire Inst_bSbox_L3 ;
    wire Inst_bSbox_L2 ;
    wire Inst_bSbox_L1 ;
    wire Inst_bSbox_L0 ;
    wire Inst_bSbox_M63 ;
    wire Inst_bSbox_M62 ;
    wire Inst_bSbox_M61 ;
    wire Inst_bSbox_M60 ;
    wire Inst_bSbox_M59 ;
    wire Inst_bSbox_M58 ;
    wire Inst_bSbox_M57 ;
    wire Inst_bSbox_M56 ;
    wire Inst_bSbox_M55 ;
    wire Inst_bSbox_M54 ;
    wire Inst_bSbox_M53 ;
    wire Inst_bSbox_M52 ;
    wire Inst_bSbox_M51 ;
    wire Inst_bSbox_M50 ;
    wire Inst_bSbox_M49 ;
    wire Inst_bSbox_M48 ;
    wire Inst_bSbox_M47 ;
    wire Inst_bSbox_M46 ;
    wire Inst_bSbox_M45 ;
    wire Inst_bSbox_M44 ;
    wire Inst_bSbox_M43 ;
    wire Inst_bSbox_M42 ;
    wire Inst_bSbox_M41 ;
    wire Inst_bSbox_M40 ;
    wire Inst_bSbox_M39 ;
    wire Inst_bSbox_M38 ;
    wire Inst_bSbox_M37 ;
    wire Inst_bSbox_M36 ;
    wire Inst_bSbox_M35 ;
    wire Inst_bSbox_M34 ;
    wire Inst_bSbox_M33 ;
    wire Inst_bSbox_M32 ;
    wire Inst_bSbox_M31 ;
    wire Inst_bSbox_M30 ;
    wire Inst_bSbox_M29 ;
    wire Inst_bSbox_M28 ;
    wire Inst_bSbox_M27 ;
    wire Inst_bSbox_M26 ;
    wire Inst_bSbox_M25 ;
    wire Inst_bSbox_M24 ;
    wire Inst_bSbox_M23 ;
    wire Inst_bSbox_M22 ;
    wire Inst_bSbox_M21 ;
    wire Inst_bSbox_M20 ;
    wire Inst_bSbox_M19 ;
    wire Inst_bSbox_M18 ;
    wire Inst_bSbox_M17 ;
    wire Inst_bSbox_M16 ;
    wire Inst_bSbox_M15 ;
    wire Inst_bSbox_M14 ;
    wire Inst_bSbox_M13 ;
    wire Inst_bSbox_M12 ;
    wire Inst_bSbox_M11 ;
    wire Inst_bSbox_M10 ;
    wire Inst_bSbox_M9 ;
    wire Inst_bSbox_M8 ;
    wire Inst_bSbox_M7 ;
    wire Inst_bSbox_M6 ;
    wire Inst_bSbox_M5 ;
    wire Inst_bSbox_M4 ;
    wire Inst_bSbox_M3 ;
    wire Inst_bSbox_M2 ;
    wire Inst_bSbox_M1 ;
    wire Inst_bSbox_T27 ;
    wire Inst_bSbox_T26 ;
    wire Inst_bSbox_T25 ;
    wire Inst_bSbox_T24 ;
    wire Inst_bSbox_T23 ;
    wire Inst_bSbox_T22 ;
    wire Inst_bSbox_T21 ;
    wire Inst_bSbox_T20 ;
    wire Inst_bSbox_T19 ;
    wire Inst_bSbox_T18 ;
    wire Inst_bSbox_T17 ;
    wire Inst_bSbox_T16 ;
    wire Inst_bSbox_T15 ;
    wire Inst_bSbox_T14 ;
    wire Inst_bSbox_T13 ;
    wire Inst_bSbox_T12 ;
    wire Inst_bSbox_T11 ;
    wire Inst_bSbox_T10 ;
    wire Inst_bSbox_T9 ;
    wire Inst_bSbox_T8 ;
    wire Inst_bSbox_T7 ;
    wire Inst_bSbox_T6 ;
    wire Inst_bSbox_T5 ;
    wire Inst_bSbox_T4 ;
    wire Inst_bSbox_T3 ;
    wire Inst_bSbox_T2 ;
    wire Inst_bSbox_T1 ;
    wire [7:0] SboxOut ;
    wire [7:0] StateOutXORroundKey ;
    wire [7:0] StateIn ;
    wire [31:0] StateInMC ;
    wire [31:0] MCout ;
    wire [7:0] keyStateIn ;
    wire [7:0] roundConstant ;
    wire [7:0] keySBIn ;
    wire [7:0] SboxIn ;
    wire [7:0] stateArray_input_MC ;
    wire [7:0] stateArray_outS30ser_MC ;
    wire [7:0] stateArray_outS20ser_MC ;
    wire [7:0] stateArray_outS10ser_MC ;
    wire [7:0] stateArray_inS33ser ;
    wire [7:0] stateArray_inS32ser ;
    wire [7:0] stateArray_inS31ser ;
    wire [7:0] stateArray_inS30ser ;
    wire [7:0] stateArray_inS23ser ;
    wire [7:0] stateArray_inS22ser ;
    wire [7:0] stateArray_inS21ser ;
    wire [7:0] stateArray_inS20ser ;
    wire [7:0] stateArray_inS13ser ;
    wire [7:0] stateArray_inS12ser ;
    wire [7:0] stateArray_inS11ser ;
    wire [7:0] stateArray_inS10ser ;
    wire [7:0] stateArray_inS03ser ;
    wire [7:0] stateArray_inS02ser ;
    wire [7:0] stateArray_inS01ser ;
    wire [7:0] stateArray_inS00ser ;
    wire [7:0] KeyArray_outS01ser_p ;
    wire [7:0] KeyArray_outS01ser_XOR_00 ;
    wire [7:0] KeyArray_outS33ser ;
    wire [7:0] KeyArray_inS33ser ;
    wire [7:0] KeyArray_outS32ser ;
    wire [7:0] KeyArray_inS32ser ;
    wire [7:0] KeyArray_outS31ser ;
    wire [7:0] KeyArray_inS31ser ;
    wire [7:0] KeyArray_outS30ser ;
    wire [7:0] KeyArray_inS30par ;
    wire [7:0] KeyArray_inS30ser ;
    wire [7:0] KeyArray_outS23ser ;
    wire [7:0] KeyArray_inS23ser ;
    wire [7:0] KeyArray_outS22ser ;
    wire [7:0] KeyArray_inS22ser ;
    wire [7:0] KeyArray_outS21ser ;
    wire [7:0] KeyArray_inS21ser ;
    wire [7:0] KeyArray_outS20ser ;
    wire [7:0] KeyArray_inS20ser ;
    wire [7:0] KeyArray_inS13ser ;
    wire [7:0] KeyArray_outS12ser ;
    wire [7:0] KeyArray_inS12ser ;
    wire [7:0] KeyArray_outS11ser ;
    wire [7:0] KeyArray_inS11ser ;
    wire [7:0] KeyArray_outS10ser ;
    wire [7:0] KeyArray_inS10ser ;
    wire [7:0] KeyArray_outS03ser ;
    wire [7:0] KeyArray_inS03ser ;
    wire [7:0] KeyArray_outS02ser ;
    wire [7:0] KeyArray_inS02ser ;
    wire [7:0] KeyArray_inS01ser ;
    wire [7:0] KeyArray_inS00ser ;
    wire [7:0] MixColumns_line0_S13 ;
    wire [4:1] MixColumns_line0_S02 ;
    wire [4:1] MixColumns_line0_timesTHREE_input2 ;
    wire [7:0] MixColumns_line1_S13 ;
    wire [4:1] MixColumns_line1_timesTHREE_input2 ;
    wire [7:0] MixColumns_line2_S13 ;
    wire [4:1] MixColumns_line2_timesTHREE_input2 ;
    wire [7:0] MixColumns_line3_S13 ;
    wire LMDPL_pre1 ;
    wire LMDPL_pre2 ;
    wire mid_rst ;
    wire new_AGEMA_signal_1987 ;
    wire new_AGEMA_signal_1988 ;
    wire new_AGEMA_signal_1989 ;
    wire new_AGEMA_signal_1990 ;
    wire new_AGEMA_signal_1991 ;
    wire new_AGEMA_signal_1993 ;
    wire new_AGEMA_signal_1994 ;
    wire new_AGEMA_signal_1995 ;
    wire new_AGEMA_signal_1996 ;
    wire new_AGEMA_signal_1997 ;
    wire new_AGEMA_signal_1999 ;
    wire new_AGEMA_signal_2000 ;
    wire new_AGEMA_signal_2001 ;
    wire new_AGEMA_signal_2002 ;
    wire new_AGEMA_signal_2003 ;
    wire new_AGEMA_signal_2005 ;
    wire new_AGEMA_signal_2006 ;
    wire new_AGEMA_signal_2007 ;
    wire new_AGEMA_signal_2008 ;
    wire new_AGEMA_signal_2009 ;
    wire new_AGEMA_signal_2011 ;
    wire new_AGEMA_signal_2012 ;
    wire new_AGEMA_signal_2013 ;
    wire new_AGEMA_signal_2014 ;
    wire new_AGEMA_signal_2015 ;
    wire new_AGEMA_signal_2017 ;
    wire new_AGEMA_signal_2018 ;
    wire new_AGEMA_signal_2019 ;
    wire new_AGEMA_signal_2020 ;
    wire new_AGEMA_signal_2021 ;
    wire new_AGEMA_signal_2023 ;
    wire new_AGEMA_signal_2024 ;
    wire new_AGEMA_signal_2025 ;
    wire new_AGEMA_signal_2026 ;
    wire new_AGEMA_signal_2027 ;
    wire new_AGEMA_signal_2029 ;
    wire new_AGEMA_signal_2030 ;
    wire new_AGEMA_signal_2031 ;
    wire new_AGEMA_signal_2032 ;
    wire new_AGEMA_signal_2033 ;
    wire new_AGEMA_signal_2034 ;
    wire new_AGEMA_signal_2035 ;
    wire new_AGEMA_signal_2036 ;
    wire new_AGEMA_signal_2037 ;
    wire new_AGEMA_signal_2038 ;
    wire new_AGEMA_signal_2039 ;
    wire new_AGEMA_signal_2040 ;
    wire new_AGEMA_signal_2041 ;
    wire new_AGEMA_signal_2042 ;
    wire new_AGEMA_signal_2043 ;
    wire new_AGEMA_signal_2044 ;
    wire new_AGEMA_signal_2045 ;
    wire new_AGEMA_signal_2046 ;
    wire new_AGEMA_signal_2047 ;
    wire new_AGEMA_signal_2048 ;
    wire new_AGEMA_signal_2049 ;
    wire new_AGEMA_signal_2050 ;
    wire new_AGEMA_signal_2051 ;
    wire new_AGEMA_signal_2052 ;
    wire new_AGEMA_signal_2053 ;
    wire new_AGEMA_signal_2054 ;
    wire new_AGEMA_signal_2055 ;
    wire new_AGEMA_signal_2056 ;
    wire new_AGEMA_signal_2057 ;
    wire new_AGEMA_signal_2058 ;
    wire new_AGEMA_signal_2059 ;
    wire new_AGEMA_signal_2060 ;
    wire new_AGEMA_signal_2061 ;
    wire new_AGEMA_signal_2062 ;
    wire new_AGEMA_signal_2063 ;
    wire new_AGEMA_signal_2064 ;
    wire new_AGEMA_signal_2065 ;
    wire new_AGEMA_signal_2067 ;
    wire new_AGEMA_signal_2069 ;
    wire new_AGEMA_signal_2070 ;
    wire new_AGEMA_signal_2071 ;
    wire new_AGEMA_signal_2073 ;
    wire new_AGEMA_signal_2075 ;
    wire new_AGEMA_signal_2076 ;
    wire new_AGEMA_signal_2077 ;
    wire new_AGEMA_signal_2079 ;
    wire new_AGEMA_signal_2081 ;
    wire new_AGEMA_signal_2082 ;
    wire new_AGEMA_signal_2083 ;
    wire new_AGEMA_signal_2085 ;
    wire new_AGEMA_signal_2087 ;
    wire new_AGEMA_signal_2088 ;
    wire new_AGEMA_signal_2089 ;
    wire new_AGEMA_signal_2091 ;
    wire new_AGEMA_signal_2093 ;
    wire new_AGEMA_signal_2094 ;
    wire new_AGEMA_signal_2095 ;
    wire new_AGEMA_signal_2097 ;
    wire new_AGEMA_signal_2099 ;
    wire new_AGEMA_signal_2100 ;
    wire new_AGEMA_signal_2101 ;
    wire new_AGEMA_signal_2103 ;
    wire new_AGEMA_signal_2105 ;
    wire new_AGEMA_signal_2106 ;
    wire new_AGEMA_signal_2107 ;
    wire new_AGEMA_signal_2109 ;
    wire new_AGEMA_signal_2111 ;
    wire new_AGEMA_signal_2112 ;
    wire new_AGEMA_signal_2113 ;
    wire new_AGEMA_signal_2114 ;
    wire new_AGEMA_signal_2115 ;
    wire new_AGEMA_signal_2116 ;
    wire new_AGEMA_signal_2117 ;
    wire new_AGEMA_signal_2118 ;
    wire new_AGEMA_signal_2119 ;
    wire new_AGEMA_signal_2121 ;
    wire new_AGEMA_signal_2123 ;
    wire new_AGEMA_signal_2124 ;
    wire new_AGEMA_signal_2125 ;
    wire new_AGEMA_signal_2127 ;
    wire new_AGEMA_signal_2128 ;
    wire new_AGEMA_signal_2129 ;
    wire new_AGEMA_signal_2131 ;
    wire new_AGEMA_signal_2132 ;
    wire new_AGEMA_signal_2133 ;
    wire new_AGEMA_signal_2135 ;
    wire new_AGEMA_signal_2137 ;
    wire new_AGEMA_signal_2138 ;
    wire new_AGEMA_signal_2139 ;
    wire new_AGEMA_signal_2141 ;
    wire new_AGEMA_signal_2142 ;
    wire new_AGEMA_signal_2143 ;
    wire new_AGEMA_signal_2145 ;
    wire new_AGEMA_signal_2146 ;
    wire new_AGEMA_signal_2147 ;
    wire new_AGEMA_signal_2148 ;
    wire new_AGEMA_signal_2149 ;
    wire new_AGEMA_signal_2150 ;
    wire new_AGEMA_signal_2151 ;
    wire new_AGEMA_signal_2152 ;
    wire new_AGEMA_signal_2153 ;
    wire new_AGEMA_signal_2154 ;
    wire new_AGEMA_signal_2155 ;
    wire new_AGEMA_signal_2156 ;
    wire new_AGEMA_signal_2157 ;
    wire new_AGEMA_signal_2158 ;
    wire new_AGEMA_signal_2159 ;
    wire new_AGEMA_signal_2160 ;
    wire new_AGEMA_signal_2161 ;
    wire new_AGEMA_signal_2162 ;
    wire new_AGEMA_signal_2163 ;
    wire new_AGEMA_signal_2164 ;
    wire new_AGEMA_signal_2165 ;
    wire new_AGEMA_signal_2166 ;
    wire new_AGEMA_signal_2167 ;
    wire new_AGEMA_signal_2168 ;
    wire new_AGEMA_signal_2169 ;
    wire new_AGEMA_signal_2170 ;
    wire new_AGEMA_signal_2171 ;
    wire new_AGEMA_signal_2172 ;
    wire new_AGEMA_signal_2173 ;
    wire new_AGEMA_signal_2174 ;
    wire new_AGEMA_signal_2175 ;
    wire new_AGEMA_signal_2176 ;
    wire new_AGEMA_signal_2177 ;
    wire new_AGEMA_signal_2178 ;
    wire new_AGEMA_signal_2179 ;
    wire new_AGEMA_signal_2180 ;
    wire new_AGEMA_signal_2181 ;
    wire new_AGEMA_signal_2182 ;
    wire new_AGEMA_signal_2183 ;
    wire new_AGEMA_signal_2184 ;
    wire new_AGEMA_signal_2185 ;
    wire new_AGEMA_signal_2186 ;
    wire new_AGEMA_signal_2187 ;
    wire new_AGEMA_signal_2188 ;
    wire new_AGEMA_signal_2189 ;
    wire new_AGEMA_signal_2190 ;
    wire new_AGEMA_signal_2191 ;
    wire new_AGEMA_signal_2192 ;
    wire new_AGEMA_signal_2193 ;
    wire new_AGEMA_signal_2194 ;
    wire new_AGEMA_signal_2195 ;
    wire new_AGEMA_signal_2196 ;
    wire new_AGEMA_signal_2197 ;
    wire new_AGEMA_signal_2198 ;
    wire new_AGEMA_signal_2199 ;
    wire new_AGEMA_signal_2200 ;
    wire new_AGEMA_signal_2201 ;
    wire new_AGEMA_signal_2202 ;
    wire new_AGEMA_signal_2203 ;
    wire new_AGEMA_signal_2204 ;
    wire new_AGEMA_signal_2205 ;
    wire new_AGEMA_signal_2206 ;
    wire new_AGEMA_signal_2207 ;
    wire new_AGEMA_signal_2208 ;
    wire new_AGEMA_signal_2209 ;
    wire new_AGEMA_signal_2210 ;
    wire new_AGEMA_signal_2211 ;
    wire new_AGEMA_signal_2212 ;
    wire new_AGEMA_signal_2213 ;
    wire new_AGEMA_signal_2214 ;
    wire new_AGEMA_signal_2215 ;
    wire new_AGEMA_signal_2216 ;
    wire new_AGEMA_signal_2217 ;
    wire new_AGEMA_signal_2218 ;
    wire new_AGEMA_signal_2219 ;
    wire new_AGEMA_signal_2220 ;
    wire new_AGEMA_signal_2221 ;
    wire new_AGEMA_signal_2222 ;
    wire new_AGEMA_signal_2223 ;
    wire new_AGEMA_signal_2224 ;
    wire new_AGEMA_signal_2225 ;
    wire new_AGEMA_signal_2226 ;
    wire new_AGEMA_signal_2227 ;
    wire new_AGEMA_signal_2228 ;
    wire new_AGEMA_signal_2229 ;
    wire new_AGEMA_signal_2230 ;
    wire new_AGEMA_signal_2231 ;
    wire new_AGEMA_signal_2232 ;
    wire new_AGEMA_signal_2233 ;
    wire new_AGEMA_signal_2234 ;
    wire new_AGEMA_signal_2235 ;
    wire new_AGEMA_signal_2236 ;
    wire new_AGEMA_signal_2237 ;
    wire new_AGEMA_signal_2238 ;
    wire new_AGEMA_signal_2239 ;
    wire new_AGEMA_signal_2240 ;
    wire new_AGEMA_signal_2241 ;
    wire new_AGEMA_signal_2242 ;
    wire new_AGEMA_signal_2243 ;
    wire new_AGEMA_signal_2244 ;
    wire new_AGEMA_signal_2245 ;
    wire new_AGEMA_signal_2246 ;
    wire new_AGEMA_signal_2247 ;
    wire new_AGEMA_signal_2248 ;
    wire new_AGEMA_signal_2249 ;
    wire new_AGEMA_signal_2250 ;
    wire new_AGEMA_signal_2251 ;
    wire new_AGEMA_signal_2252 ;
    wire new_AGEMA_signal_2253 ;
    wire new_AGEMA_signal_2254 ;
    wire new_AGEMA_signal_2255 ;
    wire new_AGEMA_signal_2256 ;
    wire new_AGEMA_signal_2257 ;
    wire new_AGEMA_signal_2258 ;
    wire new_AGEMA_signal_2259 ;
    wire new_AGEMA_signal_2260 ;
    wire new_AGEMA_signal_2261 ;
    wire new_AGEMA_signal_2262 ;
    wire new_AGEMA_signal_2263 ;
    wire new_AGEMA_signal_2264 ;
    wire new_AGEMA_signal_2265 ;
    wire new_AGEMA_signal_2266 ;
    wire new_AGEMA_signal_2267 ;
    wire new_AGEMA_signal_2268 ;
    wire new_AGEMA_signal_2269 ;
    wire new_AGEMA_signal_2270 ;
    wire new_AGEMA_signal_2271 ;
    wire new_AGEMA_signal_2272 ;
    wire new_AGEMA_signal_2273 ;
    wire new_AGEMA_signal_2274 ;
    wire new_AGEMA_signal_2275 ;
    wire new_AGEMA_signal_2276 ;
    wire new_AGEMA_signal_2277 ;
    wire new_AGEMA_signal_2278 ;
    wire new_AGEMA_signal_2279 ;
    wire new_AGEMA_signal_2280 ;
    wire new_AGEMA_signal_2281 ;
    wire new_AGEMA_signal_2282 ;
    wire new_AGEMA_signal_2283 ;
    wire new_AGEMA_signal_2284 ;
    wire new_AGEMA_signal_2285 ;
    wire new_AGEMA_signal_2286 ;
    wire new_AGEMA_signal_2287 ;
    wire new_AGEMA_signal_2288 ;
    wire new_AGEMA_signal_2289 ;
    wire new_AGEMA_signal_2290 ;
    wire new_AGEMA_signal_2291 ;
    wire new_AGEMA_signal_2292 ;
    wire new_AGEMA_signal_2293 ;
    wire new_AGEMA_signal_2294 ;
    wire new_AGEMA_signal_2295 ;
    wire new_AGEMA_signal_2296 ;
    wire new_AGEMA_signal_2297 ;
    wire new_AGEMA_signal_2298 ;
    wire new_AGEMA_signal_2299 ;
    wire new_AGEMA_signal_2300 ;
    wire new_AGEMA_signal_2301 ;
    wire new_AGEMA_signal_2302 ;
    wire new_AGEMA_signal_2303 ;
    wire new_AGEMA_signal_2304 ;
    wire new_AGEMA_signal_2305 ;
    wire new_AGEMA_signal_2306 ;
    wire new_AGEMA_signal_2307 ;
    wire new_AGEMA_signal_2308 ;
    wire new_AGEMA_signal_2309 ;
    wire new_AGEMA_signal_2310 ;
    wire new_AGEMA_signal_2311 ;
    wire new_AGEMA_signal_2312 ;
    wire new_AGEMA_signal_2313 ;
    wire new_AGEMA_signal_2314 ;
    wire new_AGEMA_signal_2315 ;
    wire new_AGEMA_signal_2316 ;
    wire new_AGEMA_signal_2317 ;
    wire new_AGEMA_signal_2318 ;
    wire new_AGEMA_signal_2319 ;
    wire new_AGEMA_signal_2320 ;
    wire new_AGEMA_signal_2321 ;
    wire new_AGEMA_signal_2322 ;
    wire new_AGEMA_signal_2323 ;
    wire new_AGEMA_signal_2324 ;
    wire new_AGEMA_signal_2325 ;
    wire new_AGEMA_signal_2326 ;
    wire new_AGEMA_signal_2327 ;
    wire new_AGEMA_signal_2328 ;
    wire new_AGEMA_signal_2329 ;
    wire new_AGEMA_signal_2330 ;
    wire new_AGEMA_signal_2331 ;
    wire new_AGEMA_signal_2332 ;
    wire new_AGEMA_signal_2333 ;
    wire new_AGEMA_signal_2335 ;
    wire new_AGEMA_signal_2336 ;
    wire new_AGEMA_signal_2337 ;
    wire new_AGEMA_signal_2338 ;
    wire new_AGEMA_signal_2339 ;
    wire new_AGEMA_signal_2341 ;
    wire new_AGEMA_signal_2342 ;
    wire new_AGEMA_signal_2343 ;
    wire new_AGEMA_signal_2344 ;
    wire new_AGEMA_signal_2345 ;
    wire new_AGEMA_signal_2347 ;
    wire new_AGEMA_signal_2348 ;
    wire new_AGEMA_signal_2349 ;
    wire new_AGEMA_signal_2350 ;
    wire new_AGEMA_signal_2351 ;
    wire new_AGEMA_signal_2353 ;
    wire new_AGEMA_signal_2354 ;
    wire new_AGEMA_signal_2355 ;
    wire new_AGEMA_signal_2356 ;
    wire new_AGEMA_signal_2357 ;
    wire new_AGEMA_signal_2359 ;
    wire new_AGEMA_signal_2360 ;
    wire new_AGEMA_signal_2361 ;
    wire new_AGEMA_signal_2362 ;
    wire new_AGEMA_signal_2363 ;
    wire new_AGEMA_signal_2365 ;
    wire new_AGEMA_signal_2366 ;
    wire new_AGEMA_signal_2367 ;
    wire new_AGEMA_signal_2368 ;
    wire new_AGEMA_signal_2369 ;
    wire new_AGEMA_signal_2371 ;
    wire new_AGEMA_signal_2372 ;
    wire new_AGEMA_signal_2373 ;
    wire new_AGEMA_signal_2374 ;
    wire new_AGEMA_signal_2375 ;
    wire new_AGEMA_signal_2377 ;
    wire new_AGEMA_signal_2378 ;
    wire new_AGEMA_signal_2379 ;
    wire new_AGEMA_signal_2380 ;
    wire new_AGEMA_signal_2381 ;
    wire new_AGEMA_signal_2383 ;
    wire new_AGEMA_signal_2384 ;
    wire new_AGEMA_signal_2385 ;
    wire new_AGEMA_signal_2386 ;
    wire new_AGEMA_signal_2387 ;
    wire new_AGEMA_signal_2389 ;
    wire new_AGEMA_signal_2390 ;
    wire new_AGEMA_signal_2391 ;
    wire new_AGEMA_signal_2392 ;
    wire new_AGEMA_signal_2393 ;
    wire new_AGEMA_signal_2395 ;
    wire new_AGEMA_signal_2396 ;
    wire new_AGEMA_signal_2397 ;
    wire new_AGEMA_signal_2398 ;
    wire new_AGEMA_signal_2399 ;
    wire new_AGEMA_signal_2401 ;
    wire new_AGEMA_signal_2402 ;
    wire new_AGEMA_signal_2403 ;
    wire new_AGEMA_signal_2404 ;
    wire new_AGEMA_signal_2405 ;
    wire new_AGEMA_signal_2407 ;
    wire new_AGEMA_signal_2408 ;
    wire new_AGEMA_signal_2409 ;
    wire new_AGEMA_signal_2410 ;
    wire new_AGEMA_signal_2411 ;
    wire new_AGEMA_signal_2413 ;
    wire new_AGEMA_signal_2414 ;
    wire new_AGEMA_signal_2415 ;
    wire new_AGEMA_signal_2416 ;
    wire new_AGEMA_signal_2417 ;
    wire new_AGEMA_signal_2419 ;
    wire new_AGEMA_signal_2420 ;
    wire new_AGEMA_signal_2421 ;
    wire new_AGEMA_signal_2422 ;
    wire new_AGEMA_signal_2423 ;
    wire new_AGEMA_signal_2425 ;
    wire new_AGEMA_signal_2426 ;
    wire new_AGEMA_signal_2427 ;
    wire new_AGEMA_signal_2428 ;
    wire new_AGEMA_signal_2429 ;
    wire new_AGEMA_signal_2430 ;
    wire new_AGEMA_signal_2431 ;
    wire new_AGEMA_signal_2433 ;
    wire new_AGEMA_signal_2434 ;
    wire new_AGEMA_signal_2435 ;
    wire new_AGEMA_signal_2436 ;
    wire new_AGEMA_signal_2437 ;
    wire new_AGEMA_signal_2439 ;
    wire new_AGEMA_signal_2440 ;
    wire new_AGEMA_signal_2441 ;
    wire new_AGEMA_signal_2442 ;
    wire new_AGEMA_signal_2443 ;
    wire new_AGEMA_signal_2445 ;
    wire new_AGEMA_signal_2446 ;
    wire new_AGEMA_signal_2447 ;
    wire new_AGEMA_signal_2448 ;
    wire new_AGEMA_signal_2449 ;
    wire new_AGEMA_signal_2451 ;
    wire new_AGEMA_signal_2452 ;
    wire new_AGEMA_signal_2453 ;
    wire new_AGEMA_signal_2454 ;
    wire new_AGEMA_signal_2455 ;
    wire new_AGEMA_signal_2457 ;
    wire new_AGEMA_signal_2458 ;
    wire new_AGEMA_signal_2459 ;
    wire new_AGEMA_signal_2460 ;
    wire new_AGEMA_signal_2461 ;
    wire new_AGEMA_signal_2463 ;
    wire new_AGEMA_signal_2464 ;
    wire new_AGEMA_signal_2465 ;
    wire new_AGEMA_signal_2466 ;
    wire new_AGEMA_signal_2467 ;
    wire new_AGEMA_signal_2469 ;
    wire new_AGEMA_signal_2470 ;
    wire new_AGEMA_signal_2471 ;
    wire new_AGEMA_signal_2472 ;
    wire new_AGEMA_signal_2473 ;
    wire new_AGEMA_signal_2475 ;
    wire new_AGEMA_signal_2476 ;
    wire new_AGEMA_signal_2477 ;
    wire new_AGEMA_signal_2478 ;
    wire new_AGEMA_signal_2479 ;
    wire new_AGEMA_signal_2480 ;
    wire new_AGEMA_signal_2481 ;
    wire new_AGEMA_signal_2483 ;
    wire new_AGEMA_signal_2484 ;
    wire new_AGEMA_signal_2485 ;
    wire new_AGEMA_signal_2486 ;
    wire new_AGEMA_signal_2487 ;
    wire new_AGEMA_signal_2489 ;
    wire new_AGEMA_signal_2490 ;
    wire new_AGEMA_signal_2491 ;
    wire new_AGEMA_signal_2492 ;
    wire new_AGEMA_signal_2493 ;
    wire new_AGEMA_signal_2495 ;
    wire new_AGEMA_signal_2496 ;
    wire new_AGEMA_signal_2497 ;
    wire new_AGEMA_signal_2498 ;
    wire new_AGEMA_signal_2499 ;
    wire new_AGEMA_signal_2501 ;
    wire new_AGEMA_signal_2502 ;
    wire new_AGEMA_signal_2503 ;
    wire new_AGEMA_signal_2504 ;
    wire new_AGEMA_signal_2505 ;
    wire new_AGEMA_signal_2507 ;
    wire new_AGEMA_signal_2508 ;
    wire new_AGEMA_signal_2509 ;
    wire new_AGEMA_signal_2510 ;
    wire new_AGEMA_signal_2511 ;
    wire new_AGEMA_signal_2513 ;
    wire new_AGEMA_signal_2514 ;
    wire new_AGEMA_signal_2515 ;
    wire new_AGEMA_signal_2516 ;
    wire new_AGEMA_signal_2517 ;
    wire new_AGEMA_signal_2519 ;
    wire new_AGEMA_signal_2520 ;
    wire new_AGEMA_signal_2521 ;
    wire new_AGEMA_signal_2522 ;
    wire new_AGEMA_signal_2523 ;
    wire new_AGEMA_signal_2525 ;
    wire new_AGEMA_signal_2526 ;
    wire new_AGEMA_signal_2527 ;
    wire new_AGEMA_signal_2528 ;
    wire new_AGEMA_signal_2529 ;
    wire new_AGEMA_signal_2531 ;
    wire new_AGEMA_signal_2532 ;
    wire new_AGEMA_signal_2533 ;
    wire new_AGEMA_signal_2534 ;
    wire new_AGEMA_signal_2535 ;
    wire new_AGEMA_signal_2537 ;
    wire new_AGEMA_signal_2538 ;
    wire new_AGEMA_signal_2539 ;
    wire new_AGEMA_signal_2540 ;
    wire new_AGEMA_signal_2541 ;
    wire new_AGEMA_signal_2543 ;
    wire new_AGEMA_signal_2544 ;
    wire new_AGEMA_signal_2545 ;
    wire new_AGEMA_signal_2546 ;
    wire new_AGEMA_signal_2547 ;
    wire new_AGEMA_signal_2549 ;
    wire new_AGEMA_signal_2550 ;
    wire new_AGEMA_signal_2551 ;
    wire new_AGEMA_signal_2552 ;
    wire new_AGEMA_signal_2553 ;
    wire new_AGEMA_signal_2555 ;
    wire new_AGEMA_signal_2556 ;
    wire new_AGEMA_signal_2557 ;
    wire new_AGEMA_signal_2558 ;
    wire new_AGEMA_signal_2559 ;
    wire new_AGEMA_signal_2561 ;
    wire new_AGEMA_signal_2562 ;
    wire new_AGEMA_signal_2563 ;
    wire new_AGEMA_signal_2564 ;
    wire new_AGEMA_signal_2565 ;
    wire new_AGEMA_signal_2567 ;
    wire new_AGEMA_signal_2568 ;
    wire new_AGEMA_signal_2569 ;
    wire new_AGEMA_signal_2570 ;
    wire new_AGEMA_signal_2571 ;
    wire new_AGEMA_signal_2573 ;
    wire new_AGEMA_signal_2574 ;
    wire new_AGEMA_signal_2575 ;
    wire new_AGEMA_signal_2576 ;
    wire new_AGEMA_signal_2577 ;
    wire new_AGEMA_signal_2578 ;
    wire new_AGEMA_signal_2579 ;
    wire new_AGEMA_signal_2581 ;
    wire new_AGEMA_signal_2582 ;
    wire new_AGEMA_signal_2583 ;
    wire new_AGEMA_signal_2584 ;
    wire new_AGEMA_signal_2585 ;
    wire new_AGEMA_signal_2587 ;
    wire new_AGEMA_signal_2588 ;
    wire new_AGEMA_signal_2589 ;
    wire new_AGEMA_signal_2590 ;
    wire new_AGEMA_signal_2591 ;
    wire new_AGEMA_signal_2593 ;
    wire new_AGEMA_signal_2594 ;
    wire new_AGEMA_signal_2595 ;
    wire new_AGEMA_signal_2596 ;
    wire new_AGEMA_signal_2597 ;
    wire new_AGEMA_signal_2599 ;
    wire new_AGEMA_signal_2600 ;
    wire new_AGEMA_signal_2601 ;
    wire new_AGEMA_signal_2602 ;
    wire new_AGEMA_signal_2603 ;
    wire new_AGEMA_signal_2605 ;
    wire new_AGEMA_signal_2606 ;
    wire new_AGEMA_signal_2607 ;
    wire new_AGEMA_signal_2608 ;
    wire new_AGEMA_signal_2609 ;
    wire new_AGEMA_signal_2611 ;
    wire new_AGEMA_signal_2612 ;
    wire new_AGEMA_signal_2613 ;
    wire new_AGEMA_signal_2614 ;
    wire new_AGEMA_signal_2615 ;
    wire new_AGEMA_signal_2617 ;
    wire new_AGEMA_signal_2618 ;
    wire new_AGEMA_signal_2619 ;
    wire new_AGEMA_signal_2620 ;
    wire new_AGEMA_signal_2621 ;
    wire new_AGEMA_signal_2623 ;
    wire new_AGEMA_signal_2624 ;
    wire new_AGEMA_signal_2625 ;
    wire new_AGEMA_signal_2626 ;
    wire new_AGEMA_signal_2627 ;
    wire new_AGEMA_signal_2628 ;
    wire new_AGEMA_signal_2629 ;
    wire new_AGEMA_signal_2631 ;
    wire new_AGEMA_signal_2632 ;
    wire new_AGEMA_signal_2633 ;
    wire new_AGEMA_signal_2634 ;
    wire new_AGEMA_signal_2635 ;
    wire new_AGEMA_signal_2637 ;
    wire new_AGEMA_signal_2638 ;
    wire new_AGEMA_signal_2639 ;
    wire new_AGEMA_signal_2640 ;
    wire new_AGEMA_signal_2641 ;
    wire new_AGEMA_signal_2643 ;
    wire new_AGEMA_signal_2644 ;
    wire new_AGEMA_signal_2645 ;
    wire new_AGEMA_signal_2646 ;
    wire new_AGEMA_signal_2647 ;
    wire new_AGEMA_signal_2649 ;
    wire new_AGEMA_signal_2650 ;
    wire new_AGEMA_signal_2651 ;
    wire new_AGEMA_signal_2652 ;
    wire new_AGEMA_signal_2653 ;
    wire new_AGEMA_signal_2655 ;
    wire new_AGEMA_signal_2656 ;
    wire new_AGEMA_signal_2657 ;
    wire new_AGEMA_signal_2658 ;
    wire new_AGEMA_signal_2659 ;
    wire new_AGEMA_signal_2661 ;
    wire new_AGEMA_signal_2662 ;
    wire new_AGEMA_signal_2663 ;
    wire new_AGEMA_signal_2664 ;
    wire new_AGEMA_signal_2665 ;
    wire new_AGEMA_signal_2667 ;
    wire new_AGEMA_signal_2668 ;
    wire new_AGEMA_signal_2669 ;
    wire new_AGEMA_signal_2670 ;
    wire new_AGEMA_signal_2671 ;
    wire new_AGEMA_signal_2673 ;
    wire new_AGEMA_signal_2674 ;
    wire new_AGEMA_signal_2675 ;
    wire new_AGEMA_signal_2676 ;
    wire new_AGEMA_signal_2677 ;
    wire new_AGEMA_signal_2679 ;
    wire new_AGEMA_signal_2680 ;
    wire new_AGEMA_signal_2681 ;
    wire new_AGEMA_signal_2682 ;
    wire new_AGEMA_signal_2683 ;
    wire new_AGEMA_signal_2685 ;
    wire new_AGEMA_signal_2686 ;
    wire new_AGEMA_signal_2687 ;
    wire new_AGEMA_signal_2688 ;
    wire new_AGEMA_signal_2689 ;
    wire new_AGEMA_signal_2691 ;
    wire new_AGEMA_signal_2692 ;
    wire new_AGEMA_signal_2693 ;
    wire new_AGEMA_signal_2694 ;
    wire new_AGEMA_signal_2695 ;
    wire new_AGEMA_signal_2697 ;
    wire new_AGEMA_signal_2698 ;
    wire new_AGEMA_signal_2699 ;
    wire new_AGEMA_signal_2700 ;
    wire new_AGEMA_signal_2701 ;
    wire new_AGEMA_signal_2703 ;
    wire new_AGEMA_signal_2704 ;
    wire new_AGEMA_signal_2705 ;
    wire new_AGEMA_signal_2706 ;
    wire new_AGEMA_signal_2707 ;
    wire new_AGEMA_signal_2709 ;
    wire new_AGEMA_signal_2710 ;
    wire new_AGEMA_signal_2711 ;
    wire new_AGEMA_signal_2712 ;
    wire new_AGEMA_signal_2713 ;
    wire new_AGEMA_signal_2715 ;
    wire new_AGEMA_signal_2716 ;
    wire new_AGEMA_signal_2717 ;
    wire new_AGEMA_signal_2718 ;
    wire new_AGEMA_signal_2719 ;
    wire new_AGEMA_signal_2721 ;
    wire new_AGEMA_signal_2722 ;
    wire new_AGEMA_signal_2723 ;
    wire new_AGEMA_signal_2724 ;
    wire new_AGEMA_signal_2725 ;
    wire new_AGEMA_signal_2726 ;
    wire new_AGEMA_signal_2727 ;
    wire new_AGEMA_signal_2729 ;
    wire new_AGEMA_signal_2730 ;
    wire new_AGEMA_signal_2731 ;
    wire new_AGEMA_signal_2732 ;
    wire new_AGEMA_signal_2733 ;
    wire new_AGEMA_signal_2735 ;
    wire new_AGEMA_signal_2736 ;
    wire new_AGEMA_signal_2737 ;
    wire new_AGEMA_signal_2738 ;
    wire new_AGEMA_signal_2739 ;
    wire new_AGEMA_signal_2741 ;
    wire new_AGEMA_signal_2742 ;
    wire new_AGEMA_signal_2743 ;
    wire new_AGEMA_signal_2744 ;
    wire new_AGEMA_signal_2745 ;
    wire new_AGEMA_signal_2747 ;
    wire new_AGEMA_signal_2748 ;
    wire new_AGEMA_signal_2749 ;
    wire new_AGEMA_signal_2750 ;
    wire new_AGEMA_signal_2751 ;
    wire new_AGEMA_signal_2753 ;
    wire new_AGEMA_signal_2754 ;
    wire new_AGEMA_signal_2755 ;
    wire new_AGEMA_signal_2756 ;
    wire new_AGEMA_signal_2757 ;
    wire new_AGEMA_signal_2759 ;
    wire new_AGEMA_signal_2760 ;
    wire new_AGEMA_signal_2761 ;
    wire new_AGEMA_signal_2762 ;
    wire new_AGEMA_signal_2763 ;
    wire new_AGEMA_signal_2765 ;
    wire new_AGEMA_signal_2766 ;
    wire new_AGEMA_signal_2767 ;
    wire new_AGEMA_signal_2768 ;
    wire new_AGEMA_signal_2769 ;
    wire new_AGEMA_signal_2771 ;
    wire new_AGEMA_signal_2772 ;
    wire new_AGEMA_signal_2773 ;
    wire new_AGEMA_signal_2774 ;
    wire new_AGEMA_signal_2775 ;
    wire new_AGEMA_signal_2776 ;
    wire new_AGEMA_signal_2777 ;
    wire new_AGEMA_signal_2779 ;
    wire new_AGEMA_signal_2780 ;
    wire new_AGEMA_signal_2781 ;
    wire new_AGEMA_signal_2782 ;
    wire new_AGEMA_signal_2783 ;
    wire new_AGEMA_signal_2785 ;
    wire new_AGEMA_signal_2786 ;
    wire new_AGEMA_signal_2787 ;
    wire new_AGEMA_signal_2788 ;
    wire new_AGEMA_signal_2789 ;
    wire new_AGEMA_signal_2791 ;
    wire new_AGEMA_signal_2792 ;
    wire new_AGEMA_signal_2793 ;
    wire new_AGEMA_signal_2794 ;
    wire new_AGEMA_signal_2795 ;
    wire new_AGEMA_signal_2797 ;
    wire new_AGEMA_signal_2798 ;
    wire new_AGEMA_signal_2799 ;
    wire new_AGEMA_signal_2800 ;
    wire new_AGEMA_signal_2801 ;
    wire new_AGEMA_signal_2803 ;
    wire new_AGEMA_signal_2804 ;
    wire new_AGEMA_signal_2805 ;
    wire new_AGEMA_signal_2806 ;
    wire new_AGEMA_signal_2807 ;
    wire new_AGEMA_signal_2809 ;
    wire new_AGEMA_signal_2810 ;
    wire new_AGEMA_signal_2811 ;
    wire new_AGEMA_signal_2812 ;
    wire new_AGEMA_signal_2813 ;
    wire new_AGEMA_signal_2815 ;
    wire new_AGEMA_signal_2816 ;
    wire new_AGEMA_signal_2817 ;
    wire new_AGEMA_signal_2818 ;
    wire new_AGEMA_signal_2819 ;
    wire new_AGEMA_signal_2821 ;
    wire new_AGEMA_signal_2822 ;
    wire new_AGEMA_signal_2823 ;
    wire new_AGEMA_signal_2824 ;
    wire new_AGEMA_signal_2825 ;
    wire new_AGEMA_signal_2827 ;
    wire new_AGEMA_signal_2828 ;
    wire new_AGEMA_signal_2829 ;
    wire new_AGEMA_signal_2830 ;
    wire new_AGEMA_signal_2831 ;
    wire new_AGEMA_signal_2833 ;
    wire new_AGEMA_signal_2834 ;
    wire new_AGEMA_signal_2835 ;
    wire new_AGEMA_signal_2836 ;
    wire new_AGEMA_signal_2837 ;
    wire new_AGEMA_signal_2839 ;
    wire new_AGEMA_signal_2840 ;
    wire new_AGEMA_signal_2841 ;
    wire new_AGEMA_signal_2842 ;
    wire new_AGEMA_signal_2843 ;
    wire new_AGEMA_signal_2845 ;
    wire new_AGEMA_signal_2846 ;
    wire new_AGEMA_signal_2847 ;
    wire new_AGEMA_signal_2848 ;
    wire new_AGEMA_signal_2849 ;
    wire new_AGEMA_signal_2851 ;
    wire new_AGEMA_signal_2852 ;
    wire new_AGEMA_signal_2853 ;
    wire new_AGEMA_signal_2854 ;
    wire new_AGEMA_signal_2855 ;
    wire new_AGEMA_signal_2857 ;
    wire new_AGEMA_signal_2858 ;
    wire new_AGEMA_signal_2859 ;
    wire new_AGEMA_signal_2860 ;
    wire new_AGEMA_signal_2861 ;
    wire new_AGEMA_signal_2863 ;
    wire new_AGEMA_signal_2864 ;
    wire new_AGEMA_signal_2865 ;
    wire new_AGEMA_signal_2866 ;
    wire new_AGEMA_signal_2867 ;
    wire new_AGEMA_signal_2869 ;
    wire new_AGEMA_signal_2870 ;
    wire new_AGEMA_signal_2871 ;
    wire new_AGEMA_signal_2872 ;
    wire new_AGEMA_signal_2873 ;
    wire new_AGEMA_signal_2874 ;
    wire new_AGEMA_signal_2875 ;
    wire new_AGEMA_signal_2877 ;
    wire new_AGEMA_signal_2878 ;
    wire new_AGEMA_signal_2879 ;
    wire new_AGEMA_signal_2880 ;
    wire new_AGEMA_signal_2881 ;
    wire new_AGEMA_signal_2883 ;
    wire new_AGEMA_signal_2884 ;
    wire new_AGEMA_signal_2885 ;
    wire new_AGEMA_signal_2886 ;
    wire new_AGEMA_signal_2887 ;
    wire new_AGEMA_signal_2889 ;
    wire new_AGEMA_signal_2890 ;
    wire new_AGEMA_signal_2891 ;
    wire new_AGEMA_signal_2892 ;
    wire new_AGEMA_signal_2893 ;
    wire new_AGEMA_signal_2895 ;
    wire new_AGEMA_signal_2896 ;
    wire new_AGEMA_signal_2897 ;
    wire new_AGEMA_signal_2898 ;
    wire new_AGEMA_signal_2899 ;
    wire new_AGEMA_signal_2901 ;
    wire new_AGEMA_signal_2902 ;
    wire new_AGEMA_signal_2903 ;
    wire new_AGEMA_signal_2904 ;
    wire new_AGEMA_signal_2905 ;
    wire new_AGEMA_signal_2907 ;
    wire new_AGEMA_signal_2908 ;
    wire new_AGEMA_signal_2909 ;
    wire new_AGEMA_signal_2910 ;
    wire new_AGEMA_signal_2911 ;
    wire new_AGEMA_signal_2913 ;
    wire new_AGEMA_signal_2914 ;
    wire new_AGEMA_signal_2915 ;
    wire new_AGEMA_signal_2916 ;
    wire new_AGEMA_signal_2917 ;
    wire new_AGEMA_signal_2919 ;
    wire new_AGEMA_signal_2920 ;
    wire new_AGEMA_signal_2921 ;
    wire new_AGEMA_signal_2922 ;
    wire new_AGEMA_signal_2923 ;
    wire new_AGEMA_signal_2924 ;
    wire new_AGEMA_signal_2925 ;
    wire new_AGEMA_signal_2926 ;
    wire new_AGEMA_signal_2927 ;
    wire new_AGEMA_signal_2928 ;
    wire new_AGEMA_signal_2929 ;
    wire new_AGEMA_signal_2930 ;
    wire new_AGEMA_signal_2931 ;
    wire new_AGEMA_signal_2932 ;
    wire new_AGEMA_signal_2933 ;
    wire new_AGEMA_signal_2934 ;
    wire new_AGEMA_signal_2935 ;
    wire new_AGEMA_signal_2936 ;
    wire new_AGEMA_signal_2937 ;
    wire new_AGEMA_signal_2938 ;
    wire new_AGEMA_signal_2939 ;
    wire new_AGEMA_signal_2940 ;
    wire new_AGEMA_signal_2941 ;
    wire new_AGEMA_signal_2942 ;
    wire new_AGEMA_signal_2943 ;
    wire new_AGEMA_signal_2944 ;
    wire new_AGEMA_signal_2945 ;
    wire new_AGEMA_signal_2946 ;
    wire new_AGEMA_signal_2947 ;
    wire new_AGEMA_signal_2948 ;
    wire new_AGEMA_signal_2949 ;
    wire new_AGEMA_signal_2950 ;
    wire new_AGEMA_signal_2951 ;
    wire new_AGEMA_signal_2952 ;
    wire new_AGEMA_signal_2953 ;
    wire new_AGEMA_signal_2954 ;
    wire new_AGEMA_signal_2955 ;
    wire new_AGEMA_signal_2956 ;
    wire new_AGEMA_signal_2957 ;
    wire new_AGEMA_signal_2958 ;
    wire new_AGEMA_signal_2959 ;
    wire new_AGEMA_signal_2960 ;
    wire new_AGEMA_signal_2961 ;
    wire new_AGEMA_signal_2962 ;
    wire new_AGEMA_signal_2963 ;
    wire new_AGEMA_signal_2964 ;
    wire new_AGEMA_signal_2965 ;
    wire new_AGEMA_signal_2966 ;
    wire new_AGEMA_signal_2967 ;
    wire new_AGEMA_signal_2968 ;
    wire new_AGEMA_signal_2969 ;
    wire new_AGEMA_signal_2970 ;
    wire new_AGEMA_signal_2971 ;
    wire new_AGEMA_signal_2972 ;
    wire new_AGEMA_signal_2973 ;
    wire new_AGEMA_signal_2974 ;
    wire new_AGEMA_signal_2975 ;
    wire new_AGEMA_signal_2976 ;
    wire new_AGEMA_signal_2977 ;
    wire new_AGEMA_signal_2978 ;
    wire new_AGEMA_signal_2979 ;
    wire new_AGEMA_signal_2980 ;
    wire new_AGEMA_signal_2981 ;
    wire new_AGEMA_signal_2982 ;
    wire new_AGEMA_signal_2983 ;
    wire new_AGEMA_signal_2984 ;
    wire new_AGEMA_signal_2985 ;
    wire new_AGEMA_signal_2986 ;
    wire new_AGEMA_signal_2987 ;
    wire new_AGEMA_signal_2988 ;
    wire new_AGEMA_signal_2989 ;
    wire new_AGEMA_signal_2990 ;
    wire new_AGEMA_signal_2991 ;
    wire new_AGEMA_signal_2992 ;
    wire new_AGEMA_signal_2993 ;
    wire new_AGEMA_signal_2994 ;
    wire new_AGEMA_signal_2995 ;
    wire new_AGEMA_signal_2996 ;
    wire new_AGEMA_signal_2997 ;
    wire new_AGEMA_signal_2998 ;
    wire new_AGEMA_signal_2999 ;
    wire new_AGEMA_signal_3000 ;
    wire new_AGEMA_signal_3001 ;
    wire new_AGEMA_signal_3002 ;
    wire new_AGEMA_signal_3003 ;
    wire new_AGEMA_signal_3004 ;
    wire new_AGEMA_signal_3005 ;
    wire new_AGEMA_signal_3006 ;
    wire new_AGEMA_signal_3007 ;
    wire new_AGEMA_signal_3008 ;
    wire new_AGEMA_signal_3009 ;
    wire new_AGEMA_signal_3010 ;
    wire new_AGEMA_signal_3011 ;
    wire new_AGEMA_signal_3012 ;
    wire new_AGEMA_signal_3013 ;
    wire new_AGEMA_signal_3014 ;
    wire new_AGEMA_signal_3015 ;
    wire new_AGEMA_signal_3016 ;
    wire new_AGEMA_signal_3017 ;
    wire new_AGEMA_signal_3018 ;
    wire new_AGEMA_signal_3019 ;
    wire new_AGEMA_signal_3020 ;
    wire new_AGEMA_signal_3021 ;
    wire new_AGEMA_signal_3022 ;
    wire new_AGEMA_signal_3023 ;
    wire new_AGEMA_signal_3024 ;
    wire new_AGEMA_signal_3025 ;
    wire new_AGEMA_signal_3026 ;
    wire new_AGEMA_signal_3027 ;
    wire new_AGEMA_signal_3028 ;
    wire new_AGEMA_signal_3029 ;
    wire new_AGEMA_signal_3030 ;
    wire new_AGEMA_signal_3031 ;
    wire new_AGEMA_signal_3032 ;
    wire new_AGEMA_signal_3033 ;
    wire new_AGEMA_signal_3034 ;
    wire new_AGEMA_signal_3035 ;
    wire new_AGEMA_signal_3036 ;
    wire new_AGEMA_signal_3037 ;
    wire new_AGEMA_signal_3038 ;
    wire new_AGEMA_signal_3039 ;
    wire new_AGEMA_signal_3040 ;
    wire new_AGEMA_signal_3041 ;
    wire new_AGEMA_signal_3042 ;
    wire new_AGEMA_signal_3043 ;
    wire new_AGEMA_signal_3044 ;
    wire new_AGEMA_signal_3045 ;
    wire new_AGEMA_signal_3046 ;
    wire new_AGEMA_signal_3047 ;
    wire new_AGEMA_signal_3048 ;
    wire new_AGEMA_signal_3049 ;
    wire new_AGEMA_signal_3050 ;
    wire new_AGEMA_signal_3051 ;
    wire new_AGEMA_signal_3052 ;
    wire new_AGEMA_signal_3053 ;
    wire new_AGEMA_signal_3054 ;
    wire new_AGEMA_signal_3055 ;
    wire new_AGEMA_signal_3056 ;
    wire new_AGEMA_signal_3057 ;
    wire new_AGEMA_signal_3058 ;
    wire new_AGEMA_signal_3059 ;
    wire new_AGEMA_signal_3060 ;
    wire new_AGEMA_signal_3061 ;
    wire new_AGEMA_signal_3062 ;
    wire new_AGEMA_signal_3063 ;
    wire new_AGEMA_signal_3064 ;
    wire new_AGEMA_signal_3065 ;
    wire new_AGEMA_signal_3066 ;
    wire new_AGEMA_signal_3067 ;
    wire new_AGEMA_signal_3068 ;
    wire new_AGEMA_signal_3069 ;
    wire new_AGEMA_signal_3070 ;
    wire new_AGEMA_signal_3071 ;
    wire new_AGEMA_signal_3072 ;
    wire new_AGEMA_signal_3073 ;
    wire new_AGEMA_signal_3074 ;
    wire new_AGEMA_signal_3075 ;
    wire new_AGEMA_signal_3076 ;
    wire new_AGEMA_signal_3077 ;
    wire new_AGEMA_signal_3078 ;
    wire new_AGEMA_signal_3079 ;
    wire new_AGEMA_signal_3080 ;
    wire new_AGEMA_signal_3081 ;
    wire new_AGEMA_signal_3082 ;
    wire new_AGEMA_signal_3083 ;
    wire new_AGEMA_signal_3084 ;
    wire new_AGEMA_signal_3085 ;
    wire new_AGEMA_signal_3086 ;
    wire new_AGEMA_signal_3087 ;
    wire new_AGEMA_signal_3088 ;
    wire new_AGEMA_signal_3089 ;
    wire new_AGEMA_signal_3090 ;
    wire new_AGEMA_signal_3091 ;
    wire new_AGEMA_signal_3092 ;
    wire new_AGEMA_signal_3093 ;
    wire new_AGEMA_signal_3094 ;
    wire new_AGEMA_signal_3095 ;
    wire new_AGEMA_signal_3096 ;
    wire new_AGEMA_signal_3097 ;
    wire new_AGEMA_signal_3098 ;
    wire new_AGEMA_signal_3099 ;
    wire new_AGEMA_signal_3100 ;
    wire new_AGEMA_signal_3101 ;
    wire new_AGEMA_signal_3102 ;
    wire new_AGEMA_signal_3103 ;
    wire new_AGEMA_signal_3104 ;
    wire new_AGEMA_signal_3105 ;
    wire new_AGEMA_signal_3106 ;
    wire new_AGEMA_signal_3107 ;
    wire new_AGEMA_signal_3108 ;
    wire new_AGEMA_signal_3109 ;
    wire new_AGEMA_signal_3110 ;
    wire new_AGEMA_signal_3111 ;
    wire new_AGEMA_signal_3112 ;
    wire new_AGEMA_signal_3113 ;
    wire new_AGEMA_signal_3114 ;
    wire new_AGEMA_signal_3115 ;
    wire new_AGEMA_signal_3116 ;
    wire new_AGEMA_signal_3117 ;
    wire new_AGEMA_signal_3118 ;
    wire new_AGEMA_signal_3119 ;
    wire new_AGEMA_signal_3120 ;
    wire new_AGEMA_signal_3121 ;
    wire new_AGEMA_signal_3122 ;
    wire new_AGEMA_signal_3123 ;
    wire new_AGEMA_signal_3124 ;
    wire new_AGEMA_signal_3125 ;
    wire new_AGEMA_signal_3126 ;
    wire new_AGEMA_signal_3127 ;
    wire new_AGEMA_signal_3128 ;
    wire new_AGEMA_signal_3129 ;
    wire new_AGEMA_signal_3130 ;
    wire new_AGEMA_signal_3131 ;
    wire new_AGEMA_signal_3132 ;
    wire new_AGEMA_signal_3133 ;
    wire new_AGEMA_signal_3134 ;
    wire new_AGEMA_signal_3135 ;
    wire new_AGEMA_signal_3136 ;
    wire new_AGEMA_signal_3137 ;
    wire new_AGEMA_signal_3138 ;
    wire new_AGEMA_signal_3139 ;
    wire new_AGEMA_signal_3140 ;
    wire new_AGEMA_signal_3141 ;
    wire new_AGEMA_signal_3142 ;
    wire new_AGEMA_signal_3143 ;
    wire new_AGEMA_signal_3144 ;
    wire new_AGEMA_signal_3145 ;
    wire new_AGEMA_signal_3146 ;
    wire new_AGEMA_signal_3147 ;
    wire new_AGEMA_signal_3148 ;
    wire new_AGEMA_signal_3149 ;
    wire new_AGEMA_signal_3150 ;
    wire new_AGEMA_signal_3151 ;
    wire new_AGEMA_signal_3152 ;
    wire new_AGEMA_signal_3153 ;
    wire new_AGEMA_signal_3154 ;
    wire new_AGEMA_signal_3155 ;
    wire new_AGEMA_signal_3156 ;
    wire new_AGEMA_signal_3157 ;
    wire new_AGEMA_signal_3158 ;
    wire new_AGEMA_signal_3159 ;
    wire new_AGEMA_signal_3160 ;
    wire new_AGEMA_signal_3161 ;
    wire new_AGEMA_signal_3162 ;
    wire new_AGEMA_signal_3163 ;
    wire new_AGEMA_signal_3164 ;
    wire new_AGEMA_signal_3165 ;
    wire new_AGEMA_signal_3166 ;
    wire new_AGEMA_signal_3167 ;
    wire new_AGEMA_signal_3168 ;
    wire new_AGEMA_signal_3169 ;
    wire new_AGEMA_signal_3170 ;
    wire new_AGEMA_signal_3171 ;
    wire new_AGEMA_signal_3172 ;
    wire new_AGEMA_signal_3173 ;
    wire new_AGEMA_signal_3174 ;
    wire new_AGEMA_signal_3175 ;
    wire new_AGEMA_signal_3176 ;
    wire new_AGEMA_signal_3177 ;
    wire new_AGEMA_signal_3178 ;
    wire new_AGEMA_signal_3179 ;
    wire new_AGEMA_signal_3180 ;
    wire new_AGEMA_signal_3181 ;
    wire new_AGEMA_signal_3182 ;
    wire new_AGEMA_signal_3183 ;
    wire new_AGEMA_signal_3184 ;
    wire new_AGEMA_signal_3185 ;
    wire new_AGEMA_signal_3186 ;
    wire new_AGEMA_signal_3187 ;
    wire new_AGEMA_signal_3188 ;
    wire new_AGEMA_signal_3189 ;
    wire new_AGEMA_signal_3190 ;
    wire new_AGEMA_signal_3191 ;
    wire new_AGEMA_signal_3192 ;
    wire new_AGEMA_signal_3193 ;
    wire new_AGEMA_signal_3194 ;
    wire new_AGEMA_signal_3195 ;
    wire new_AGEMA_signal_3196 ;
    wire new_AGEMA_signal_3197 ;
    wire new_AGEMA_signal_3198 ;
    wire new_AGEMA_signal_3199 ;
    wire new_AGEMA_signal_3200 ;
    wire new_AGEMA_signal_3201 ;
    wire new_AGEMA_signal_3202 ;
    wire new_AGEMA_signal_3203 ;
    wire new_AGEMA_signal_3204 ;
    wire new_AGEMA_signal_3205 ;
    wire new_AGEMA_signal_3206 ;
    wire new_AGEMA_signal_3207 ;
    wire new_AGEMA_signal_3208 ;
    wire new_AGEMA_signal_3209 ;
    wire new_AGEMA_signal_3210 ;
    wire new_AGEMA_signal_3211 ;
    wire new_AGEMA_signal_3212 ;
    wire new_AGEMA_signal_3213 ;
    wire new_AGEMA_signal_3214 ;
    wire new_AGEMA_signal_3215 ;
    wire new_AGEMA_signal_3216 ;
    wire new_AGEMA_signal_3217 ;
    wire new_AGEMA_signal_3218 ;
    wire new_AGEMA_signal_3219 ;
    wire new_AGEMA_signal_3220 ;
    wire new_AGEMA_signal_3221 ;
    wire new_AGEMA_signal_3222 ;
    wire new_AGEMA_signal_3223 ;
    wire new_AGEMA_signal_3224 ;
    wire new_AGEMA_signal_3225 ;
    wire new_AGEMA_signal_3226 ;
    wire new_AGEMA_signal_3227 ;
    wire new_AGEMA_signal_3228 ;
    wire new_AGEMA_signal_3229 ;
    wire new_AGEMA_signal_3230 ;
    wire new_AGEMA_signal_3231 ;
    wire new_AGEMA_signal_3232 ;
    wire new_AGEMA_signal_3233 ;
    wire new_AGEMA_signal_3234 ;
    wire new_AGEMA_signal_3235 ;
    wire new_AGEMA_signal_3236 ;
    wire new_AGEMA_signal_3237 ;
    wire new_AGEMA_signal_3238 ;
    wire new_AGEMA_signal_3239 ;
    wire new_AGEMA_signal_3240 ;
    wire new_AGEMA_signal_3241 ;
    wire new_AGEMA_signal_3242 ;
    wire new_AGEMA_signal_3243 ;
    wire new_AGEMA_signal_3244 ;
    wire new_AGEMA_signal_3245 ;
    wire new_AGEMA_signal_3246 ;
    wire new_AGEMA_signal_3247 ;
    wire new_AGEMA_signal_3248 ;
    wire new_AGEMA_signal_3249 ;
    wire new_AGEMA_signal_3250 ;
    wire new_AGEMA_signal_3251 ;
    wire new_AGEMA_signal_3252 ;
    wire new_AGEMA_signal_3253 ;
    wire new_AGEMA_signal_3254 ;
    wire new_AGEMA_signal_3255 ;
    wire new_AGEMA_signal_3256 ;
    wire new_AGEMA_signal_3257 ;
    wire new_AGEMA_signal_3258 ;
    wire new_AGEMA_signal_3259 ;
    wire new_AGEMA_signal_3260 ;
    wire new_AGEMA_signal_3261 ;
    wire new_AGEMA_signal_3262 ;
    wire new_AGEMA_signal_3263 ;
    wire new_AGEMA_signal_3264 ;
    wire new_AGEMA_signal_3265 ;
    wire new_AGEMA_signal_3266 ;
    wire new_AGEMA_signal_3267 ;
    wire new_AGEMA_signal_3268 ;
    wire new_AGEMA_signal_3269 ;
    wire new_AGEMA_signal_3270 ;
    wire new_AGEMA_signal_3271 ;
    wire new_AGEMA_signal_3272 ;
    wire new_AGEMA_signal_3273 ;
    wire new_AGEMA_signal_3274 ;
    wire new_AGEMA_signal_3275 ;
    wire new_AGEMA_signal_3276 ;
    wire new_AGEMA_signal_3277 ;
    wire new_AGEMA_signal_3278 ;
    wire new_AGEMA_signal_3279 ;
    wire new_AGEMA_signal_3280 ;
    wire new_AGEMA_signal_3281 ;
    wire new_AGEMA_signal_3282 ;
    wire new_AGEMA_signal_3283 ;
    wire new_AGEMA_signal_3284 ;
    wire new_AGEMA_signal_3285 ;
    wire new_AGEMA_signal_3286 ;
    wire new_AGEMA_signal_3287 ;
    wire new_AGEMA_signal_3288 ;
    wire new_AGEMA_signal_3289 ;
    wire new_AGEMA_signal_3290 ;
    wire new_AGEMA_signal_3291 ;
    wire new_AGEMA_signal_3292 ;
    wire new_AGEMA_signal_3293 ;
    wire new_AGEMA_signal_3294 ;
    wire new_AGEMA_signal_3295 ;
    wire new_AGEMA_signal_3296 ;
    wire new_AGEMA_signal_3297 ;
    wire new_AGEMA_signal_3298 ;
    wire new_AGEMA_signal_3299 ;
    wire new_AGEMA_signal_3300 ;
    wire new_AGEMA_signal_3301 ;
    wire new_AGEMA_signal_3302 ;
    wire new_AGEMA_signal_3303 ;
    wire new_AGEMA_signal_3304 ;
    wire new_AGEMA_signal_3305 ;
    wire new_AGEMA_signal_3306 ;
    wire new_AGEMA_signal_3307 ;
    wire new_AGEMA_signal_3308 ;
    wire new_AGEMA_signal_3309 ;
    wire new_AGEMA_signal_3310 ;
    wire new_AGEMA_signal_3311 ;
    wire new_AGEMA_signal_3312 ;
    wire new_AGEMA_signal_3313 ;
    wire new_AGEMA_signal_3314 ;
    wire new_AGEMA_signal_3315 ;
    wire new_AGEMA_signal_3316 ;
    wire new_AGEMA_signal_3317 ;
    wire new_AGEMA_signal_3318 ;
    wire new_AGEMA_signal_3319 ;
    wire new_AGEMA_signal_3320 ;
    wire new_AGEMA_signal_3321 ;
    wire new_AGEMA_signal_3322 ;
    wire new_AGEMA_signal_3323 ;
    wire new_AGEMA_signal_3324 ;
    wire new_AGEMA_signal_3325 ;
    wire new_AGEMA_signal_3326 ;
    wire new_AGEMA_signal_3327 ;
    wire new_AGEMA_signal_3328 ;
    wire new_AGEMA_signal_3329 ;
    wire new_AGEMA_signal_3330 ;
    wire new_AGEMA_signal_3331 ;
    wire new_AGEMA_signal_3332 ;
    wire new_AGEMA_signal_3333 ;
    wire new_AGEMA_signal_3334 ;
    wire new_AGEMA_signal_3335 ;
    wire new_AGEMA_signal_3336 ;
    wire new_AGEMA_signal_3337 ;
    wire new_AGEMA_signal_3338 ;
    wire new_AGEMA_signal_3339 ;
    wire new_AGEMA_signal_3340 ;
    wire new_AGEMA_signal_3341 ;
    wire new_AGEMA_signal_3342 ;
    wire new_AGEMA_signal_3343 ;
    wire new_AGEMA_signal_3344 ;
    wire new_AGEMA_signal_3345 ;
    wire new_AGEMA_signal_3346 ;
    wire new_AGEMA_signal_3347 ;
    wire new_AGEMA_signal_3348 ;
    wire new_AGEMA_signal_3349 ;
    wire new_AGEMA_signal_3350 ;
    wire new_AGEMA_signal_3351 ;
    wire new_AGEMA_signal_3352 ;
    wire new_AGEMA_signal_3353 ;
    wire new_AGEMA_signal_3354 ;
    wire new_AGEMA_signal_3355 ;
    wire new_AGEMA_signal_3356 ;
    wire new_AGEMA_signal_3357 ;
    wire new_AGEMA_signal_3358 ;
    wire new_AGEMA_signal_3359 ;
    wire new_AGEMA_signal_3360 ;
    wire new_AGEMA_signal_3361 ;
    wire new_AGEMA_signal_3362 ;
    wire new_AGEMA_signal_3363 ;
    wire new_AGEMA_signal_3364 ;
    wire new_AGEMA_signal_3365 ;
    wire new_AGEMA_signal_3366 ;
    wire new_AGEMA_signal_3367 ;
    wire new_AGEMA_signal_3368 ;
    wire new_AGEMA_signal_3369 ;
    wire new_AGEMA_signal_3370 ;
    wire new_AGEMA_signal_3371 ;
    wire new_AGEMA_signal_3372 ;
    wire new_AGEMA_signal_3373 ;
    wire new_AGEMA_signal_3374 ;
    wire new_AGEMA_signal_3375 ;
    wire new_AGEMA_signal_3376 ;
    wire new_AGEMA_signal_3377 ;
    wire new_AGEMA_signal_3378 ;
    wire new_AGEMA_signal_3379 ;
    wire new_AGEMA_signal_3380 ;
    wire new_AGEMA_signal_3381 ;
    wire new_AGEMA_signal_3382 ;
    wire new_AGEMA_signal_3383 ;
    wire new_AGEMA_signal_3384 ;
    wire new_AGEMA_signal_3385 ;
    wire new_AGEMA_signal_3386 ;
    wire new_AGEMA_signal_3387 ;
    wire new_AGEMA_signal_3388 ;
    wire new_AGEMA_signal_3389 ;
    wire new_AGEMA_signal_3390 ;
    wire new_AGEMA_signal_3391 ;
    wire new_AGEMA_signal_3392 ;
    wire new_AGEMA_signal_3393 ;
    wire new_AGEMA_signal_3394 ;
    wire new_AGEMA_signal_3395 ;
    wire new_AGEMA_signal_3396 ;
    wire new_AGEMA_signal_3397 ;
    wire new_AGEMA_signal_3398 ;
    wire new_AGEMA_signal_3399 ;
    wire new_AGEMA_signal_3400 ;
    wire new_AGEMA_signal_3401 ;
    wire new_AGEMA_signal_3402 ;
    wire new_AGEMA_signal_3403 ;
    wire new_AGEMA_signal_3404 ;
    wire new_AGEMA_signal_3405 ;
    wire new_AGEMA_signal_3406 ;
    wire new_AGEMA_signal_3407 ;
    wire new_AGEMA_signal_3408 ;
    wire new_AGEMA_signal_3409 ;
    wire new_AGEMA_signal_3410 ;
    wire new_AGEMA_signal_3411 ;
    wire new_AGEMA_signal_3412 ;
    wire new_AGEMA_signal_3413 ;
    wire new_AGEMA_signal_3414 ;
    wire new_AGEMA_signal_3415 ;
    wire new_AGEMA_signal_3416 ;
    wire new_AGEMA_signal_3417 ;
    wire new_AGEMA_signal_3418 ;
    wire new_AGEMA_signal_3419 ;
    wire new_AGEMA_signal_3420 ;
    wire new_AGEMA_signal_3421 ;
    wire new_AGEMA_signal_3422 ;
    wire new_AGEMA_signal_3423 ;
    wire new_AGEMA_signal_3424 ;
    wire new_AGEMA_signal_3425 ;
    wire new_AGEMA_signal_3426 ;
    wire new_AGEMA_signal_3427 ;
    wire new_AGEMA_signal_3428 ;
    wire new_AGEMA_signal_3429 ;
    wire new_AGEMA_signal_3430 ;
    wire new_AGEMA_signal_3431 ;
    wire new_AGEMA_signal_3432 ;
    wire new_AGEMA_signal_3433 ;
    wire new_AGEMA_signal_3434 ;
    wire new_AGEMA_signal_3435 ;
    wire new_AGEMA_signal_3436 ;
    wire new_AGEMA_signal_3437 ;
    wire new_AGEMA_signal_3438 ;
    wire new_AGEMA_signal_3439 ;
    wire new_AGEMA_signal_3440 ;
    wire new_AGEMA_signal_3441 ;
    wire new_AGEMA_signal_3442 ;
    wire new_AGEMA_signal_3443 ;
    wire new_AGEMA_signal_3444 ;
    wire new_AGEMA_signal_3445 ;
    wire new_AGEMA_signal_3446 ;
    wire new_AGEMA_signal_3447 ;
    wire new_AGEMA_signal_3448 ;
    wire new_AGEMA_signal_3449 ;
    wire new_AGEMA_signal_3450 ;
    wire new_AGEMA_signal_3451 ;
    wire new_AGEMA_signal_3452 ;
    wire new_AGEMA_signal_3453 ;
    wire new_AGEMA_signal_3454 ;
    wire new_AGEMA_signal_3455 ;
    wire new_AGEMA_signal_3456 ;
    wire new_AGEMA_signal_3457 ;
    wire new_AGEMA_signal_3458 ;
    wire new_AGEMA_signal_3459 ;
    wire new_AGEMA_signal_3460 ;
    wire new_AGEMA_signal_3461 ;
    wire new_AGEMA_signal_3462 ;
    wire new_AGEMA_signal_3463 ;
    wire new_AGEMA_signal_3464 ;
    wire new_AGEMA_signal_3465 ;
    wire new_AGEMA_signal_3466 ;
    wire new_AGEMA_signal_3467 ;
    wire new_AGEMA_signal_3468 ;
    wire new_AGEMA_signal_3469 ;
    wire new_AGEMA_signal_3470 ;
    wire new_AGEMA_signal_3471 ;
    wire new_AGEMA_signal_3472 ;
    wire new_AGEMA_signal_3473 ;
    wire new_AGEMA_signal_3474 ;
    wire new_AGEMA_signal_3475 ;
    wire new_AGEMA_signal_3476 ;
    wire new_AGEMA_signal_3477 ;
    wire new_AGEMA_signal_3478 ;
    wire new_AGEMA_signal_3479 ;
    wire new_AGEMA_signal_3480 ;
    wire new_AGEMA_signal_3481 ;
    wire new_AGEMA_signal_3482 ;
    wire new_AGEMA_signal_3483 ;
    wire new_AGEMA_signal_3484 ;
    wire new_AGEMA_signal_3485 ;
    wire new_AGEMA_signal_3486 ;
    wire new_AGEMA_signal_3487 ;
    wire new_AGEMA_signal_3488 ;
    wire new_AGEMA_signal_3489 ;
    wire new_AGEMA_signal_3490 ;
    wire new_AGEMA_signal_3491 ;
    wire new_AGEMA_signal_3492 ;
    wire new_AGEMA_signal_3493 ;
    wire new_AGEMA_signal_3494 ;
    wire new_AGEMA_signal_3495 ;
    wire new_AGEMA_signal_3496 ;
    wire new_AGEMA_signal_3497 ;
    wire new_AGEMA_signal_3498 ;
    wire new_AGEMA_signal_3499 ;
    wire new_AGEMA_signal_3500 ;
    wire new_AGEMA_signal_3501 ;
    wire new_AGEMA_signal_3502 ;
    wire new_AGEMA_signal_3503 ;
    wire new_AGEMA_signal_3504 ;
    wire new_AGEMA_signal_3505 ;
    wire new_AGEMA_signal_3506 ;
    wire new_AGEMA_signal_3507 ;
    wire new_AGEMA_signal_3508 ;
    wire new_AGEMA_signal_3509 ;
    wire new_AGEMA_signal_3510 ;
    wire new_AGEMA_signal_3511 ;
    wire new_AGEMA_signal_3512 ;
    wire new_AGEMA_signal_3513 ;
    wire new_AGEMA_signal_3514 ;
    wire new_AGEMA_signal_3515 ;
    wire new_AGEMA_signal_3516 ;
    wire new_AGEMA_signal_3517 ;
    wire new_AGEMA_signal_3518 ;
    wire new_AGEMA_signal_3519 ;
    wire new_AGEMA_signal_3520 ;
    wire new_AGEMA_signal_3521 ;
    wire new_AGEMA_signal_3522 ;
    wire new_AGEMA_signal_3523 ;
    wire new_AGEMA_signal_3524 ;
    wire new_AGEMA_signal_3525 ;
    wire new_AGEMA_signal_3526 ;
    wire new_AGEMA_signal_3527 ;
    wire new_AGEMA_signal_3528 ;
    wire new_AGEMA_signal_3529 ;
    wire new_AGEMA_signal_3530 ;
    wire new_AGEMA_signal_3531 ;
    wire new_AGEMA_signal_3532 ;
    wire new_AGEMA_signal_3533 ;
    wire new_AGEMA_signal_3534 ;
    wire new_AGEMA_signal_3535 ;
    wire new_AGEMA_signal_3536 ;
    wire new_AGEMA_signal_3537 ;
    wire new_AGEMA_signal_3538 ;
    wire new_AGEMA_signal_3539 ;
    wire new_AGEMA_signal_3540 ;
    wire new_AGEMA_signal_3541 ;
    wire new_AGEMA_signal_3542 ;
    wire new_AGEMA_signal_3543 ;
    wire new_AGEMA_signal_3544 ;
    wire new_AGEMA_signal_3545 ;
    wire new_AGEMA_signal_3546 ;
    wire new_AGEMA_signal_3547 ;
    wire new_AGEMA_signal_3548 ;
    wire new_AGEMA_signal_3549 ;
    wire new_AGEMA_signal_3550 ;
    wire new_AGEMA_signal_3551 ;
    wire new_AGEMA_signal_3552 ;
    wire new_AGEMA_signal_3553 ;
    wire new_AGEMA_signal_3554 ;
    wire new_AGEMA_signal_3555 ;
    wire new_AGEMA_signal_3556 ;
    wire new_AGEMA_signal_3557 ;
    wire new_AGEMA_signal_3558 ;
    wire new_AGEMA_signal_3559 ;
    wire new_AGEMA_signal_3560 ;
    wire new_AGEMA_signal_3561 ;
    wire new_AGEMA_signal_3562 ;
    wire new_AGEMA_signal_3563 ;
    wire new_AGEMA_signal_3564 ;
    wire new_AGEMA_signal_3565 ;
    wire new_AGEMA_signal_3566 ;
    wire new_AGEMA_signal_3567 ;
    wire new_AGEMA_signal_3568 ;
    wire new_AGEMA_signal_3569 ;
    wire new_AGEMA_signal_3570 ;
    wire new_AGEMA_signal_3571 ;
    wire new_AGEMA_signal_3572 ;
    wire new_AGEMA_signal_3573 ;
    wire new_AGEMA_signal_3574 ;
    wire new_AGEMA_signal_3575 ;
    wire new_AGEMA_signal_3576 ;
    wire new_AGEMA_signal_3577 ;
    wire new_AGEMA_signal_3578 ;
    wire new_AGEMA_signal_3579 ;
    wire new_AGEMA_signal_3580 ;
    wire new_AGEMA_signal_3581 ;
    wire new_AGEMA_signal_3582 ;
    wire new_AGEMA_signal_3583 ;
    wire new_AGEMA_signal_3584 ;
    wire new_AGEMA_signal_3585 ;
    wire new_AGEMA_signal_3586 ;
    wire new_AGEMA_signal_3587 ;
    wire new_AGEMA_signal_3588 ;
    wire new_AGEMA_signal_3589 ;
    wire new_AGEMA_signal_3590 ;
    wire new_AGEMA_signal_3591 ;
    wire new_AGEMA_signal_3592 ;
    wire new_AGEMA_signal_3593 ;
    wire new_AGEMA_signal_3594 ;
    wire new_AGEMA_signal_3595 ;
    wire new_AGEMA_signal_3596 ;
    wire new_AGEMA_signal_3597 ;
    wire new_AGEMA_signal_3598 ;
    wire new_AGEMA_signal_3599 ;
    wire new_AGEMA_signal_3600 ;
    wire new_AGEMA_signal_3601 ;
    wire new_AGEMA_signal_3602 ;
    wire new_AGEMA_signal_3603 ;
    wire new_AGEMA_signal_3604 ;
    wire new_AGEMA_signal_3605 ;
    wire new_AGEMA_signal_3606 ;
    wire new_AGEMA_signal_3607 ;
    wire new_AGEMA_signal_3608 ;
    wire new_AGEMA_signal_3609 ;
    wire new_AGEMA_signal_3610 ;
    wire new_AGEMA_signal_3611 ;
    wire new_AGEMA_signal_3612 ;
    wire new_AGEMA_signal_3613 ;
    wire new_AGEMA_signal_3614 ;
    wire new_AGEMA_signal_3615 ;
    wire new_AGEMA_signal_3616 ;
    wire new_AGEMA_signal_3617 ;
    wire new_AGEMA_signal_3618 ;
    wire new_AGEMA_signal_3619 ;
    wire new_AGEMA_signal_3620 ;
    wire new_AGEMA_signal_3621 ;
    wire new_AGEMA_signal_3622 ;
    wire new_AGEMA_signal_3623 ;
    wire new_AGEMA_signal_3624 ;
    wire new_AGEMA_signal_3625 ;
    wire new_AGEMA_signal_3626 ;
    wire new_AGEMA_signal_3627 ;
    wire new_AGEMA_signal_3628 ;
    wire new_AGEMA_signal_3629 ;
    wire new_AGEMA_signal_3630 ;
    wire new_AGEMA_signal_3631 ;
    wire new_AGEMA_signal_3632 ;
    wire new_AGEMA_signal_3633 ;
    wire new_AGEMA_signal_3634 ;
    wire new_AGEMA_signal_3635 ;
    wire new_AGEMA_signal_3636 ;
    wire new_AGEMA_signal_3637 ;
    wire new_AGEMA_signal_3638 ;
    wire new_AGEMA_signal_3639 ;
    wire new_AGEMA_signal_3640 ;
    wire new_AGEMA_signal_3641 ;
    wire new_AGEMA_signal_3642 ;
    wire new_AGEMA_signal_3643 ;
    wire new_AGEMA_signal_3644 ;
    wire new_AGEMA_signal_3645 ;
    wire new_AGEMA_signal_3646 ;
    wire new_AGEMA_signal_3647 ;
    wire new_AGEMA_signal_3648 ;
    wire new_AGEMA_signal_3649 ;
    wire new_AGEMA_signal_3650 ;
    wire new_AGEMA_signal_3651 ;
    wire new_AGEMA_signal_3652 ;
    wire new_AGEMA_signal_3653 ;
    wire new_AGEMA_signal_3654 ;
    wire new_AGEMA_signal_3655 ;
    wire new_AGEMA_signal_3656 ;
    wire new_AGEMA_signal_3657 ;
    wire new_AGEMA_signal_3658 ;
    wire new_AGEMA_signal_3659 ;
    wire new_AGEMA_signal_3660 ;
    wire new_AGEMA_signal_3661 ;
    wire new_AGEMA_signal_3662 ;
    wire new_AGEMA_signal_3663 ;
    wire new_AGEMA_signal_3664 ;
    wire new_AGEMA_signal_3665 ;
    wire new_AGEMA_signal_3666 ;
    wire new_AGEMA_signal_3667 ;
    wire new_AGEMA_signal_3668 ;
    wire new_AGEMA_signal_3669 ;
    wire new_AGEMA_signal_3670 ;
    wire new_AGEMA_signal_3671 ;
    wire new_AGEMA_signal_3672 ;
    wire new_AGEMA_signal_3673 ;
    wire new_AGEMA_signal_3674 ;
    wire new_AGEMA_signal_3675 ;
    wire new_AGEMA_signal_3676 ;
    wire new_AGEMA_signal_3677 ;
    wire new_AGEMA_signal_3678 ;
    wire new_AGEMA_signal_3679 ;
    wire new_AGEMA_signal_3680 ;
    wire new_AGEMA_signal_3681 ;
    wire new_AGEMA_signal_3682 ;
    wire new_AGEMA_signal_3683 ;
    wire new_AGEMA_signal_3684 ;
    wire new_AGEMA_signal_3685 ;
    wire new_AGEMA_signal_3686 ;
    wire new_AGEMA_signal_3687 ;
    wire new_AGEMA_signal_3688 ;
    wire new_AGEMA_signal_3689 ;
    wire new_AGEMA_signal_3690 ;
    wire new_AGEMA_signal_3691 ;
    wire new_AGEMA_signal_3692 ;
    wire new_AGEMA_signal_3693 ;
    wire new_AGEMA_signal_3694 ;
    wire new_AGEMA_signal_3695 ;
    wire new_AGEMA_signal_3696 ;
    wire new_AGEMA_signal_3697 ;
    wire new_AGEMA_signal_3698 ;
    wire new_AGEMA_signal_3699 ;
    wire new_AGEMA_signal_3700 ;
    wire new_AGEMA_signal_3701 ;
    wire new_AGEMA_signal_3702 ;
    wire new_AGEMA_signal_3703 ;
    wire new_AGEMA_signal_3704 ;
    wire new_AGEMA_signal_3705 ;
    wire new_AGEMA_signal_3706 ;
    wire new_AGEMA_signal_3707 ;
    wire new_AGEMA_signal_3708 ;
    wire new_AGEMA_signal_3709 ;
    wire new_AGEMA_signal_3710 ;
    wire new_AGEMA_signal_3711 ;
    wire new_AGEMA_signal_3712 ;
    wire new_AGEMA_signal_3713 ;
    wire new_AGEMA_signal_3714 ;
    wire new_AGEMA_signal_3715 ;
    wire new_AGEMA_signal_3716 ;
    wire new_AGEMA_signal_3717 ;
    wire new_AGEMA_signal_3718 ;
    wire new_AGEMA_signal_3719 ;
    wire new_AGEMA_signal_3720 ;
    wire new_AGEMA_signal_3721 ;
    wire new_AGEMA_signal_3722 ;
    wire new_AGEMA_signal_3723 ;
    wire new_AGEMA_signal_3724 ;
    wire new_AGEMA_signal_3725 ;
    wire new_AGEMA_signal_3726 ;
    wire new_AGEMA_signal_3727 ;
    wire new_AGEMA_signal_3728 ;
    wire new_AGEMA_signal_3729 ;
    wire new_AGEMA_signal_3730 ;
    wire new_AGEMA_signal_3731 ;
    wire new_AGEMA_signal_3732 ;
    wire new_AGEMA_signal_3733 ;
    wire new_AGEMA_signal_3734 ;
    wire new_AGEMA_signal_3735 ;
    wire new_AGEMA_signal_3736 ;
    wire new_AGEMA_signal_3737 ;
    wire new_AGEMA_signal_3738 ;
    wire new_AGEMA_signal_3739 ;
    wire new_AGEMA_signal_3740 ;
    wire new_AGEMA_signal_3741 ;
    wire new_AGEMA_signal_3742 ;
    wire new_AGEMA_signal_3743 ;
    wire new_AGEMA_signal_3744 ;
    wire new_AGEMA_signal_3745 ;
    wire new_AGEMA_signal_3746 ;
    wire new_AGEMA_signal_3747 ;
    wire new_AGEMA_signal_3748 ;
    wire new_AGEMA_signal_3749 ;
    wire new_AGEMA_signal_3750 ;
    wire new_AGEMA_signal_3751 ;
    wire new_AGEMA_signal_3752 ;
    wire new_AGEMA_signal_3753 ;
    wire new_AGEMA_signal_3754 ;
    wire new_AGEMA_signal_3755 ;
    wire new_AGEMA_signal_3756 ;
    wire new_AGEMA_signal_3757 ;
    wire new_AGEMA_signal_3758 ;
    wire new_AGEMA_signal_3759 ;
    wire new_AGEMA_signal_3760 ;
    wire new_AGEMA_signal_3761 ;
    wire new_AGEMA_signal_3762 ;
    wire new_AGEMA_signal_3763 ;
    wire new_AGEMA_signal_3764 ;
    wire new_AGEMA_signal_3765 ;
    wire new_AGEMA_signal_3766 ;
    wire new_AGEMA_signal_3767 ;
    wire new_AGEMA_signal_3768 ;
    wire new_AGEMA_signal_3769 ;
    wire new_AGEMA_signal_3770 ;
    wire new_AGEMA_signal_3771 ;
    wire new_AGEMA_signal_3772 ;
    wire new_AGEMA_signal_3773 ;
    wire new_AGEMA_signal_3774 ;
    wire new_AGEMA_signal_3775 ;
    wire new_AGEMA_signal_3776 ;
    wire new_AGEMA_signal_3777 ;
    wire new_AGEMA_signal_3778 ;
    wire new_AGEMA_signal_3779 ;
    wire new_AGEMA_signal_3780 ;
    wire new_AGEMA_signal_3781 ;
    wire new_AGEMA_signal_3782 ;
    wire new_AGEMA_signal_3783 ;
    wire new_AGEMA_signal_3784 ;
    wire new_AGEMA_signal_3785 ;
    wire new_AGEMA_signal_3786 ;
    wire new_AGEMA_signal_3787 ;
    wire new_AGEMA_signal_3788 ;
    wire new_AGEMA_signal_3789 ;
    wire new_AGEMA_signal_3790 ;
    wire new_AGEMA_signal_3791 ;
    wire new_AGEMA_signal_3792 ;
    wire new_AGEMA_signal_3793 ;
    wire new_AGEMA_signal_3794 ;
    wire new_AGEMA_signal_3795 ;
    wire new_AGEMA_signal_3796 ;
    wire new_AGEMA_signal_3797 ;
    wire new_AGEMA_signal_3798 ;
    wire new_AGEMA_signal_3799 ;
    wire new_AGEMA_signal_3800 ;
    wire new_AGEMA_signal_3801 ;
    wire new_AGEMA_signal_3802 ;
    wire new_AGEMA_signal_3803 ;
    wire new_AGEMA_signal_3804 ;
    wire new_AGEMA_signal_3805 ;
    wire new_AGEMA_signal_3806 ;
    wire new_AGEMA_signal_3807 ;
    wire new_AGEMA_signal_3808 ;
    wire new_AGEMA_signal_3809 ;
    wire new_AGEMA_signal_3810 ;
    wire new_AGEMA_signal_3811 ;
    wire new_AGEMA_signal_3812 ;
    wire new_AGEMA_signal_3813 ;
    wire new_AGEMA_signal_3814 ;
    wire new_AGEMA_signal_3815 ;
    wire new_AGEMA_signal_3816 ;
    wire new_AGEMA_signal_3817 ;
    wire new_AGEMA_signal_3818 ;
    wire new_AGEMA_signal_3819 ;
    wire new_AGEMA_signal_3820 ;
    wire new_AGEMA_signal_3821 ;
    wire new_AGEMA_signal_3822 ;
    wire new_AGEMA_signal_3823 ;
    wire new_AGEMA_signal_3824 ;
    wire new_AGEMA_signal_3825 ;
    wire new_AGEMA_signal_3826 ;
    wire new_AGEMA_signal_3827 ;
    wire new_AGEMA_signal_3828 ;
    wire new_AGEMA_signal_3829 ;
    wire new_AGEMA_signal_3830 ;
    wire new_AGEMA_signal_3831 ;
    wire new_AGEMA_signal_3832 ;
    wire new_AGEMA_signal_3833 ;
    wire new_AGEMA_signal_3834 ;
    wire new_AGEMA_signal_3835 ;
    wire new_AGEMA_signal_3836 ;
    wire new_AGEMA_signal_3837 ;
    wire new_AGEMA_signal_3838 ;
    wire new_AGEMA_signal_3839 ;
    wire new_AGEMA_signal_3840 ;
    wire new_AGEMA_signal_3841 ;
    wire new_AGEMA_signal_3842 ;
    wire new_AGEMA_signal_3843 ;
    wire new_AGEMA_signal_3844 ;
    wire new_AGEMA_signal_3845 ;
    wire new_AGEMA_signal_3846 ;
    wire new_AGEMA_signal_3847 ;
    wire new_AGEMA_signal_3848 ;
    wire new_AGEMA_signal_3849 ;
    wire new_AGEMA_signal_3850 ;
    wire new_AGEMA_signal_3851 ;
    wire new_AGEMA_signal_3852 ;
    wire new_AGEMA_signal_3853 ;
    wire new_AGEMA_signal_3854 ;
    wire new_AGEMA_signal_3855 ;
    wire new_AGEMA_signal_3856 ;
    wire new_AGEMA_signal_3857 ;
    wire new_AGEMA_signal_3858 ;
    wire new_AGEMA_signal_3859 ;
    wire new_AGEMA_signal_3860 ;
    wire new_AGEMA_signal_3861 ;
    wire new_AGEMA_signal_3862 ;
    wire new_AGEMA_signal_3863 ;
    wire new_AGEMA_signal_3864 ;
    wire new_AGEMA_signal_3865 ;
    wire new_AGEMA_signal_3866 ;
    wire new_AGEMA_signal_3867 ;
    wire new_AGEMA_signal_3868 ;
    wire new_AGEMA_signal_3869 ;
    wire new_AGEMA_signal_3870 ;
    wire new_AGEMA_signal_3871 ;
    wire new_AGEMA_signal_3872 ;
    wire new_AGEMA_signal_3873 ;
    wire new_AGEMA_signal_3874 ;
    wire new_AGEMA_signal_3875 ;
    wire new_AGEMA_signal_3876 ;
    wire new_AGEMA_signal_3877 ;
    wire new_AGEMA_signal_3878 ;
    wire new_AGEMA_signal_3879 ;
    wire new_AGEMA_signal_3880 ;
    wire new_AGEMA_signal_3881 ;
    wire new_AGEMA_signal_3882 ;
    wire new_AGEMA_signal_3883 ;
    wire new_AGEMA_signal_3884 ;
    wire new_AGEMA_signal_3885 ;
    wire new_AGEMA_signal_3886 ;
    wire new_AGEMA_signal_3887 ;
    wire new_AGEMA_signal_3888 ;
    wire new_AGEMA_signal_3889 ;
    wire new_AGEMA_signal_3890 ;
    wire new_AGEMA_signal_3891 ;
    wire new_AGEMA_signal_3892 ;
    wire new_AGEMA_signal_3893 ;
    wire new_AGEMA_signal_3894 ;
    wire new_AGEMA_signal_3895 ;
    wire new_AGEMA_signal_3896 ;
    wire new_AGEMA_signal_3897 ;
    wire new_AGEMA_signal_3898 ;
    wire new_AGEMA_signal_3899 ;
    wire new_AGEMA_signal_3900 ;
    wire new_AGEMA_signal_3901 ;
    wire new_AGEMA_signal_3902 ;
    wire new_AGEMA_signal_3903 ;
    wire new_AGEMA_signal_3904 ;
    wire new_AGEMA_signal_3905 ;
    wire new_AGEMA_signal_3906 ;
    wire new_AGEMA_signal_3907 ;
    wire new_AGEMA_signal_3908 ;
    wire new_AGEMA_signal_3909 ;
    wire new_AGEMA_signal_3910 ;
    wire new_AGEMA_signal_3911 ;
    wire new_AGEMA_signal_3912 ;
    wire new_AGEMA_signal_3913 ;
    wire new_AGEMA_signal_3914 ;
    wire new_AGEMA_signal_3915 ;
    wire new_AGEMA_signal_3916 ;
    wire new_AGEMA_signal_3917 ;
    wire new_AGEMA_signal_3918 ;
    wire new_AGEMA_signal_3919 ;
    wire new_AGEMA_signal_3920 ;
    wire new_AGEMA_signal_3921 ;
    wire new_AGEMA_signal_3922 ;
    wire new_AGEMA_signal_3923 ;
    wire new_AGEMA_signal_3924 ;
    wire new_AGEMA_signal_3925 ;
    wire new_AGEMA_signal_3926 ;
    wire new_AGEMA_signal_3927 ;
    wire new_AGEMA_signal_3928 ;
    wire new_AGEMA_signal_3929 ;
    wire new_AGEMA_signal_3930 ;
    wire new_AGEMA_signal_3931 ;
    wire new_AGEMA_signal_3932 ;
    wire new_AGEMA_signal_3933 ;
    wire new_AGEMA_signal_3934 ;
    wire new_AGEMA_signal_3935 ;
    wire new_AGEMA_signal_3936 ;
    wire new_AGEMA_signal_3937 ;
    wire new_AGEMA_signal_3938 ;
    wire new_AGEMA_signal_3939 ;
    wire new_AGEMA_signal_3940 ;
    wire new_AGEMA_signal_3941 ;
    wire new_AGEMA_signal_3942 ;
    wire new_AGEMA_signal_3943 ;
    wire new_AGEMA_signal_3944 ;
    wire new_AGEMA_signal_3945 ;
    wire new_AGEMA_signal_3946 ;
    wire new_AGEMA_signal_3947 ;
    wire new_AGEMA_signal_3948 ;
    wire new_AGEMA_signal_3949 ;
    wire new_AGEMA_signal_3950 ;
    wire new_AGEMA_signal_3951 ;
    wire new_AGEMA_signal_3952 ;
    wire new_AGEMA_signal_3953 ;
    wire new_AGEMA_signal_3954 ;
    wire new_AGEMA_signal_3955 ;
    wire new_AGEMA_signal_3956 ;
    wire new_AGEMA_signal_3957 ;
    wire new_AGEMA_signal_3958 ;
    wire new_AGEMA_signal_3959 ;
    wire new_AGEMA_signal_3960 ;
    wire new_AGEMA_signal_3961 ;
    wire new_AGEMA_signal_3962 ;
    wire new_AGEMA_signal_3963 ;
    wire new_AGEMA_signal_3964 ;
    wire new_AGEMA_signal_3965 ;
    wire new_AGEMA_signal_3966 ;
    wire new_AGEMA_signal_3967 ;
    wire new_AGEMA_signal_3968 ;
    wire new_AGEMA_signal_3969 ;
    wire new_AGEMA_signal_3970 ;
    wire new_AGEMA_signal_3971 ;
    wire new_AGEMA_signal_3972 ;
    wire new_AGEMA_signal_3973 ;
    wire new_AGEMA_signal_3974 ;
    wire new_AGEMA_signal_3975 ;
    wire new_AGEMA_signal_3976 ;
    wire new_AGEMA_signal_3977 ;
    wire new_AGEMA_signal_3978 ;
    wire new_AGEMA_signal_3979 ;
    wire new_AGEMA_signal_3980 ;
    wire new_AGEMA_signal_3981 ;
    wire new_AGEMA_signal_3982 ;
    wire new_AGEMA_signal_3983 ;
    wire new_AGEMA_signal_3984 ;
    wire new_AGEMA_signal_3985 ;
    wire new_AGEMA_signal_3986 ;
    wire new_AGEMA_signal_3987 ;
    wire new_AGEMA_signal_3988 ;
    wire new_AGEMA_signal_3989 ;
    wire new_AGEMA_signal_3990 ;
    wire new_AGEMA_signal_3991 ;
    wire new_AGEMA_signal_3992 ;
    wire new_AGEMA_signal_3993 ;
    wire new_AGEMA_signal_3994 ;
    wire new_AGEMA_signal_3995 ;
    wire new_AGEMA_signal_3996 ;
    wire new_AGEMA_signal_3997 ;
    wire new_AGEMA_signal_3998 ;
    wire new_AGEMA_signal_3999 ;
    wire new_AGEMA_signal_4000 ;
    wire new_AGEMA_signal_4001 ;
    wire new_AGEMA_signal_4002 ;
    wire new_AGEMA_signal_4003 ;
    wire new_AGEMA_signal_4004 ;
    wire new_AGEMA_signal_4005 ;
    wire new_AGEMA_signal_4006 ;
    wire new_AGEMA_signal_4007 ;
    wire new_AGEMA_signal_4008 ;
    wire new_AGEMA_signal_4009 ;
    wire new_AGEMA_signal_4010 ;
    wire new_AGEMA_signal_4011 ;
    wire new_AGEMA_signal_4012 ;
    wire new_AGEMA_signal_4013 ;
    wire new_AGEMA_signal_4014 ;
    wire new_AGEMA_signal_4015 ;
    wire new_AGEMA_signal_4016 ;
    wire new_AGEMA_signal_4017 ;
    wire new_AGEMA_signal_4018 ;
    wire new_AGEMA_signal_4019 ;
    wire new_AGEMA_signal_4020 ;
    wire new_AGEMA_signal_4021 ;
    wire new_AGEMA_signal_4022 ;
    wire new_AGEMA_signal_4023 ;
    wire new_AGEMA_signal_4024 ;
    wire new_AGEMA_signal_4025 ;
    wire new_AGEMA_signal_4026 ;
    wire new_AGEMA_signal_4027 ;
    wire new_AGEMA_signal_4028 ;
    wire new_AGEMA_signal_4029 ;
    wire new_AGEMA_signal_4030 ;
    wire new_AGEMA_signal_4031 ;
    wire new_AGEMA_signal_4032 ;
    wire new_AGEMA_signal_4033 ;
    wire new_AGEMA_signal_4034 ;
    wire new_AGEMA_signal_4035 ;
    wire new_AGEMA_signal_4036 ;
    wire new_AGEMA_signal_4037 ;
    wire new_AGEMA_signal_4038 ;
    wire new_AGEMA_signal_4039 ;
    wire new_AGEMA_signal_4040 ;
    wire new_AGEMA_signal_4041 ;
    wire new_AGEMA_signal_4042 ;
    wire new_AGEMA_signal_4043 ;
    wire new_AGEMA_signal_4044 ;
    wire new_AGEMA_signal_4045 ;
    wire new_AGEMA_signal_4046 ;
    wire new_AGEMA_signal_4047 ;
    wire new_AGEMA_signal_4048 ;
    wire new_AGEMA_signal_4049 ;
    wire new_AGEMA_signal_4050 ;
    wire new_AGEMA_signal_4051 ;
    wire new_AGEMA_signal_4052 ;
    wire new_AGEMA_signal_4053 ;
    wire new_AGEMA_signal_4054 ;
    wire new_AGEMA_signal_4055 ;
    wire new_AGEMA_signal_4056 ;
    wire new_AGEMA_signal_4057 ;
    wire new_AGEMA_signal_4058 ;
    wire new_AGEMA_signal_4059 ;
    wire new_AGEMA_signal_4060 ;
    wire new_AGEMA_signal_4061 ;
    wire new_AGEMA_signal_4062 ;
    wire new_AGEMA_signal_4063 ;
    wire new_AGEMA_signal_4064 ;
    wire new_AGEMA_signal_4065 ;
    wire new_AGEMA_signal_4066 ;
    wire new_AGEMA_signal_4067 ;
    wire new_AGEMA_signal_4068 ;
    wire new_AGEMA_signal_4069 ;
    wire new_AGEMA_signal_4070 ;
    wire new_AGEMA_signal_4071 ;
    wire new_AGEMA_signal_4072 ;
    wire new_AGEMA_signal_4073 ;
    wire new_AGEMA_signal_4074 ;
    wire new_AGEMA_signal_4075 ;
    wire new_AGEMA_signal_4076 ;
    wire new_AGEMA_signal_4077 ;
    wire new_AGEMA_signal_4078 ;
    wire new_AGEMA_signal_4079 ;
    wire new_AGEMA_signal_4080 ;
    wire new_AGEMA_signal_4081 ;
    wire new_AGEMA_signal_4082 ;
    wire new_AGEMA_signal_4083 ;
    wire new_AGEMA_signal_4084 ;
    wire new_AGEMA_signal_4085 ;
    wire new_AGEMA_signal_4086 ;
    wire new_AGEMA_signal_4087 ;
    wire new_AGEMA_signal_4088 ;
    wire new_AGEMA_signal_4089 ;
    wire new_AGEMA_signal_4090 ;
    wire new_AGEMA_signal_4091 ;
    wire new_AGEMA_signal_4092 ;
    wire new_AGEMA_signal_4093 ;
    wire new_AGEMA_signal_4094 ;
    wire new_AGEMA_signal_4095 ;
    wire new_AGEMA_signal_4096 ;
    wire new_AGEMA_signal_4097 ;
    wire new_AGEMA_signal_4098 ;
    wire new_AGEMA_signal_4099 ;
    wire new_AGEMA_signal_4100 ;
    wire new_AGEMA_signal_4101 ;
    wire new_AGEMA_signal_4102 ;
    wire new_AGEMA_signal_4103 ;
    wire new_AGEMA_signal_4104 ;
    wire new_AGEMA_signal_4105 ;
    wire new_AGEMA_signal_4106 ;
    wire new_AGEMA_signal_4107 ;
    wire new_AGEMA_signal_4108 ;
    wire new_AGEMA_signal_4109 ;
    wire new_AGEMA_signal_4110 ;
    wire new_AGEMA_signal_4111 ;
    wire new_AGEMA_signal_4112 ;
    wire new_AGEMA_signal_4113 ;
    wire new_AGEMA_signal_4114 ;
    wire new_AGEMA_signal_4115 ;
    wire new_AGEMA_signal_4116 ;
    wire new_AGEMA_signal_4117 ;
    wire new_AGEMA_signal_4118 ;
    wire new_AGEMA_signal_4119 ;
    wire new_AGEMA_signal_4120 ;
    wire new_AGEMA_signal_4121 ;
    wire new_AGEMA_signal_4122 ;
    wire new_AGEMA_signal_4123 ;
    wire new_AGEMA_signal_4124 ;
    wire new_AGEMA_signal_4125 ;
    wire new_AGEMA_signal_4126 ;
    wire new_AGEMA_signal_4127 ;
    wire new_AGEMA_signal_4128 ;
    wire new_AGEMA_signal_4129 ;
    wire new_AGEMA_signal_4130 ;
    wire new_AGEMA_signal_4131 ;
    wire new_AGEMA_signal_4132 ;
    wire new_AGEMA_signal_4133 ;
    wire new_AGEMA_signal_4134 ;
    wire new_AGEMA_signal_4135 ;
    wire new_AGEMA_signal_4136 ;
    wire new_AGEMA_signal_4137 ;
    wire new_AGEMA_signal_4138 ;
    wire new_AGEMA_signal_4139 ;
    wire new_AGEMA_signal_4140 ;
    wire new_AGEMA_signal_4141 ;
    wire new_AGEMA_signal_4142 ;
    wire new_AGEMA_signal_4143 ;
    wire new_AGEMA_signal_4144 ;
    wire new_AGEMA_signal_4145 ;
    wire new_AGEMA_signal_4146 ;
    wire new_AGEMA_signal_4147 ;
    wire new_AGEMA_signal_4148 ;
    wire new_AGEMA_signal_4149 ;
    wire new_AGEMA_signal_4150 ;
    wire new_AGEMA_signal_4151 ;
    wire new_AGEMA_signal_4152 ;
    wire new_AGEMA_signal_4153 ;
    wire new_AGEMA_signal_4154 ;
    wire new_AGEMA_signal_4155 ;
    wire new_AGEMA_signal_4156 ;
    wire new_AGEMA_signal_4157 ;
    wire new_AGEMA_signal_4158 ;
    wire new_AGEMA_signal_4159 ;
    wire new_AGEMA_signal_4160 ;
    wire new_AGEMA_signal_4161 ;
    wire new_AGEMA_signal_4162 ;
    wire new_AGEMA_signal_4163 ;
    wire new_AGEMA_signal_4164 ;
    wire new_AGEMA_signal_4165 ;
    wire new_AGEMA_signal_4166 ;
    wire new_AGEMA_signal_4167 ;
    wire new_AGEMA_signal_4168 ;
    wire new_AGEMA_signal_4169 ;
    wire new_AGEMA_signal_4170 ;
    wire new_AGEMA_signal_4171 ;
    wire new_AGEMA_signal_4172 ;
    wire new_AGEMA_signal_4173 ;
    wire new_AGEMA_signal_4174 ;
    wire new_AGEMA_signal_4175 ;
    wire new_AGEMA_signal_4176 ;
    wire new_AGEMA_signal_4177 ;
    wire new_AGEMA_signal_4178 ;
    wire new_AGEMA_signal_4179 ;
    wire new_AGEMA_signal_4180 ;
    wire new_AGEMA_signal_4181 ;
    wire new_AGEMA_signal_4182 ;
    wire new_AGEMA_signal_4183 ;
    wire new_AGEMA_signal_4184 ;
    wire new_AGEMA_signal_4185 ;
    wire new_AGEMA_signal_4186 ;
    wire new_AGEMA_signal_4187 ;
    wire new_AGEMA_signal_4188 ;
    wire new_AGEMA_signal_4189 ;
    wire new_AGEMA_signal_4190 ;
    wire new_AGEMA_signal_4191 ;
    wire new_AGEMA_signal_4192 ;
    wire new_AGEMA_signal_4193 ;
    wire new_AGEMA_signal_4194 ;
    wire new_AGEMA_signal_4195 ;
    wire new_AGEMA_signal_4196 ;
    wire new_AGEMA_signal_4197 ;
    wire new_AGEMA_signal_4198 ;
    wire new_AGEMA_signal_4199 ;
    wire new_AGEMA_signal_4200 ;
    wire new_AGEMA_signal_4201 ;
    wire new_AGEMA_signal_4202 ;
    wire new_AGEMA_signal_4203 ;
    wire new_AGEMA_signal_4204 ;
    wire new_AGEMA_signal_4205 ;
    wire new_AGEMA_signal_4206 ;
    wire new_AGEMA_signal_4207 ;
    wire new_AGEMA_signal_4208 ;
    wire new_AGEMA_signal_4209 ;
    wire new_AGEMA_signal_4210 ;
    wire new_AGEMA_signal_4211 ;
    wire new_AGEMA_signal_4212 ;
    wire new_AGEMA_signal_4213 ;
    wire new_AGEMA_signal_4214 ;
    wire new_AGEMA_signal_4215 ;
    wire new_AGEMA_signal_4216 ;
    wire new_AGEMA_signal_4217 ;
    wire new_AGEMA_signal_4218 ;
    wire new_AGEMA_signal_4219 ;
    wire new_AGEMA_signal_4220 ;
    wire new_AGEMA_signal_4221 ;
    wire new_AGEMA_signal_4222 ;
    wire new_AGEMA_signal_4223 ;
    wire new_AGEMA_signal_4224 ;
    wire new_AGEMA_signal_4225 ;
    wire new_AGEMA_signal_4226 ;
    wire new_AGEMA_signal_4227 ;
    wire new_AGEMA_signal_4228 ;
    wire new_AGEMA_signal_4229 ;
    wire new_AGEMA_signal_4230 ;
    wire new_AGEMA_signal_4231 ;
    wire new_AGEMA_signal_4232 ;
    wire new_AGEMA_signal_4233 ;
    wire new_AGEMA_signal_4234 ;
    wire new_AGEMA_signal_4235 ;
    wire new_AGEMA_signal_4236 ;
    wire new_AGEMA_signal_4237 ;
    wire new_AGEMA_signal_4238 ;
    wire new_AGEMA_signal_4239 ;
    wire new_AGEMA_signal_4240 ;
    wire new_AGEMA_signal_4241 ;
    wire new_AGEMA_signal_4242 ;
    wire new_AGEMA_signal_4243 ;
    wire new_AGEMA_signal_4244 ;
    wire new_AGEMA_signal_4245 ;
    wire new_AGEMA_signal_4246 ;
    wire new_AGEMA_signal_4247 ;
    wire new_AGEMA_signal_4248 ;
    wire new_AGEMA_signal_4249 ;
    wire new_AGEMA_signal_4250 ;
    wire new_AGEMA_signal_4251 ;
    wire new_AGEMA_signal_4252 ;
    wire new_AGEMA_signal_4253 ;
    wire new_AGEMA_signal_4254 ;
    wire new_AGEMA_signal_4255 ;
    wire new_AGEMA_signal_4256 ;
    wire new_AGEMA_signal_4257 ;
    wire new_AGEMA_signal_4258 ;
    wire new_AGEMA_signal_4259 ;
    wire new_AGEMA_signal_4260 ;
    wire new_AGEMA_signal_4261 ;
    wire new_AGEMA_signal_4262 ;
    wire new_AGEMA_signal_4263 ;
    wire new_AGEMA_signal_4264 ;
    wire new_AGEMA_signal_4265 ;
    wire new_AGEMA_signal_4266 ;
    wire new_AGEMA_signal_4267 ;
    wire new_AGEMA_signal_4268 ;
    wire new_AGEMA_signal_4269 ;
    wire new_AGEMA_signal_4270 ;
    wire new_AGEMA_signal_4271 ;
    wire new_AGEMA_signal_4272 ;
    wire new_AGEMA_signal_4273 ;
    wire new_AGEMA_signal_4274 ;
    wire new_AGEMA_signal_4275 ;
    wire new_AGEMA_signal_4276 ;
    wire new_AGEMA_signal_4277 ;
    wire new_AGEMA_signal_4278 ;
    wire new_AGEMA_signal_4279 ;
    wire new_AGEMA_signal_4280 ;
    wire new_AGEMA_signal_4281 ;
    wire new_AGEMA_signal_4282 ;
    wire new_AGEMA_signal_4283 ;
    wire new_AGEMA_signal_4284 ;
    wire new_AGEMA_signal_4285 ;
    wire new_AGEMA_signal_4286 ;
    wire new_AGEMA_signal_4287 ;
    wire new_AGEMA_signal_4288 ;
    wire new_AGEMA_signal_4289 ;
    wire new_AGEMA_signal_4290 ;
    wire new_AGEMA_signal_4291 ;
    wire new_AGEMA_signal_4292 ;
    wire new_AGEMA_signal_4293 ;
    wire new_AGEMA_signal_4294 ;
    wire new_AGEMA_signal_4295 ;
    wire new_AGEMA_signal_4296 ;
    wire new_AGEMA_signal_4297 ;
    wire new_AGEMA_signal_4298 ;
    wire new_AGEMA_signal_4299 ;
    wire new_AGEMA_signal_4300 ;
    wire new_AGEMA_signal_4301 ;
    wire new_AGEMA_signal_4302 ;
    wire new_AGEMA_signal_4303 ;
    wire new_AGEMA_signal_4304 ;
    wire new_AGEMA_signal_4305 ;
    wire new_AGEMA_signal_4306 ;
    wire new_AGEMA_signal_4307 ;
    wire new_AGEMA_signal_4308 ;
    wire new_AGEMA_signal_4309 ;
    wire new_AGEMA_signal_4310 ;
    wire new_AGEMA_signal_4311 ;
    wire new_AGEMA_signal_4312 ;
    wire new_AGEMA_signal_4313 ;
    wire new_AGEMA_signal_4314 ;
    wire new_AGEMA_signal_4315 ;
    wire new_AGEMA_signal_4316 ;
    wire new_AGEMA_signal_4317 ;
    wire new_AGEMA_signal_4318 ;
    wire new_AGEMA_signal_4319 ;
    wire new_AGEMA_signal_4320 ;
    wire new_AGEMA_signal_4321 ;
    wire new_AGEMA_signal_4322 ;
    wire new_AGEMA_signal_4323 ;
    wire new_AGEMA_signal_4324 ;
    wire new_AGEMA_signal_4325 ;
    wire new_AGEMA_signal_4326 ;
    wire new_AGEMA_signal_4327 ;
    wire new_AGEMA_signal_4328 ;
    wire new_AGEMA_signal_4329 ;
    wire new_AGEMA_signal_4330 ;
    wire new_AGEMA_signal_4331 ;
    wire new_AGEMA_signal_4332 ;
    wire new_AGEMA_signal_4333 ;
    wire new_AGEMA_signal_4334 ;
    wire new_AGEMA_signal_4335 ;
    wire new_AGEMA_signal_4336 ;
    wire new_AGEMA_signal_4337 ;
    wire new_AGEMA_signal_4338 ;
    wire new_AGEMA_signal_4339 ;
    wire new_AGEMA_signal_4340 ;
    wire new_AGEMA_signal_4341 ;
    wire new_AGEMA_signal_4342 ;
    wire new_AGEMA_signal_4343 ;
    wire new_AGEMA_signal_4344 ;
    wire new_AGEMA_signal_4345 ;
    wire new_AGEMA_signal_4346 ;
    wire new_AGEMA_signal_4347 ;
    wire new_AGEMA_signal_4348 ;
    wire new_AGEMA_signal_4349 ;
    wire new_AGEMA_signal_4350 ;
    wire new_AGEMA_signal_4351 ;
    wire new_AGEMA_signal_4352 ;
    wire new_AGEMA_signal_4353 ;
    wire new_AGEMA_signal_4354 ;
    wire new_AGEMA_signal_4355 ;
    wire new_AGEMA_signal_4356 ;
    wire new_AGEMA_signal_4357 ;
    wire new_AGEMA_signal_4358 ;
    wire new_AGEMA_signal_4359 ;
    wire new_AGEMA_signal_4360 ;
    wire new_AGEMA_signal_4361 ;
    wire new_AGEMA_signal_4362 ;
    wire new_AGEMA_signal_4363 ;
    wire new_AGEMA_signal_4364 ;
    wire new_AGEMA_signal_4365 ;
    wire new_AGEMA_signal_4366 ;
    wire new_AGEMA_signal_4367 ;
    wire new_AGEMA_signal_4368 ;
    wire new_AGEMA_signal_4369 ;
    wire new_AGEMA_signal_4370 ;
    wire new_AGEMA_signal_4371 ;
    wire new_AGEMA_signal_4372 ;
    wire new_AGEMA_signal_4373 ;
    wire new_AGEMA_signal_4374 ;
    wire new_AGEMA_signal_4375 ;
    wire new_AGEMA_signal_4376 ;
    wire new_AGEMA_signal_4377 ;
    wire new_AGEMA_signal_4378 ;
    wire new_AGEMA_signal_4379 ;
    wire new_AGEMA_signal_4380 ;
    wire new_AGEMA_signal_4381 ;
    wire new_AGEMA_signal_4382 ;
    wire new_AGEMA_signal_4383 ;
    wire new_AGEMA_signal_4384 ;
    wire new_AGEMA_signal_4385 ;
    wire new_AGEMA_signal_4386 ;
    wire new_AGEMA_signal_4387 ;
    wire new_AGEMA_signal_4388 ;
    wire new_AGEMA_signal_4389 ;
    wire new_AGEMA_signal_4390 ;
    wire new_AGEMA_signal_4391 ;
    wire new_AGEMA_signal_4392 ;
    wire new_AGEMA_signal_4393 ;
    wire new_AGEMA_signal_4394 ;
    wire new_AGEMA_signal_4395 ;
    wire new_AGEMA_signal_4396 ;
    wire new_AGEMA_signal_4397 ;
    wire new_AGEMA_signal_4398 ;
    wire new_AGEMA_signal_4399 ;
    wire new_AGEMA_signal_4400 ;
    wire new_AGEMA_signal_4401 ;
    wire new_AGEMA_signal_4402 ;
    wire new_AGEMA_signal_4403 ;
    wire new_AGEMA_signal_4404 ;
    wire new_AGEMA_signal_4405 ;
    wire new_AGEMA_signal_4406 ;
    wire new_AGEMA_signal_4407 ;
    wire new_AGEMA_signal_4408 ;
    wire new_AGEMA_signal_4409 ;
    wire new_AGEMA_signal_4410 ;
    wire new_AGEMA_signal_4411 ;
    wire new_AGEMA_signal_4412 ;
    wire new_AGEMA_signal_4413 ;
    wire new_AGEMA_signal_4414 ;
    wire new_AGEMA_signal_4415 ;
    wire new_AGEMA_signal_4416 ;
    wire new_AGEMA_signal_4417 ;
    wire new_AGEMA_signal_4418 ;
    wire new_AGEMA_signal_4419 ;
    wire new_AGEMA_signal_4420 ;
    wire new_AGEMA_signal_4421 ;
    wire new_AGEMA_signal_4422 ;
    wire new_AGEMA_signal_4423 ;
    wire new_AGEMA_signal_4424 ;
    wire new_AGEMA_signal_4425 ;
    wire new_AGEMA_signal_4426 ;
    wire new_AGEMA_signal_4427 ;
    wire new_AGEMA_signal_4428 ;
    wire new_AGEMA_signal_4429 ;
    wire new_AGEMA_signal_4430 ;
    wire new_AGEMA_signal_4431 ;
    wire new_AGEMA_signal_4432 ;
    wire new_AGEMA_signal_4433 ;
    wire new_AGEMA_signal_4434 ;
    wire new_AGEMA_signal_4435 ;
    wire new_AGEMA_signal_4436 ;
    wire new_AGEMA_signal_4437 ;
    wire new_AGEMA_signal_4438 ;
    wire new_AGEMA_signal_4439 ;
    wire new_AGEMA_signal_4440 ;
    wire new_AGEMA_signal_4441 ;
    wire new_AGEMA_signal_4442 ;
    wire new_AGEMA_signal_4443 ;
    wire new_AGEMA_signal_4444 ;
    wire new_AGEMA_signal_4445 ;
    wire new_AGEMA_signal_4446 ;
    wire new_AGEMA_signal_4447 ;
    wire new_AGEMA_signal_4448 ;
    wire new_AGEMA_signal_4449 ;
    wire new_AGEMA_signal_4450 ;
    wire new_AGEMA_signal_4451 ;
    wire new_AGEMA_signal_4452 ;
    wire new_AGEMA_signal_4453 ;
    wire new_AGEMA_signal_4454 ;
    wire new_AGEMA_signal_4455 ;
    wire new_AGEMA_signal_4456 ;
    wire new_AGEMA_signal_4457 ;
    wire new_AGEMA_signal_4458 ;
    wire new_AGEMA_signal_4459 ;
    wire new_AGEMA_signal_4460 ;
    wire new_AGEMA_signal_4461 ;
    wire new_AGEMA_signal_4462 ;
    wire new_AGEMA_signal_4463 ;
    wire new_AGEMA_signal_4464 ;
    wire new_AGEMA_signal_4465 ;
    wire new_AGEMA_signal_4466 ;
    wire new_AGEMA_signal_4467 ;
    wire new_AGEMA_signal_4468 ;
    wire new_AGEMA_signal_4469 ;
    wire new_AGEMA_signal_4470 ;
    wire new_AGEMA_signal_4471 ;
    wire new_AGEMA_signal_4472 ;
    wire new_AGEMA_signal_4473 ;
    wire new_AGEMA_signal_4474 ;
    wire new_AGEMA_signal_4475 ;
    wire new_AGEMA_signal_4476 ;
    wire new_AGEMA_signal_4477 ;
    wire new_AGEMA_signal_4478 ;
    wire new_AGEMA_signal_4479 ;
    wire new_AGEMA_signal_4480 ;
    wire new_AGEMA_signal_4481 ;
    wire new_AGEMA_signal_4482 ;
    wire new_AGEMA_signal_4483 ;
    wire new_AGEMA_signal_4484 ;
    wire new_AGEMA_signal_4485 ;
    wire new_AGEMA_signal_4486 ;
    wire new_AGEMA_signal_4487 ;
    wire new_AGEMA_signal_4488 ;
    wire new_AGEMA_signal_4489 ;
    wire new_AGEMA_signal_4490 ;
    wire new_AGEMA_signal_4491 ;
    wire new_AGEMA_signal_4492 ;
    wire new_AGEMA_signal_4493 ;
    wire new_AGEMA_signal_4494 ;
    wire new_AGEMA_signal_4495 ;
    wire new_AGEMA_signal_4496 ;
    wire new_AGEMA_signal_4497 ;
    wire new_AGEMA_signal_4498 ;
    wire new_AGEMA_signal_4499 ;
    wire new_AGEMA_signal_4500 ;
    wire new_AGEMA_signal_4501 ;
    wire new_AGEMA_signal_4502 ;
    wire new_AGEMA_signal_4503 ;
    wire new_AGEMA_signal_4504 ;
    wire new_AGEMA_signal_4505 ;
    wire new_AGEMA_signal_4506 ;
    wire new_AGEMA_signal_4507 ;
    wire new_AGEMA_signal_4508 ;
    wire new_AGEMA_signal_4509 ;
    wire new_AGEMA_signal_4510 ;
    wire new_AGEMA_signal_4511 ;
    wire new_AGEMA_signal_4512 ;
    wire new_AGEMA_signal_4513 ;
    wire new_AGEMA_signal_4514 ;
    wire new_AGEMA_signal_4515 ;
    wire new_AGEMA_signal_4516 ;
    wire new_AGEMA_signal_4517 ;
    wire new_AGEMA_signal_4518 ;
    wire new_AGEMA_signal_4519 ;
    wire new_AGEMA_signal_4520 ;
    wire new_AGEMA_signal_4521 ;
    wire new_AGEMA_signal_4522 ;
    wire new_AGEMA_signal_4523 ;
    wire new_AGEMA_signal_4524 ;
    wire new_AGEMA_signal_4525 ;
    wire new_AGEMA_signal_4526 ;
    wire new_AGEMA_signal_4527 ;
    wire new_AGEMA_signal_4528 ;
    wire new_AGEMA_signal_4529 ;
    wire new_AGEMA_signal_4530 ;
    wire new_AGEMA_signal_4531 ;
    wire new_AGEMA_signal_4532 ;
    wire new_AGEMA_signal_4533 ;
    wire new_AGEMA_signal_4534 ;
    wire new_AGEMA_signal_4535 ;
    wire new_AGEMA_signal_4536 ;
    wire new_AGEMA_signal_4537 ;
    wire new_AGEMA_signal_4538 ;
    wire new_AGEMA_signal_4539 ;
    wire new_AGEMA_signal_4540 ;
    wire new_AGEMA_signal_4541 ;
    wire new_AGEMA_signal_4542 ;
    wire new_AGEMA_signal_4543 ;
    wire new_AGEMA_signal_4544 ;
    wire new_AGEMA_signal_4545 ;
    wire new_AGEMA_signal_4546 ;
    wire new_AGEMA_signal_4547 ;
    wire new_AGEMA_signal_4548 ;
    wire new_AGEMA_signal_4549 ;
    wire new_AGEMA_signal_4550 ;
    wire new_AGEMA_signal_4551 ;
    wire new_AGEMA_signal_4552 ;
    wire new_AGEMA_signal_4553 ;
    wire new_AGEMA_signal_4554 ;
    wire new_AGEMA_signal_4555 ;
    wire new_AGEMA_signal_4556 ;
    wire new_AGEMA_signal_4557 ;
    wire new_AGEMA_signal_4558 ;
    wire new_AGEMA_signal_4559 ;
    wire new_AGEMA_signal_4560 ;
    wire new_AGEMA_signal_4561 ;
    wire new_AGEMA_signal_4562 ;
    wire new_AGEMA_signal_4563 ;
    wire new_AGEMA_signal_4564 ;
    wire new_AGEMA_signal_4565 ;
    wire new_AGEMA_signal_4566 ;
    wire new_AGEMA_signal_4567 ;
    wire new_AGEMA_signal_4568 ;
    wire new_AGEMA_signal_4569 ;
    wire new_AGEMA_signal_4570 ;
    wire new_AGEMA_signal_4571 ;
    wire new_AGEMA_signal_4572 ;
    wire new_AGEMA_signal_4573 ;
    wire new_AGEMA_signal_4574 ;
    wire new_AGEMA_signal_4575 ;
    wire new_AGEMA_signal_4576 ;
    wire new_AGEMA_signal_4577 ;
    wire new_AGEMA_signal_4578 ;
    wire new_AGEMA_signal_4579 ;
    wire new_AGEMA_signal_4580 ;
    wire new_AGEMA_signal_4581 ;
    wire new_AGEMA_signal_4582 ;
    wire new_AGEMA_signal_4583 ;
    wire new_AGEMA_signal_4584 ;
    wire new_AGEMA_signal_4585 ;
    wire new_AGEMA_signal_4586 ;
    wire new_AGEMA_signal_4587 ;
    wire new_AGEMA_signal_4588 ;
    wire new_AGEMA_signal_4589 ;
    wire new_AGEMA_signal_4590 ;
    wire new_AGEMA_signal_4591 ;
    wire new_AGEMA_signal_4592 ;
    wire new_AGEMA_signal_4593 ;
    wire new_AGEMA_signal_4594 ;
    wire new_AGEMA_signal_4595 ;
    wire new_AGEMA_signal_4596 ;
    wire new_AGEMA_signal_4597 ;
    wire new_AGEMA_signal_4598 ;
    wire new_AGEMA_signal_4599 ;
    wire new_AGEMA_signal_4600 ;
    wire new_AGEMA_signal_4601 ;
    wire new_AGEMA_signal_4602 ;
    wire new_AGEMA_signal_4603 ;
    wire new_AGEMA_signal_4604 ;
    wire new_AGEMA_signal_4605 ;
    wire new_AGEMA_signal_4606 ;
    wire new_AGEMA_signal_4607 ;
    wire new_AGEMA_signal_4608 ;
    wire new_AGEMA_signal_4609 ;
    wire new_AGEMA_signal_4610 ;
    wire new_AGEMA_signal_4611 ;
    wire new_AGEMA_signal_4612 ;
    wire new_AGEMA_signal_4613 ;
    wire new_AGEMA_signal_4614 ;
    wire new_AGEMA_signal_4615 ;
    wire new_AGEMA_signal_4616 ;
    wire new_AGEMA_signal_4617 ;
    wire new_AGEMA_signal_4618 ;
    wire new_AGEMA_signal_4619 ;
    wire new_AGEMA_signal_4620 ;
    wire new_AGEMA_signal_4621 ;
    wire new_AGEMA_signal_4622 ;
    wire new_AGEMA_signal_4623 ;
    wire new_AGEMA_signal_4624 ;
    wire new_AGEMA_signal_4625 ;
    wire new_AGEMA_signal_4626 ;
    wire new_AGEMA_signal_4627 ;
    wire new_AGEMA_signal_4628 ;
    wire new_AGEMA_signal_4629 ;
    wire new_AGEMA_signal_4630 ;
    wire new_AGEMA_signal_4631 ;
    wire new_AGEMA_signal_4632 ;
    wire new_AGEMA_signal_4633 ;
    wire new_AGEMA_signal_4634 ;
    wire new_AGEMA_signal_4635 ;
    wire new_AGEMA_signal_4636 ;
    wire new_AGEMA_signal_4637 ;
    wire new_AGEMA_signal_4638 ;
    wire new_AGEMA_signal_4639 ;
    wire new_AGEMA_signal_4640 ;
    wire new_AGEMA_signal_4641 ;
    wire new_AGEMA_signal_4642 ;
    wire new_AGEMA_signal_4643 ;
    wire new_AGEMA_signal_4644 ;
    wire new_AGEMA_signal_4645 ;
    wire new_AGEMA_signal_4646 ;
    wire new_AGEMA_signal_4647 ;
    wire new_AGEMA_signal_4648 ;
    wire new_AGEMA_signal_4649 ;
    wire new_AGEMA_signal_4650 ;
    wire new_AGEMA_signal_4651 ;
    wire new_AGEMA_signal_4652 ;
    wire new_AGEMA_signal_4653 ;
    wire new_AGEMA_signal_4654 ;
    wire new_AGEMA_signal_4655 ;
    wire new_AGEMA_signal_4656 ;
    wire new_AGEMA_signal_4657 ;
    wire new_AGEMA_signal_4658 ;
    wire new_AGEMA_signal_4659 ;
    wire new_AGEMA_signal_4660 ;
    wire new_AGEMA_signal_4661 ;
    wire new_AGEMA_signal_4662 ;
    wire new_AGEMA_signal_4663 ;
    wire new_AGEMA_signal_4664 ;
    wire new_AGEMA_signal_4665 ;
    wire new_AGEMA_signal_4666 ;
    wire new_AGEMA_signal_4667 ;
    wire new_AGEMA_signal_4668 ;
    wire new_AGEMA_signal_4669 ;
    wire new_AGEMA_signal_4670 ;
    wire new_AGEMA_signal_4671 ;
    wire new_AGEMA_signal_4672 ;
    wire new_AGEMA_signal_4673 ;
    wire new_AGEMA_signal_4674 ;
    wire new_AGEMA_signal_4675 ;
    wire new_AGEMA_signal_4676 ;
    wire new_AGEMA_signal_4677 ;
    wire new_AGEMA_signal_4678 ;
    wire new_AGEMA_signal_4679 ;
    wire new_AGEMA_signal_4680 ;
    wire new_AGEMA_signal_4681 ;
    wire new_AGEMA_signal_4682 ;
    wire new_AGEMA_signal_4683 ;
    wire new_AGEMA_signal_4684 ;
    wire new_AGEMA_signal_4685 ;
    wire new_AGEMA_signal_4686 ;
    wire new_AGEMA_signal_4687 ;
    wire new_AGEMA_signal_4688 ;
    wire new_AGEMA_signal_4689 ;
    wire new_AGEMA_signal_4690 ;
    wire new_AGEMA_signal_4691 ;
    wire new_AGEMA_signal_4692 ;
    wire new_AGEMA_signal_4693 ;
    wire new_AGEMA_signal_4694 ;
    wire new_AGEMA_signal_4695 ;
    wire new_AGEMA_signal_4696 ;
    wire new_AGEMA_signal_4697 ;
    wire new_AGEMA_signal_4698 ;
    wire new_AGEMA_signal_4699 ;
    wire new_AGEMA_signal_4700 ;
    wire new_AGEMA_signal_4701 ;
    wire new_AGEMA_signal_4702 ;
    wire new_AGEMA_signal_4703 ;
    wire new_AGEMA_signal_4704 ;
    wire new_AGEMA_signal_4705 ;
    wire new_AGEMA_signal_4706 ;
    wire new_AGEMA_signal_4707 ;
    wire new_AGEMA_signal_4708 ;
    wire new_AGEMA_signal_4709 ;
    wire new_AGEMA_signal_4710 ;
    wire new_AGEMA_signal_4711 ;
    wire new_AGEMA_signal_4712 ;
    wire new_AGEMA_signal_4713 ;
    wire new_AGEMA_signal_4714 ;
    wire new_AGEMA_signal_4715 ;
    wire new_AGEMA_signal_4716 ;
    wire new_AGEMA_signal_4717 ;
    wire new_AGEMA_signal_4718 ;
    wire new_AGEMA_signal_4719 ;
    wire new_AGEMA_signal_4720 ;
    wire new_AGEMA_signal_4721 ;
    wire new_AGEMA_signal_4722 ;
    wire new_AGEMA_signal_4723 ;
    wire new_AGEMA_signal_4724 ;
    wire new_AGEMA_signal_4725 ;
    wire new_AGEMA_signal_4726 ;
    wire new_AGEMA_signal_4727 ;
    wire new_AGEMA_signal_4728 ;
    wire new_AGEMA_signal_4729 ;
    wire new_AGEMA_signal_4730 ;
    wire new_AGEMA_signal_4731 ;
    wire new_AGEMA_signal_4732 ;
    wire new_AGEMA_signal_4733 ;
    wire new_AGEMA_signal_4734 ;
    wire new_AGEMA_signal_4735 ;
    wire new_AGEMA_signal_4736 ;
    wire new_AGEMA_signal_4737 ;
    wire new_AGEMA_signal_4738 ;
    wire new_AGEMA_signal_4739 ;
    wire new_AGEMA_signal_4740 ;
    wire new_AGEMA_signal_4741 ;
    wire new_AGEMA_signal_4742 ;
    wire new_AGEMA_signal_4743 ;
    wire new_AGEMA_signal_4744 ;
    wire new_AGEMA_signal_4745 ;
    wire new_AGEMA_signal_4746 ;
    wire new_AGEMA_signal_4747 ;
    wire new_AGEMA_signal_4748 ;
    wire new_AGEMA_signal_4749 ;
    wire new_AGEMA_signal_4750 ;
    wire new_AGEMA_signal_4751 ;
    wire new_AGEMA_signal_4752 ;
    wire new_AGEMA_signal_4753 ;
    wire new_AGEMA_signal_4754 ;
    wire new_AGEMA_signal_4755 ;
    wire new_AGEMA_signal_4756 ;
    wire new_AGEMA_signal_4757 ;
    wire new_AGEMA_signal_4758 ;
    wire new_AGEMA_signal_4759 ;
    wire new_AGEMA_signal_4760 ;
    wire new_AGEMA_signal_4761 ;
    wire new_AGEMA_signal_4762 ;
    wire new_AGEMA_signal_4763 ;
    wire new_AGEMA_signal_4764 ;
    wire new_AGEMA_signal_4765 ;
    wire new_AGEMA_signal_4766 ;
    wire new_AGEMA_signal_4767 ;
    wire new_AGEMA_signal_4768 ;
    wire new_AGEMA_signal_4769 ;
    wire new_AGEMA_signal_4770 ;
    wire new_AGEMA_signal_4771 ;
    wire new_AGEMA_signal_4772 ;
    wire new_AGEMA_signal_4773 ;
    wire new_AGEMA_signal_4774 ;
    wire new_AGEMA_signal_4775 ;
    wire new_AGEMA_signal_4776 ;
    wire new_AGEMA_signal_4777 ;
    wire new_AGEMA_signal_4778 ;
    wire new_AGEMA_signal_4779 ;
    wire new_AGEMA_signal_4780 ;
    wire new_AGEMA_signal_4781 ;
    wire new_AGEMA_signal_4782 ;
    wire new_AGEMA_signal_4783 ;
    wire new_AGEMA_signal_4784 ;
    wire new_AGEMA_signal_4785 ;
    wire new_AGEMA_signal_4786 ;
    wire new_AGEMA_signal_4787 ;
    wire new_AGEMA_signal_4788 ;
    wire new_AGEMA_signal_4789 ;
    wire new_AGEMA_signal_4790 ;
    wire new_AGEMA_signal_4791 ;
    wire new_AGEMA_signal_4792 ;
    wire new_AGEMA_signal_4793 ;
    wire new_AGEMA_signal_4794 ;
    wire new_AGEMA_signal_4795 ;
    wire new_AGEMA_signal_4796 ;
    wire new_AGEMA_signal_4797 ;
    wire new_AGEMA_signal_4798 ;
    wire new_AGEMA_signal_4799 ;
    wire new_AGEMA_signal_4800 ;
    wire new_AGEMA_signal_4801 ;
    wire new_AGEMA_signal_4802 ;
    wire new_AGEMA_signal_4803 ;
    wire new_AGEMA_signal_4804 ;
    wire new_AGEMA_signal_4805 ;
    wire new_AGEMA_signal_4806 ;
    wire new_AGEMA_signal_4807 ;
    wire new_AGEMA_signal_4808 ;
    wire new_AGEMA_signal_4809 ;
    wire new_AGEMA_signal_4810 ;
    wire new_AGEMA_signal_4811 ;
    wire new_AGEMA_signal_4812 ;
    wire new_AGEMA_signal_4813 ;
    wire new_AGEMA_signal_4814 ;
    wire new_AGEMA_signal_4815 ;
    wire new_AGEMA_signal_4816 ;
    wire new_AGEMA_signal_4817 ;
    wire new_AGEMA_signal_4818 ;
    wire new_AGEMA_signal_4819 ;
    wire new_AGEMA_signal_4820 ;
    wire new_AGEMA_signal_4821 ;
    wire new_AGEMA_signal_4822 ;
    wire new_AGEMA_signal_4823 ;
    wire new_AGEMA_signal_4824 ;
    wire new_AGEMA_signal_4825 ;
    wire new_AGEMA_signal_4826 ;
    wire new_AGEMA_signal_4827 ;
    wire new_AGEMA_signal_4828 ;
    wire new_AGEMA_signal_4829 ;
    wire new_AGEMA_signal_4830 ;
    wire new_AGEMA_signal_4831 ;
    wire new_AGEMA_signal_4832 ;
    wire new_AGEMA_signal_4833 ;
    wire new_AGEMA_signal_4834 ;
    wire new_AGEMA_signal_4835 ;
    wire new_AGEMA_signal_4836 ;
    wire new_AGEMA_signal_4837 ;
    wire new_AGEMA_signal_4838 ;
    wire new_AGEMA_signal_4839 ;
    wire new_AGEMA_signal_4840 ;
    wire new_AGEMA_signal_4841 ;
    wire new_AGEMA_signal_4842 ;
    wire new_AGEMA_signal_4843 ;
    wire new_AGEMA_signal_4844 ;
    wire new_AGEMA_signal_4845 ;
    wire new_AGEMA_signal_4846 ;
    wire new_AGEMA_signal_4847 ;
    wire new_AGEMA_signal_4848 ;
    wire new_AGEMA_signal_4849 ;
    wire new_AGEMA_signal_4850 ;
    wire new_AGEMA_signal_4851 ;
    wire new_AGEMA_signal_4852 ;
    wire new_AGEMA_signal_4853 ;
    wire new_AGEMA_signal_4854 ;
    wire new_AGEMA_signal_4855 ;
    wire new_AGEMA_signal_4856 ;
    wire new_AGEMA_signal_4857 ;
    wire new_AGEMA_signal_4858 ;
    wire new_AGEMA_signal_4859 ;
    wire new_AGEMA_signal_4860 ;
    wire new_AGEMA_signal_4861 ;
    wire new_AGEMA_signal_4862 ;
    wire new_AGEMA_signal_4863 ;
    wire new_AGEMA_signal_4864 ;
    wire new_AGEMA_signal_4865 ;
    wire new_AGEMA_signal_4866 ;
    wire new_AGEMA_signal_4867 ;
    wire new_AGEMA_signal_4868 ;
    wire new_AGEMA_signal_4869 ;
    wire new_AGEMA_signal_4870 ;
    wire new_AGEMA_signal_4871 ;
    wire new_AGEMA_signal_4872 ;
    wire new_AGEMA_signal_4873 ;
    wire new_AGEMA_signal_4874 ;
    wire new_AGEMA_signal_4875 ;
    wire new_AGEMA_signal_4876 ;
    wire new_AGEMA_signal_4877 ;
    wire new_AGEMA_signal_4878 ;
    wire new_AGEMA_signal_4879 ;
    wire new_AGEMA_signal_4880 ;
    wire new_AGEMA_signal_4881 ;
    wire new_AGEMA_signal_4882 ;
    wire new_AGEMA_signal_4883 ;
    wire new_AGEMA_signal_4884 ;
    wire new_AGEMA_signal_4885 ;
    wire new_AGEMA_signal_4886 ;
    wire new_AGEMA_signal_4887 ;
    wire new_AGEMA_signal_4888 ;
    wire new_AGEMA_signal_4889 ;
    wire new_AGEMA_signal_4890 ;
    wire new_AGEMA_signal_4891 ;
    wire new_AGEMA_signal_4892 ;
    wire new_AGEMA_signal_4893 ;
    wire new_AGEMA_signal_4894 ;
    wire new_AGEMA_signal_4895 ;
    wire new_AGEMA_signal_4896 ;
    wire new_AGEMA_signal_4897 ;
    wire new_AGEMA_signal_4898 ;
    wire new_AGEMA_signal_4899 ;
    wire new_AGEMA_signal_4900 ;
    wire new_AGEMA_signal_4901 ;
    wire new_AGEMA_signal_4902 ;
    wire new_AGEMA_signal_4903 ;
    wire new_AGEMA_signal_4904 ;
    wire new_AGEMA_signal_4905 ;
    wire new_AGEMA_signal_4906 ;
    wire new_AGEMA_signal_4907 ;
    wire new_AGEMA_signal_4908 ;
    wire new_AGEMA_signal_4909 ;
    wire new_AGEMA_signal_4910 ;
    wire new_AGEMA_signal_4911 ;
    wire new_AGEMA_signal_4912 ;
    wire new_AGEMA_signal_4913 ;
    wire new_AGEMA_signal_4914 ;
    wire new_AGEMA_signal_4915 ;
    wire new_AGEMA_signal_4916 ;
    wire new_AGEMA_signal_4917 ;
    wire new_AGEMA_signal_4918 ;
    wire new_AGEMA_signal_4919 ;
    wire new_AGEMA_signal_4920 ;
    wire new_AGEMA_signal_4921 ;
    wire new_AGEMA_signal_4922 ;
    wire new_AGEMA_signal_4923 ;
    wire new_AGEMA_signal_4924 ;
    wire new_AGEMA_signal_4925 ;
    wire new_AGEMA_signal_4926 ;
    wire new_AGEMA_signal_4927 ;
    wire new_AGEMA_signal_4928 ;
    wire new_AGEMA_signal_4929 ;
    wire new_AGEMA_signal_4930 ;
    wire new_AGEMA_signal_4931 ;
    wire new_AGEMA_signal_4932 ;
    wire new_AGEMA_signal_4933 ;
    wire new_AGEMA_signal_4934 ;
    wire new_AGEMA_signal_4935 ;
    wire new_AGEMA_signal_4936 ;
    wire new_AGEMA_signal_4937 ;
    wire new_AGEMA_signal_4938 ;
    wire new_AGEMA_signal_4939 ;
    wire new_AGEMA_signal_4940 ;
    wire new_AGEMA_signal_4941 ;
    wire new_AGEMA_signal_4942 ;
    wire new_AGEMA_signal_4943 ;
    wire new_AGEMA_signal_4944 ;
    wire new_AGEMA_signal_4945 ;
    wire new_AGEMA_signal_4946 ;
    wire new_AGEMA_signal_4947 ;
    wire new_AGEMA_signal_4948 ;
    wire new_AGEMA_signal_4949 ;
    wire new_AGEMA_signal_4950 ;
    wire new_AGEMA_signal_4951 ;
    wire new_AGEMA_signal_4952 ;
    wire new_AGEMA_signal_4953 ;
    wire new_AGEMA_signal_4954 ;
    wire new_AGEMA_signal_4955 ;
    wire new_AGEMA_signal_4956 ;
    wire new_AGEMA_signal_4957 ;
    wire new_AGEMA_signal_4958 ;
    wire new_AGEMA_signal_4959 ;
    wire new_AGEMA_signal_4960 ;
    wire new_AGEMA_signal_4961 ;
    wire new_AGEMA_signal_4962 ;
    wire new_AGEMA_signal_4963 ;
    wire new_AGEMA_signal_4964 ;
    wire new_AGEMA_signal_4965 ;
    wire new_AGEMA_signal_4966 ;
    wire new_AGEMA_signal_4967 ;
    wire new_AGEMA_signal_4968 ;
    wire new_AGEMA_signal_4969 ;
    wire new_AGEMA_signal_4970 ;
    wire new_AGEMA_signal_4971 ;
    wire new_AGEMA_signal_4972 ;
    wire new_AGEMA_signal_4973 ;
    wire new_AGEMA_signal_4974 ;
    wire new_AGEMA_signal_4975 ;
    wire new_AGEMA_signal_4976 ;
    wire new_AGEMA_signal_4977 ;
    wire new_AGEMA_signal_4978 ;
    wire new_AGEMA_signal_4979 ;
    wire new_AGEMA_signal_4980 ;
    wire new_AGEMA_signal_4981 ;
    wire new_AGEMA_signal_4982 ;
    wire new_AGEMA_signal_4983 ;
    wire new_AGEMA_signal_4984 ;
    wire new_AGEMA_signal_4985 ;
    wire new_AGEMA_signal_4986 ;
    wire new_AGEMA_signal_4987 ;
    wire new_AGEMA_signal_4988 ;
    wire new_AGEMA_signal_4989 ;
    wire new_AGEMA_signal_4990 ;
    wire new_AGEMA_signal_4991 ;
    wire new_AGEMA_signal_4992 ;
    wire new_AGEMA_signal_4993 ;
    wire new_AGEMA_signal_4994 ;
    wire new_AGEMA_signal_4995 ;
    wire new_AGEMA_signal_4996 ;
    wire new_AGEMA_signal_4997 ;
    wire new_AGEMA_signal_4998 ;
    wire new_AGEMA_signal_4999 ;
    wire new_AGEMA_signal_5000 ;
    wire new_AGEMA_signal_5001 ;
    wire new_AGEMA_signal_5002 ;
    wire new_AGEMA_signal_5003 ;
    wire new_AGEMA_signal_5004 ;
    wire new_AGEMA_signal_5005 ;
    wire new_AGEMA_signal_5006 ;
    wire new_AGEMA_signal_5007 ;
    wire new_AGEMA_signal_5008 ;
    wire new_AGEMA_signal_5009 ;
    wire new_AGEMA_signal_5010 ;
    wire new_AGEMA_signal_5011 ;
    wire new_AGEMA_signal_5012 ;
    wire new_AGEMA_signal_5013 ;
    wire new_AGEMA_signal_5014 ;
    wire new_AGEMA_signal_5015 ;
    wire new_AGEMA_signal_5016 ;
    wire new_AGEMA_signal_5017 ;
    wire new_AGEMA_signal_5018 ;
    wire new_AGEMA_signal_5019 ;
    wire new_AGEMA_signal_5020 ;
    wire new_AGEMA_signal_5021 ;
    wire new_AGEMA_signal_5022 ;
    wire new_AGEMA_signal_5023 ;
    wire new_AGEMA_signal_5024 ;
    wire new_AGEMA_signal_5025 ;
    wire new_AGEMA_signal_5026 ;
    wire new_AGEMA_signal_5027 ;
    wire new_AGEMA_signal_5028 ;
    wire new_AGEMA_signal_5029 ;
    wire new_AGEMA_signal_5030 ;
    wire new_AGEMA_signal_5031 ;
    wire new_AGEMA_signal_5032 ;
    wire new_AGEMA_signal_5033 ;
    wire new_AGEMA_signal_5034 ;
    wire new_AGEMA_signal_5035 ;
    wire new_AGEMA_signal_5036 ;
    wire new_AGEMA_signal_5037 ;
    wire new_AGEMA_signal_5038 ;
    wire new_AGEMA_signal_5039 ;
    wire new_AGEMA_signal_5040 ;
    wire new_AGEMA_signal_5041 ;
    wire new_AGEMA_signal_5042 ;
    wire new_AGEMA_signal_5043 ;
    wire new_AGEMA_signal_5044 ;
    wire new_AGEMA_signal_5045 ;
    wire new_AGEMA_signal_5046 ;
    wire new_AGEMA_signal_5047 ;
    wire new_AGEMA_signal_5048 ;
    wire new_AGEMA_signal_5049 ;
    wire new_AGEMA_signal_5050 ;
    wire new_AGEMA_signal_5051 ;
    wire new_AGEMA_signal_5052 ;
    wire new_AGEMA_signal_5053 ;
    wire new_AGEMA_signal_5054 ;
    wire new_AGEMA_signal_5055 ;
    wire new_AGEMA_signal_5056 ;
    wire new_AGEMA_signal_5057 ;
    wire new_AGEMA_signal_5058 ;
    wire new_AGEMA_signal_5059 ;
    wire new_AGEMA_signal_5060 ;
    wire new_AGEMA_signal_5061 ;
    wire new_AGEMA_signal_5062 ;
    wire new_AGEMA_signal_5063 ;
    wire new_AGEMA_signal_5064 ;
    wire new_AGEMA_signal_5065 ;
    wire new_AGEMA_signal_5066 ;
    wire new_AGEMA_signal_5067 ;
    wire new_AGEMA_signal_5068 ;
    wire new_AGEMA_signal_5069 ;
    wire new_AGEMA_signal_5070 ;
    wire new_AGEMA_signal_5071 ;
    wire new_AGEMA_signal_5072 ;
    wire new_AGEMA_signal_5073 ;
    wire new_AGEMA_signal_5074 ;
    wire new_AGEMA_signal_5075 ;
    wire new_AGEMA_signal_5076 ;
    wire new_AGEMA_signal_5077 ;
    wire new_AGEMA_signal_5078 ;
    wire new_AGEMA_signal_5079 ;
    wire new_AGEMA_signal_5080 ;
    wire new_AGEMA_signal_5081 ;
    wire new_AGEMA_signal_5082 ;
    wire new_AGEMA_signal_5083 ;
    wire new_AGEMA_signal_5084 ;
    wire new_AGEMA_signal_5085 ;
    wire new_AGEMA_signal_5086 ;
    wire new_AGEMA_signal_5087 ;
    wire new_AGEMA_signal_5088 ;
    wire new_AGEMA_signal_5089 ;
    wire new_AGEMA_signal_5090 ;
    wire new_AGEMA_signal_5091 ;
    wire new_AGEMA_signal_5092 ;
    wire new_AGEMA_signal_5093 ;
    wire new_AGEMA_signal_5094 ;
    wire new_AGEMA_signal_5095 ;
    wire new_AGEMA_signal_5096 ;
    wire new_AGEMA_signal_5097 ;
    wire new_AGEMA_signal_5098 ;
    wire new_AGEMA_signal_5099 ;
    wire new_AGEMA_signal_5100 ;
    wire new_AGEMA_signal_5101 ;
    wire new_AGEMA_signal_5102 ;
    wire new_AGEMA_signal_5103 ;
    wire new_AGEMA_signal_5104 ;
    wire new_AGEMA_signal_5105 ;
    wire new_AGEMA_signal_5106 ;
    wire new_AGEMA_signal_5107 ;
    wire new_AGEMA_signal_5108 ;
    wire new_AGEMA_signal_5109 ;
    wire new_AGEMA_signal_5110 ;
    wire new_AGEMA_signal_5111 ;
    wire new_AGEMA_signal_5112 ;
    wire new_AGEMA_signal_5113 ;
    wire new_AGEMA_signal_5114 ;
    wire new_AGEMA_signal_5115 ;
    wire new_AGEMA_signal_5116 ;
    wire new_AGEMA_signal_5117 ;
    wire new_AGEMA_signal_5118 ;
    wire new_AGEMA_signal_5119 ;
    wire new_AGEMA_signal_5120 ;
    wire new_AGEMA_signal_5121 ;
    wire new_AGEMA_signal_5122 ;
    wire new_AGEMA_signal_5123 ;
    wire new_AGEMA_signal_5124 ;
    wire new_AGEMA_signal_5125 ;
    wire new_AGEMA_signal_5126 ;
    wire new_AGEMA_signal_5127 ;
    wire new_AGEMA_signal_5128 ;
    wire new_AGEMA_signal_5129 ;
    wire new_AGEMA_signal_5130 ;
    wire new_AGEMA_signal_5131 ;
    wire new_AGEMA_signal_5132 ;
    wire new_AGEMA_signal_5133 ;
    wire new_AGEMA_signal_5134 ;
    wire new_AGEMA_signal_5135 ;
    wire new_AGEMA_signal_5136 ;
    wire new_AGEMA_signal_5137 ;
    wire new_AGEMA_signal_5138 ;
    wire new_AGEMA_signal_5139 ;
    wire new_AGEMA_signal_5140 ;
    wire new_AGEMA_signal_5141 ;
    wire new_AGEMA_signal_5142 ;
    wire new_AGEMA_signal_5143 ;
    wire new_AGEMA_signal_5144 ;
    wire new_AGEMA_signal_5145 ;
    wire new_AGEMA_signal_5146 ;
    wire new_AGEMA_signal_5147 ;
    wire new_AGEMA_signal_5148 ;
    wire new_AGEMA_signal_5149 ;
    wire new_AGEMA_signal_5150 ;
    wire new_AGEMA_signal_5151 ;
    wire new_AGEMA_signal_5152 ;
    wire new_AGEMA_signal_5153 ;
    wire new_AGEMA_signal_5154 ;
    wire new_AGEMA_signal_5155 ;
    wire new_AGEMA_signal_5156 ;
    wire new_AGEMA_signal_5157 ;
    wire new_AGEMA_signal_5158 ;
    wire new_AGEMA_signal_5159 ;
    wire new_AGEMA_signal_5160 ;
    wire new_AGEMA_signal_5161 ;
    wire new_AGEMA_signal_5162 ;
    wire new_AGEMA_signal_5163 ;
    wire new_AGEMA_signal_5164 ;
    wire new_AGEMA_signal_5165 ;
    wire new_AGEMA_signal_5166 ;
    wire new_AGEMA_signal_5167 ;
    wire new_AGEMA_signal_5168 ;
    wire new_AGEMA_signal_5169 ;
    wire new_AGEMA_signal_5170 ;
    wire new_AGEMA_signal_5171 ;
    wire new_AGEMA_signal_5172 ;
    wire new_AGEMA_signal_5173 ;
    wire new_AGEMA_signal_5174 ;
    wire new_AGEMA_signal_5175 ;
    wire new_AGEMA_signal_5176 ;
    wire new_AGEMA_signal_5177 ;
    wire new_AGEMA_signal_5178 ;
    wire new_AGEMA_signal_5179 ;
    wire new_AGEMA_signal_5180 ;
    wire new_AGEMA_signal_5181 ;
    wire new_AGEMA_signal_5182 ;
    wire new_AGEMA_signal_5183 ;

    /* cells in depth 0 */
    INV_X1 U28 ( .A (selSR), .ZN (n12) ) ;
    linear_LMDPL #(.CONF(1'b0)) U29 ( .a ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, keyStateIn[0]}), .c ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, StateOutXORroundKey[0]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U30 ( .a ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .c ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, StateOutXORroundKey[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U31 ( .a ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, keyStateIn[2]}), .c ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, StateOutXORroundKey[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U32 ( .a ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, keyStateIn[3]}), .c ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, StateOutXORroundKey[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U33 ( .a ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[4]}), .c ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, StateOutXORroundKey[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U34 ( .a ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, keyStateIn[5]}), .c ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, StateOutXORroundKey[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U35 ( .a ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, keyStateIn[6]}), .c ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, StateOutXORroundKey[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) U36 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[7]}), .c ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, StateOutXORroundKey[7]}) ) ;
    NAND2_X1 U37 ( .A1 (intFinal), .A2 (finalStep), .ZN (n13) ) ;
    NOR2_X1 U38 ( .A1 (n10), .A2 (n13), .ZN (done) ) ;
    AND2_X1 U39 ( .A1 (notFirst), .A2 (selXOR), .ZN (intselXOR) ) ;
    INV_X1 U40 ( .A (start), .ZN (n9) ) ;
    NOR2_X1 ctrl_U20 ( .A1 (ctrl_n16), .A2 (ctrl_n4), .ZN (ctrl_nRstSeq4) ) ;
    XNOR2_X1 ctrl_U19 ( .A (ctrl_seq6Out_4_), .B (ctrl_seq6In_1_), .ZN (ctrl_n13) ) ;
    NOR2_X1 ctrl_U18 ( .A1 (ctrl_n15), .A2 (ctrl_n14), .ZN (finalStep) ) ;
    NAND2_X1 ctrl_U17 ( .A1 (ctrl_seq4In_1_), .A2 (ctrl_n2), .ZN (ctrl_n14) ) ;
    INV_X1 ctrl_U16 ( .A (ctrl_n16), .ZN (ctrl_n15) ) ;
    INV_X1 ctrl_U15 ( .A (ctrl_seq4Out_1_), .ZN (ctrl_n2) ) ;
    NAND2_X1 ctrl_U14 ( .A1 (ctrl_n11), .A2 (ctrl_n10), .ZN (ctrl_N14) ) ;
    NAND2_X1 ctrl_U13 ( .A1 (selXOR), .A2 (ctrl_n6), .ZN (ctrl_n11) ) ;
    NOR2_X1 ctrl_U12 ( .A1 (ctrl_seq6In_3_), .A2 (ctrl_seq6Out_4_), .ZN (ctrl_n7) ) ;
    NOR2_X1 ctrl_U11 ( .A1 (ctrl_seq6In_1_), .A2 (ctrl_seq6In_4_), .ZN (ctrl_n8) ) ;
    NOR2_X1 ctrl_U10 ( .A1 (ctrl_n4), .A2 (ctrl_n5), .ZN (selXOR) ) ;
    NOR2_X1 ctrl_U9 ( .A1 (ctrl_seq4Out_1_), .A2 (ctrl_seq4In_1_), .ZN (ctrl_n5) ) ;
    INV_X1 ctrl_U8 ( .A (nReset), .ZN (ctrl_n4) ) ;
    NAND2_X1 ctrl_U7 ( .A1 (ctrl_n8), .A2 (ctrl_n7), .ZN (ctrl_n9) ) ;
    NOR2_X1 ctrl_U6 ( .A1 (ctrl_seq6In_2_), .A2 (ctrl_n9), .ZN (ctrl_n16) ) ;
    NAND2_X1 ctrl_U5 ( .A1 (nReset), .A2 (ctrl_n16), .ZN (ctrl_n10) ) ;
    INV_X1 ctrl_U4 ( .A (ctrl_n10), .ZN (selSR) ) ;
    NOR2_X1 ctrl_U3 ( .A1 (ctrl_n12), .A2 (ctrl_n4), .ZN (selMC) ) ;
    MUX2_X1 ctrl_seq6_SFF_0_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_n13), .Z (ctrl_seq6_SFF_0_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_1_MUXInst_U1 ( .S (nReset), .A (1'b0), .B (ctrl_seq6In_1_), .Z (ctrl_seq6_SFF_1_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_2_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_seq6In_2_), .Z (ctrl_seq6_SFF_2_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_3_MUXInst_U1 ( .S (nReset), .A (1'b0), .B (ctrl_seq6In_3_), .Z (ctrl_seq6_SFF_3_QD) ) ;
    MUX2_X1 ctrl_seq6_SFF_4_MUXInst_U1 ( .S (nReset), .A (1'b1), .B (ctrl_seq6In_4_), .Z (ctrl_seq6_SFF_4_QD) ) ;
    MUX2_X1 ctrl_seq4_SFF_0_MUXInst_U1 ( .S (ctrl_nRstSeq4), .A (1'b1), .B (ctrl_n2), .Z (ctrl_seq4_SFF_0_QD) ) ;
    MUX2_X1 ctrl_seq4_SFF_1_MUXInst_U1 ( .S (ctrl_nRstSeq4), .A (1'b0), .B (ctrl_seq4In_1_), .Z (ctrl_seq4_SFF_1_QD) ) ;
    INV_X1 ctrl_CSselMC_reg_U1 ( .A (ctrl_n6), .ZN (ctrl_n12) ) ;
    mux2_masked_LMDPL MUX_StateIn_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, SboxOut[0]}), .a ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, StateOutXORroundKey[0]}), .c ({new_AGEMA_signal_5027, new_AGEMA_signal_5026, StateIn[0]}) ) ;
    mux2_masked_LMDPL MUX_StateIn_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, SboxOut[1]}), .a ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, StateOutXORroundKey[1]}), .c ({new_AGEMA_signal_5045, new_AGEMA_signal_5044, StateIn[1]}) ) ;
    mux2_masked_LMDPL MUX_StateIn_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, SboxOut[2]}), .a ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, StateOutXORroundKey[2]}), .c ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, StateIn[2]}) ) ;
    mux2_masked_LMDPL MUX_StateIn_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, SboxOut[3]}), .a ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, StateOutXORroundKey[3]}), .c ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, StateIn[3]}) ) ;
    mux2_masked_LMDPL MUX_StateIn_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, SboxOut[4]}), .a ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, StateOutXORroundKey[4]}), .c ({new_AGEMA_signal_5051, new_AGEMA_signal_5050, StateIn[4]}) ) ;
    mux2_masked_LMDPL MUX_StateIn_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, SboxOut[5]}), .a ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, StateOutXORroundKey[5]}), .c ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, StateIn[5]}) ) ;
    mux2_masked_LMDPL MUX_StateIn_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, SboxOut[6]}), .a ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, StateOutXORroundKey[6]}), .c ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, StateIn[6]}) ) ;
    mux2_masked_LMDPL MUX_StateIn_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, SboxOut[7]}), .a ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, StateOutXORroundKey[7]}), .c ({new_AGEMA_signal_5057, new_AGEMA_signal_5056, StateIn[7]}) ) ;
    INV_X1 stateArray_U21 ( .A (selMC), .ZN (stateArray_n24) ) ;
    INV_X1 stateArray_U20 ( .A (stateArray_n24), .ZN (stateArray_n22) ) ;
    INV_X1 stateArray_U19 ( .A (nReset), .ZN (stateArray_n33) ) ;
    INV_X1 stateArray_U18 ( .A (stateArray_n33), .ZN (stateArray_n25) ) ;
    INV_X1 stateArray_U17 ( .A (stateArray_n21), .ZN (stateArray_n13) ) ;
    INV_X1 stateArray_U16 ( .A (stateArray_n24), .ZN (stateArray_n23) ) ;
    INV_X1 stateArray_U15 ( .A (stateArray_n33), .ZN (stateArray_n29) ) ;
    INV_X1 stateArray_U14 ( .A (stateArray_n21), .ZN (stateArray_n17) ) ;
    INV_X1 stateArray_U13 ( .A (stateArray_n33), .ZN (stateArray_n31) ) ;
    INV_X1 stateArray_U12 ( .A (stateArray_n21), .ZN (stateArray_n19) ) ;
    INV_X1 stateArray_U11 ( .A (stateArray_n33), .ZN (stateArray_n27) ) ;
    INV_X1 stateArray_U10 ( .A (stateArray_n21), .ZN (stateArray_n15) ) ;
    INV_X1 stateArray_U9 ( .A (stateArray_n33), .ZN (stateArray_n32) ) ;
    INV_X1 stateArray_U8 ( .A (stateArray_n21), .ZN (stateArray_n20) ) ;
    INV_X1 stateArray_U7 ( .A (stateArray_n33), .ZN (stateArray_n30) ) ;
    INV_X1 stateArray_U6 ( .A (stateArray_n21), .ZN (stateArray_n18) ) ;
    INV_X1 stateArray_U5 ( .A (stateArray_n33), .ZN (stateArray_n28) ) ;
    INV_X1 stateArray_U4 ( .A (stateArray_n21), .ZN (stateArray_n16) ) ;
    INV_X1 stateArray_U3 ( .A (stateArray_n33), .ZN (stateArray_n26) ) ;
    INV_X1 stateArray_U2 ( .A (stateArray_n21), .ZN (stateArray_n14) ) ;
    INV_X1 stateArray_U1 ( .A (selSR), .ZN (stateArray_n21) ) ;
    mux2_masked_LMDPL stateArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, stateArray_inS00ser[0]}), .a ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, stateArray_S00reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, stateArray_inS00ser[1]}), .a ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_4343, new_AGEMA_signal_4342, stateArray_S00reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, stateArray_inS00ser[2]}), .a ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, stateArray_S00reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, stateArray_inS00ser[3]}), .a ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, stateArray_S00reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, stateArray_inS00ser[4]}), .a ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_4349, new_AGEMA_signal_4348, stateArray_S00reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, stateArray_inS00ser[5]}), .a ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_4351, new_AGEMA_signal_4350, stateArray_S00reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, stateArray_inS00ser[6]}), .a ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, stateArray_S00reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, stateArray_inS00ser[7]}), .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, stateArray_S00reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, stateArray_inS01ser[0]}), .a ({new_AGEMA_signal_2335, ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, stateArray_S01reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, stateArray_inS01ser[1]}), .a ({new_AGEMA_signal_2341, ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, stateArray_S01reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, stateArray_inS01ser[2]}), .a ({new_AGEMA_signal_2347, ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, stateArray_S01reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, stateArray_inS01ser[3]}), .a ({new_AGEMA_signal_2353, ciphertext_s1[115], ciphertext_s0[115]}), .c ({new_AGEMA_signal_4363, new_AGEMA_signal_4362, stateArray_S01reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, stateArray_inS01ser[4]}), .a ({new_AGEMA_signal_2359, ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, stateArray_S01reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, stateArray_inS01ser[5]}), .a ({new_AGEMA_signal_2365, ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_4367, new_AGEMA_signal_4366, stateArray_S01reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, stateArray_inS01ser[6]}), .a ({new_AGEMA_signal_2371, ciphertext_s1[118], ciphertext_s0[118]}), .c ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, stateArray_S01reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4339, new_AGEMA_signal_4338, stateArray_n20}), .b ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, stateArray_inS01ser[7]}), .a ({new_AGEMA_signal_2377, ciphertext_s1[119], ciphertext_s0[119]}), .c ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, stateArray_S01reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, stateArray_inS02ser[0]}), .a ({new_AGEMA_signal_2383, ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_4375, new_AGEMA_signal_4374, stateArray_S02reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, stateArray_inS02ser[1]}), .a ({new_AGEMA_signal_2389, ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, stateArray_S02reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, stateArray_inS02ser[2]}), .a ({new_AGEMA_signal_2395, ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_4379, new_AGEMA_signal_4378, stateArray_S02reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, stateArray_inS02ser[3]}), .a ({new_AGEMA_signal_2401, ciphertext_s1[107], ciphertext_s0[107]}), .c ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, stateArray_S02reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, stateArray_inS02ser[4]}), .a ({new_AGEMA_signal_2407, ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, stateArray_S02reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, stateArray_inS02ser[5]}), .a ({new_AGEMA_signal_2413, ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, stateArray_S02reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, stateArray_inS02ser[6]}), .a ({new_AGEMA_signal_2419, ciphertext_s1[110], ciphertext_s0[110]}), .c ({new_AGEMA_signal_4387, new_AGEMA_signal_4386, stateArray_S02reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, stateArray_inS02ser[7]}), .a ({new_AGEMA_signal_2425, ciphertext_s1[111], ciphertext_s0[111]}), .c ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, stateArray_S02reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_4175, new_AGEMA_signal_4174, stateArray_inS03ser[0]}), .a ({new_AGEMA_signal_2433, ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_4391, new_AGEMA_signal_4390, stateArray_S03reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, stateArray_inS03ser[1]}), .a ({new_AGEMA_signal_2439, ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, stateArray_S03reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_4183, new_AGEMA_signal_4182, stateArray_inS03ser[2]}), .a ({new_AGEMA_signal_2445, ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, stateArray_S03reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_4187, new_AGEMA_signal_4186, stateArray_inS03ser[3]}), .a ({new_AGEMA_signal_2451, ciphertext_s1[99], ciphertext_s0[99]}), .c ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, stateArray_S03reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, stateArray_inS03ser[4]}), .a ({new_AGEMA_signal_2457, ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, stateArray_S03reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, stateArray_inS03ser[5]}), .a ({new_AGEMA_signal_2463, ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, stateArray_S03reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_4199, new_AGEMA_signal_4198, stateArray_inS03ser[6]}), .a ({new_AGEMA_signal_2469, ciphertext_s1[102], ciphertext_s0[102]}), .c ({new_AGEMA_signal_4403, new_AGEMA_signal_4402, stateArray_S03reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4373, new_AGEMA_signal_4372, stateArray_n19}), .b ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, stateArray_inS03ser[7]}), .a ({new_AGEMA_signal_2475, ciphertext_s1[103], ciphertext_s0[103]}), .c ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, stateArray_S03reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, stateArray_inS10ser[0]}), .a ({new_AGEMA_signal_2483, ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, stateArray_S10reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, stateArray_inS10ser[1]}), .a ({new_AGEMA_signal_2489, ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, stateArray_S10reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, stateArray_inS10ser[2]}), .a ({new_AGEMA_signal_2495, ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, stateArray_S10reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, stateArray_inS10ser[3]}), .a ({new_AGEMA_signal_2501, ciphertext_s1[83], ciphertext_s0[83]}), .c ({new_AGEMA_signal_4415, new_AGEMA_signal_4414, stateArray_S10reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, stateArray_inS10ser[4]}), .a ({new_AGEMA_signal_2507, ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, stateArray_S10reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, stateArray_inS10ser[5]}), .a ({new_AGEMA_signal_2513, ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, stateArray_S10reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, stateArray_inS10ser[6]}), .a ({new_AGEMA_signal_2519, ciphertext_s1[86], ciphertext_s0[86]}), .c ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, stateArray_S10reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, stateArray_inS10ser[7]}), .a ({new_AGEMA_signal_2525, ciphertext_s1[87], ciphertext_s0[87]}), .c ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, stateArray_S10reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, stateArray_inS11ser[0]}), .a ({new_AGEMA_signal_2531, ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, stateArray_S11reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, stateArray_inS11ser[1]}), .a ({new_AGEMA_signal_2537, ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_4427, new_AGEMA_signal_4426, stateArray_S11reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, stateArray_inS11ser[2]}), .a ({new_AGEMA_signal_2543, ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, stateArray_S11reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, stateArray_inS11ser[3]}), .a ({new_AGEMA_signal_2549, ciphertext_s1[75], ciphertext_s0[75]}), .c ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, stateArray_S11reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, stateArray_inS11ser[4]}), .a ({new_AGEMA_signal_2555, ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, stateArray_S11reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, stateArray_inS11ser[5]}), .a ({new_AGEMA_signal_2561, ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, stateArray_S11reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, stateArray_inS11ser[6]}), .a ({new_AGEMA_signal_2567, ciphertext_s1[78], ciphertext_s0[78]}), .c ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, stateArray_S11reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4407, new_AGEMA_signal_4406, stateArray_n18}), .b ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, stateArray_inS11ser[7]}), .a ({new_AGEMA_signal_2573, ciphertext_s1[79], ciphertext_s0[79]}), .c ({new_AGEMA_signal_4439, new_AGEMA_signal_4438, stateArray_S11reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, stateArray_inS12ser[0]}), .a ({new_AGEMA_signal_2581, ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, stateArray_S12reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, stateArray_inS12ser[1]}), .a ({new_AGEMA_signal_2587, ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, stateArray_S12reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, stateArray_inS12ser[2]}), .a ({new_AGEMA_signal_2593, ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, stateArray_S12reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, stateArray_inS12ser[3]}), .a ({new_AGEMA_signal_2599, ciphertext_s1[67], ciphertext_s0[67]}), .c ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, stateArray_S12reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, stateArray_inS12ser[4]}), .a ({new_AGEMA_signal_2605, ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_4451, new_AGEMA_signal_4450, stateArray_S12reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, stateArray_inS12ser[5]}), .a ({new_AGEMA_signal_2611, ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, stateArray_S12reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, stateArray_inS12ser[6]}), .a ({new_AGEMA_signal_2617, ciphertext_s1[70], ciphertext_s0[70]}), .c ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, stateArray_S12reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, stateArray_inS12ser[7]}), .a ({new_AGEMA_signal_2623, ciphertext_s1[71], ciphertext_s0[71]}), .c ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, stateArray_S12reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_4207, new_AGEMA_signal_4206, stateArray_inS13ser[0]}), .a ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, stateArray_S13reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_4211, new_AGEMA_signal_4210, stateArray_inS13ser[1]}), .a ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, stateArray_S13reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, stateArray_inS13ser[2]}), .a ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_4463, new_AGEMA_signal_4462, stateArray_S13reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_4219, new_AGEMA_signal_4218, stateArray_inS13ser[3]}), .a ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, stateArray_S13reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_4223, new_AGEMA_signal_4222, stateArray_inS13ser[4]}), .a ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, stateArray_S13reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, stateArray_inS13ser[5]}), .a ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, stateArray_S13reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, stateArray_inS13ser[6]}), .a ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, stateArray_S13reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4441, new_AGEMA_signal_4440, stateArray_n17}), .b ({new_AGEMA_signal_4235, new_AGEMA_signal_4234, stateArray_inS13ser[7]}), .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, stateArray_S13reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, stateArray_inS20ser[0]}), .a ({new_AGEMA_signal_2679, ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, stateArray_S20reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, stateArray_inS20ser[1]}), .a ({new_AGEMA_signal_2685, ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, stateArray_S20reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, stateArray_inS20ser[2]}), .a ({new_AGEMA_signal_2691, ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, stateArray_S20reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, stateArray_inS20ser[3]}), .a ({new_AGEMA_signal_2697, ciphertext_s1[43], ciphertext_s0[43]}), .c ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, stateArray_S20reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, stateArray_inS20ser[4]}), .a ({new_AGEMA_signal_2703, ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, stateArray_S20reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, stateArray_inS20ser[5]}), .a ({new_AGEMA_signal_2709, ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_4487, new_AGEMA_signal_4486, stateArray_S20reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, stateArray_inS20ser[6]}), .a ({new_AGEMA_signal_2715, ciphertext_s1[46], ciphertext_s0[46]}), .c ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, stateArray_S20reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, stateArray_inS20ser[7]}), .a ({new_AGEMA_signal_2721, ciphertext_s1[47], ciphertext_s0[47]}), .c ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, stateArray_S20reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, stateArray_inS21ser[0]}), .a ({new_AGEMA_signal_2729, ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_4493, new_AGEMA_signal_4492, stateArray_S21reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, stateArray_inS21ser[1]}), .a ({new_AGEMA_signal_2735, ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, stateArray_S21reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, stateArray_inS21ser[2]}), .a ({new_AGEMA_signal_2741, ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, stateArray_S21reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, stateArray_inS21ser[3]}), .a ({new_AGEMA_signal_2747, ciphertext_s1[35], ciphertext_s0[35]}), .c ({new_AGEMA_signal_4499, new_AGEMA_signal_4498, stateArray_S21reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, stateArray_inS21ser[4]}), .a ({new_AGEMA_signal_2753, ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, stateArray_S21reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, stateArray_inS21ser[5]}), .a ({new_AGEMA_signal_2759, ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, stateArray_S21reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, stateArray_inS21ser[6]}), .a ({new_AGEMA_signal_2765, ciphertext_s1[38], ciphertext_s0[38]}), .c ({new_AGEMA_signal_4505, new_AGEMA_signal_4504, stateArray_S21reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4475, new_AGEMA_signal_4474, stateArray_n16}), .b ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, stateArray_inS21ser[7]}), .a ({new_AGEMA_signal_2771, ciphertext_s1[39], ciphertext_s0[39]}), .c ({new_AGEMA_signal_4507, new_AGEMA_signal_4506, stateArray_S21reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, stateArray_inS22ser[0]}), .a ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_4511, new_AGEMA_signal_4510, stateArray_S22reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, stateArray_inS22ser[1]}), .a ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, stateArray_S22reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, stateArray_inS22ser[2]}), .a ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, stateArray_S22reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, stateArray_inS22ser[3]}), .a ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, stateArray_S22reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, stateArray_inS22ser[4]}), .a ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, stateArray_S22reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, stateArray_inS22ser[5]}), .a ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, stateArray_S22reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, stateArray_inS22ser[6]}), .a ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_4523, new_AGEMA_signal_4522, stateArray_S22reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, stateArray_inS22ser[7]}), .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, stateArray_S22reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, stateArray_inS23ser[0]}), .a ({new_AGEMA_signal_2631, ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, stateArray_S23reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_4243, new_AGEMA_signal_4242, stateArray_inS23ser[1]}), .a ({new_AGEMA_signal_2637, ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_4529, new_AGEMA_signal_4528, stateArray_S23reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_4247, new_AGEMA_signal_4246, stateArray_inS23ser[2]}), .a ({new_AGEMA_signal_2643, ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, stateArray_S23reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, stateArray_inS23ser[3]}), .a ({new_AGEMA_signal_2649, ciphertext_s1[51], ciphertext_s0[51]}), .c ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, stateArray_S23reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, stateArray_inS23ser[4]}), .a ({new_AGEMA_signal_2655, ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_4535, new_AGEMA_signal_4534, stateArray_S23reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, stateArray_inS23ser[5]}), .a ({new_AGEMA_signal_2661, ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, stateArray_S23reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, stateArray_inS23ser[6]}), .a ({new_AGEMA_signal_2667, ciphertext_s1[54], ciphertext_s0[54]}), .c ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, stateArray_S23reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4509, new_AGEMA_signal_4508, stateArray_n15}), .b ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, stateArray_inS23ser[7]}), .a ({new_AGEMA_signal_2673, ciphertext_s1[55], ciphertext_s0[55]}), .c ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, stateArray_S23reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, stateArray_inS30ser[0]}), .a ({new_AGEMA_signal_2877, ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, stateArray_S30reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, stateArray_inS30ser[1]}), .a ({new_AGEMA_signal_2883, ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_4547, new_AGEMA_signal_4546, stateArray_S30reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, stateArray_inS30ser[2]}), .a ({new_AGEMA_signal_2889, ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, stateArray_S30reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, stateArray_inS30ser[3]}), .a ({new_AGEMA_signal_2895, ciphertext_s1[3], ciphertext_s0[3]}), .c ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, stateArray_S30reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, stateArray_inS30ser[4]}), .a ({new_AGEMA_signal_2901, ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_4553, new_AGEMA_signal_4552, stateArray_S30reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, stateArray_inS30ser[5]}), .a ({new_AGEMA_signal_2907, ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, stateArray_S30reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, stateArray_inS30ser[6]}), .a ({new_AGEMA_signal_2913, ciphertext_s1[6], ciphertext_s0[6]}), .c ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, stateArray_S30reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, stateArray_inS30ser[7]}), .a ({new_AGEMA_signal_2919, ciphertext_s1[7], ciphertext_s0[7]}), .c ({new_AGEMA_signal_4559, new_AGEMA_signal_4558, stateArray_S30reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, stateArray_inS31ser[0]}), .a ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, stateArray_S31reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, stateArray_inS31ser[1]}), .a ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, stateArray_S31reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, stateArray_inS31ser[2]}), .a ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, stateArray_S31reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, stateArray_inS31ser[3]}), .a ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_4567, new_AGEMA_signal_4566, stateArray_S31reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, stateArray_inS31ser[4]}), .a ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, stateArray_S31reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, stateArray_inS31ser[5]}), .a ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_4571, new_AGEMA_signal_4570, stateArray_S31reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, stateArray_inS31ser[6]}), .a ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, stateArray_S31reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4543, new_AGEMA_signal_4542, stateArray_n14}), .b ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, stateArray_inS31ser[7]}), .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, stateArray_S31reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, stateArray_inS32ser[0]}), .a ({new_AGEMA_signal_2779, ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, stateArray_S32reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, stateArray_inS32ser[1]}), .a ({new_AGEMA_signal_2785, ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, stateArray_S32reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, stateArray_inS32ser[2]}), .a ({new_AGEMA_signal_2791, ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_4583, new_AGEMA_signal_4582, stateArray_S32reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, stateArray_inS32ser[3]}), .a ({new_AGEMA_signal_2797, ciphertext_s1[19], ciphertext_s0[19]}), .c ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, stateArray_S32reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, stateArray_inS32ser[4]}), .a ({new_AGEMA_signal_2803, ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, stateArray_S32reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, stateArray_inS32ser[5]}), .a ({new_AGEMA_signal_2809, ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_4589, new_AGEMA_signal_4588, stateArray_S32reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, stateArray_inS32ser[6]}), .a ({new_AGEMA_signal_2815, ciphertext_s1[22], ciphertext_s0[22]}), .c ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, stateArray_S32reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, stateArray_inS32ser[7]}), .a ({new_AGEMA_signal_2821, ciphertext_s1[23], ciphertext_s0[23]}), .c ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, stateArray_S32reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_5093, new_AGEMA_signal_5092, stateArray_inS33ser[0]}), .a ({new_AGEMA_signal_2827, ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_5111, new_AGEMA_signal_5110, stateArray_S33reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL stateArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, stateArray_inS33ser[1]}), .a ({new_AGEMA_signal_2833, ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, stateArray_S33reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL stateArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_5119, new_AGEMA_signal_5118, stateArray_inS33ser[2]}), .a ({new_AGEMA_signal_2839, ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_5159, new_AGEMA_signal_5158, stateArray_S33reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL stateArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_5123, new_AGEMA_signal_5122, stateArray_inS33ser[3]}), .a ({new_AGEMA_signal_2845, ciphertext_s1[11], ciphertext_s0[11]}), .c ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, stateArray_S33reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL stateArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, stateArray_inS33ser[4]}), .a ({new_AGEMA_signal_2851, ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, stateArray_S33reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL stateArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_5131, new_AGEMA_signal_5130, stateArray_inS33ser[5]}), .a ({new_AGEMA_signal_2857, ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_5165, new_AGEMA_signal_5164, stateArray_S33reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL stateArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_5135, new_AGEMA_signal_5134, stateArray_inS33ser[6]}), .a ({new_AGEMA_signal_2863, ciphertext_s1[14], ciphertext_s0[14]}), .c ({new_AGEMA_signal_5167, new_AGEMA_signal_5166, stateArray_S33reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL stateArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4577, new_AGEMA_signal_4576, stateArray_n13}), .b ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, stateArray_inS33ser[7]}), .a ({new_AGEMA_signal_2869, ciphertext_s1[15], ciphertext_s0[15]}), .c ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, stateArray_S33reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS00ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2333, new_AGEMA_signal_2332, plaintext_s0[120]}), .a ({new_AGEMA_signal_2335, ciphertext_s1[112], ciphertext_s0[112]}), .c ({new_AGEMA_signal_2337, new_AGEMA_signal_2336, stateArray_inS00ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS00ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2339, new_AGEMA_signal_2338, plaintext_s0[121]}), .a ({new_AGEMA_signal_2341, ciphertext_s1[113], ciphertext_s0[113]}), .c ({new_AGEMA_signal_2343, new_AGEMA_signal_2342, stateArray_inS00ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS00ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2345, new_AGEMA_signal_2344, plaintext_s0[122]}), .a ({new_AGEMA_signal_2347, ciphertext_s1[114], ciphertext_s0[114]}), .c ({new_AGEMA_signal_2349, new_AGEMA_signal_2348, stateArray_inS00ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS00ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2351, new_AGEMA_signal_2350, plaintext_s0[123]}), .a ({new_AGEMA_signal_2353, ciphertext_s1[115], ciphertext_s0[115]}), .c ({new_AGEMA_signal_2355, new_AGEMA_signal_2354, stateArray_inS00ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS00ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2357, new_AGEMA_signal_2356, plaintext_s0[124]}), .a ({new_AGEMA_signal_2359, ciphertext_s1[116], ciphertext_s0[116]}), .c ({new_AGEMA_signal_2361, new_AGEMA_signal_2360, stateArray_inS00ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS00ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2363, new_AGEMA_signal_2362, plaintext_s0[125]}), .a ({new_AGEMA_signal_2365, ciphertext_s1[117], ciphertext_s0[117]}), .c ({new_AGEMA_signal_2367, new_AGEMA_signal_2366, stateArray_inS00ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS00ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2369, new_AGEMA_signal_2368, plaintext_s0[126]}), .a ({new_AGEMA_signal_2371, ciphertext_s1[118], ciphertext_s0[118]}), .c ({new_AGEMA_signal_2373, new_AGEMA_signal_2372, stateArray_inS00ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS00ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2375, new_AGEMA_signal_2374, plaintext_s0[127]}), .a ({new_AGEMA_signal_2377, ciphertext_s1[119], ciphertext_s0[119]}), .c ({new_AGEMA_signal_2379, new_AGEMA_signal_2378, stateArray_inS00ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS01ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2381, new_AGEMA_signal_2380, plaintext_s0[112]}), .a ({new_AGEMA_signal_2383, ciphertext_s1[104], ciphertext_s0[104]}), .c ({new_AGEMA_signal_2385, new_AGEMA_signal_2384, stateArray_inS01ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS01ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2387, new_AGEMA_signal_2386, plaintext_s0[113]}), .a ({new_AGEMA_signal_2389, ciphertext_s1[105], ciphertext_s0[105]}), .c ({new_AGEMA_signal_2391, new_AGEMA_signal_2390, stateArray_inS01ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS01ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2393, new_AGEMA_signal_2392, plaintext_s0[114]}), .a ({new_AGEMA_signal_2395, ciphertext_s1[106], ciphertext_s0[106]}), .c ({new_AGEMA_signal_2397, new_AGEMA_signal_2396, stateArray_inS01ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS01ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2399, new_AGEMA_signal_2398, plaintext_s0[115]}), .a ({new_AGEMA_signal_2401, ciphertext_s1[107], ciphertext_s0[107]}), .c ({new_AGEMA_signal_2403, new_AGEMA_signal_2402, stateArray_inS01ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS01ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2405, new_AGEMA_signal_2404, plaintext_s0[116]}), .a ({new_AGEMA_signal_2407, ciphertext_s1[108], ciphertext_s0[108]}), .c ({new_AGEMA_signal_2409, new_AGEMA_signal_2408, stateArray_inS01ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS01ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2411, new_AGEMA_signal_2410, plaintext_s0[117]}), .a ({new_AGEMA_signal_2413, ciphertext_s1[109], ciphertext_s0[109]}), .c ({new_AGEMA_signal_2415, new_AGEMA_signal_2414, stateArray_inS01ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS01ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2417, new_AGEMA_signal_2416, plaintext_s0[118]}), .a ({new_AGEMA_signal_2419, ciphertext_s1[110], ciphertext_s0[110]}), .c ({new_AGEMA_signal_2421, new_AGEMA_signal_2420, stateArray_inS01ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS01ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2331, new_AGEMA_signal_2330, stateArray_n32}), .b ({new_AGEMA_signal_2423, new_AGEMA_signal_2422, plaintext_s0[119]}), .a ({new_AGEMA_signal_2425, ciphertext_s1[111], ciphertext_s0[111]}), .c ({new_AGEMA_signal_2427, new_AGEMA_signal_2426, stateArray_inS01ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS02ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_2431, new_AGEMA_signal_2430, plaintext_s0[104]}), .a ({new_AGEMA_signal_2433, ciphertext_s1[96], ciphertext_s0[96]}), .c ({new_AGEMA_signal_2435, new_AGEMA_signal_2434, stateArray_inS02ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS02ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_2437, new_AGEMA_signal_2436, plaintext_s0[105]}), .a ({new_AGEMA_signal_2439, ciphertext_s1[97], ciphertext_s0[97]}), .c ({new_AGEMA_signal_2441, new_AGEMA_signal_2440, stateArray_inS02ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS02ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_2443, new_AGEMA_signal_2442, plaintext_s0[106]}), .a ({new_AGEMA_signal_2445, ciphertext_s1[98], ciphertext_s0[98]}), .c ({new_AGEMA_signal_2447, new_AGEMA_signal_2446, stateArray_inS02ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS02ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_2449, new_AGEMA_signal_2448, plaintext_s0[107]}), .a ({new_AGEMA_signal_2451, ciphertext_s1[99], ciphertext_s0[99]}), .c ({new_AGEMA_signal_2453, new_AGEMA_signal_2452, stateArray_inS02ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS02ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_2455, new_AGEMA_signal_2454, plaintext_s0[108]}), .a ({new_AGEMA_signal_2457, ciphertext_s1[100], ciphertext_s0[100]}), .c ({new_AGEMA_signal_2459, new_AGEMA_signal_2458, stateArray_inS02ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS02ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_2461, new_AGEMA_signal_2460, plaintext_s0[109]}), .a ({new_AGEMA_signal_2463, ciphertext_s1[101], ciphertext_s0[101]}), .c ({new_AGEMA_signal_2465, new_AGEMA_signal_2464, stateArray_inS02ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS02ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_2467, new_AGEMA_signal_2466, plaintext_s0[110]}), .a ({new_AGEMA_signal_2469, ciphertext_s1[102], ciphertext_s0[102]}), .c ({new_AGEMA_signal_2471, new_AGEMA_signal_2470, stateArray_inS02ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS02ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_2473, new_AGEMA_signal_2472, plaintext_s0[111]}), .a ({new_AGEMA_signal_2475, ciphertext_s1[103], ciphertext_s0[103]}), .c ({new_AGEMA_signal_2477, new_AGEMA_signal_2476, stateArray_inS02ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS10_MC_mux_inst_0_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}), .a ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, StateInMC[24]}), .c ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, stateArray_outS10ser_MC[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS10_MC_mux_inst_1_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}), .a ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, StateInMC[25]}), .c ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, stateArray_outS10ser_MC[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS10_MC_mux_inst_2_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}), .a ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, StateInMC[26]}), .c ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, stateArray_outS10ser_MC[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS10_MC_mux_inst_3_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}), .a ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, StateInMC[27]}), .c ({new_AGEMA_signal_4103, new_AGEMA_signal_4102, stateArray_outS10ser_MC[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS10_MC_mux_inst_4_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}), .a ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, StateInMC[28]}), .c ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, stateArray_outS10ser_MC[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS10_MC_mux_inst_5_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}), .a ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, StateInMC[29]}), .c ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, stateArray_outS10ser_MC[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS10_MC_mux_inst_6_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}), .a ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, StateInMC[30]}), .c ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, stateArray_outS10ser_MC[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS10_MC_mux_inst_7_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .a ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, StateInMC[31]}), .c ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, stateArray_outS10ser_MC[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS03ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_4173, new_AGEMA_signal_4172, plaintext_s0[96]}), .a ({new_AGEMA_signal_4097, new_AGEMA_signal_4096, stateArray_outS10ser_MC[0]}), .c ({new_AGEMA_signal_4175, new_AGEMA_signal_4174, stateArray_inS03ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS03ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_4177, new_AGEMA_signal_4176, plaintext_s0[97]}), .a ({new_AGEMA_signal_4099, new_AGEMA_signal_4098, stateArray_outS10ser_MC[1]}), .c ({new_AGEMA_signal_4179, new_AGEMA_signal_4178, stateArray_inS03ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS03ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_4181, new_AGEMA_signal_4180, plaintext_s0[98]}), .a ({new_AGEMA_signal_4101, new_AGEMA_signal_4100, stateArray_outS10ser_MC[2]}), .c ({new_AGEMA_signal_4183, new_AGEMA_signal_4182, stateArray_inS03ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS03ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_4185, new_AGEMA_signal_4184, plaintext_s0[99]}), .a ({new_AGEMA_signal_4103, new_AGEMA_signal_4102, stateArray_outS10ser_MC[3]}), .c ({new_AGEMA_signal_4187, new_AGEMA_signal_4186, stateArray_inS03ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS03ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_4189, new_AGEMA_signal_4188, plaintext_s0[100]}), .a ({new_AGEMA_signal_4105, new_AGEMA_signal_4104, stateArray_outS10ser_MC[4]}), .c ({new_AGEMA_signal_4191, new_AGEMA_signal_4190, stateArray_inS03ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS03ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_4193, new_AGEMA_signal_4192, plaintext_s0[101]}), .a ({new_AGEMA_signal_4107, new_AGEMA_signal_4106, stateArray_outS10ser_MC[5]}), .c ({new_AGEMA_signal_4195, new_AGEMA_signal_4194, stateArray_inS03ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS03ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_4197, new_AGEMA_signal_4196, plaintext_s0[102]}), .a ({new_AGEMA_signal_4109, new_AGEMA_signal_4108, stateArray_outS10ser_MC[6]}), .c ({new_AGEMA_signal_4199, new_AGEMA_signal_4198, stateArray_inS03ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS03ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2429, new_AGEMA_signal_2428, stateArray_n31}), .b ({new_AGEMA_signal_4201, new_AGEMA_signal_4200, plaintext_s0[103]}), .a ({new_AGEMA_signal_4111, new_AGEMA_signal_4110, stateArray_outS10ser_MC[7]}), .c ({new_AGEMA_signal_4203, new_AGEMA_signal_4202, stateArray_inS03ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS10ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2481, new_AGEMA_signal_2480, plaintext_s0[88]}), .a ({new_AGEMA_signal_2483, ciphertext_s1[80], ciphertext_s0[80]}), .c ({new_AGEMA_signal_2485, new_AGEMA_signal_2484, stateArray_inS10ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS10ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2487, new_AGEMA_signal_2486, plaintext_s0[89]}), .a ({new_AGEMA_signal_2489, ciphertext_s1[81], ciphertext_s0[81]}), .c ({new_AGEMA_signal_2491, new_AGEMA_signal_2490, stateArray_inS10ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS10ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2493, new_AGEMA_signal_2492, plaintext_s0[90]}), .a ({new_AGEMA_signal_2495, ciphertext_s1[82], ciphertext_s0[82]}), .c ({new_AGEMA_signal_2497, new_AGEMA_signal_2496, stateArray_inS10ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS10ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2499, new_AGEMA_signal_2498, plaintext_s0[91]}), .a ({new_AGEMA_signal_2501, ciphertext_s1[83], ciphertext_s0[83]}), .c ({new_AGEMA_signal_2503, new_AGEMA_signal_2502, stateArray_inS10ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS10ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2505, new_AGEMA_signal_2504, plaintext_s0[92]}), .a ({new_AGEMA_signal_2507, ciphertext_s1[84], ciphertext_s0[84]}), .c ({new_AGEMA_signal_2509, new_AGEMA_signal_2508, stateArray_inS10ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS10ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2511, new_AGEMA_signal_2510, plaintext_s0[93]}), .a ({new_AGEMA_signal_2513, ciphertext_s1[85], ciphertext_s0[85]}), .c ({new_AGEMA_signal_2515, new_AGEMA_signal_2514, stateArray_inS10ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS10ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2517, new_AGEMA_signal_2516, plaintext_s0[94]}), .a ({new_AGEMA_signal_2519, ciphertext_s1[86], ciphertext_s0[86]}), .c ({new_AGEMA_signal_2521, new_AGEMA_signal_2520, stateArray_inS10ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS10ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2523, new_AGEMA_signal_2522, plaintext_s0[95]}), .a ({new_AGEMA_signal_2525, ciphertext_s1[87], ciphertext_s0[87]}), .c ({new_AGEMA_signal_2527, new_AGEMA_signal_2526, stateArray_inS10ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS11ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2529, new_AGEMA_signal_2528, plaintext_s0[80]}), .a ({new_AGEMA_signal_2531, ciphertext_s1[72], ciphertext_s0[72]}), .c ({new_AGEMA_signal_2533, new_AGEMA_signal_2532, stateArray_inS11ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS11ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2535, new_AGEMA_signal_2534, plaintext_s0[81]}), .a ({new_AGEMA_signal_2537, ciphertext_s1[73], ciphertext_s0[73]}), .c ({new_AGEMA_signal_2539, new_AGEMA_signal_2538, stateArray_inS11ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS11ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2541, new_AGEMA_signal_2540, plaintext_s0[82]}), .a ({new_AGEMA_signal_2543, ciphertext_s1[74], ciphertext_s0[74]}), .c ({new_AGEMA_signal_2545, new_AGEMA_signal_2544, stateArray_inS11ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS11ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2547, new_AGEMA_signal_2546, plaintext_s0[83]}), .a ({new_AGEMA_signal_2549, ciphertext_s1[75], ciphertext_s0[75]}), .c ({new_AGEMA_signal_2551, new_AGEMA_signal_2550, stateArray_inS11ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS11ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2553, new_AGEMA_signal_2552, plaintext_s0[84]}), .a ({new_AGEMA_signal_2555, ciphertext_s1[76], ciphertext_s0[76]}), .c ({new_AGEMA_signal_2557, new_AGEMA_signal_2556, stateArray_inS11ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS11ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2559, new_AGEMA_signal_2558, plaintext_s0[85]}), .a ({new_AGEMA_signal_2561, ciphertext_s1[77], ciphertext_s0[77]}), .c ({new_AGEMA_signal_2563, new_AGEMA_signal_2562, stateArray_inS11ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS11ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2565, new_AGEMA_signal_2564, plaintext_s0[86]}), .a ({new_AGEMA_signal_2567, ciphertext_s1[78], ciphertext_s0[78]}), .c ({new_AGEMA_signal_2569, new_AGEMA_signal_2568, stateArray_inS11ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS11ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2479, new_AGEMA_signal_2478, stateArray_n30}), .b ({new_AGEMA_signal_2571, new_AGEMA_signal_2570, plaintext_s0[87]}), .a ({new_AGEMA_signal_2573, ciphertext_s1[79], ciphertext_s0[79]}), .c ({new_AGEMA_signal_2575, new_AGEMA_signal_2574, stateArray_inS11ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS12ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_2579, new_AGEMA_signal_2578, plaintext_s0[72]}), .a ({new_AGEMA_signal_2581, ciphertext_s1[64], ciphertext_s0[64]}), .c ({new_AGEMA_signal_2583, new_AGEMA_signal_2582, stateArray_inS12ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS12ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_2585, new_AGEMA_signal_2584, plaintext_s0[73]}), .a ({new_AGEMA_signal_2587, ciphertext_s1[65], ciphertext_s0[65]}), .c ({new_AGEMA_signal_2589, new_AGEMA_signal_2588, stateArray_inS12ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS12ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_2591, new_AGEMA_signal_2590, plaintext_s0[74]}), .a ({new_AGEMA_signal_2593, ciphertext_s1[66], ciphertext_s0[66]}), .c ({new_AGEMA_signal_2595, new_AGEMA_signal_2594, stateArray_inS12ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS12ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_2597, new_AGEMA_signal_2596, plaintext_s0[75]}), .a ({new_AGEMA_signal_2599, ciphertext_s1[67], ciphertext_s0[67]}), .c ({new_AGEMA_signal_2601, new_AGEMA_signal_2600, stateArray_inS12ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS12ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_2603, new_AGEMA_signal_2602, plaintext_s0[76]}), .a ({new_AGEMA_signal_2605, ciphertext_s1[68], ciphertext_s0[68]}), .c ({new_AGEMA_signal_2607, new_AGEMA_signal_2606, stateArray_inS12ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS12ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_2609, new_AGEMA_signal_2608, plaintext_s0[77]}), .a ({new_AGEMA_signal_2611, ciphertext_s1[69], ciphertext_s0[69]}), .c ({new_AGEMA_signal_2613, new_AGEMA_signal_2612, stateArray_inS12ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS12ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_2615, new_AGEMA_signal_2614, plaintext_s0[78]}), .a ({new_AGEMA_signal_2617, ciphertext_s1[70], ciphertext_s0[70]}), .c ({new_AGEMA_signal_2619, new_AGEMA_signal_2618, stateArray_inS12ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS12ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_2621, new_AGEMA_signal_2620, plaintext_s0[79]}), .a ({new_AGEMA_signal_2623, ciphertext_s1[71], ciphertext_s0[71]}), .c ({new_AGEMA_signal_2625, new_AGEMA_signal_2624, stateArray_inS12ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS20_MC_mux_inst_0_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}), .a ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, StateInMC[16]}), .c ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, stateArray_outS20ser_MC[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS20_MC_mux_inst_1_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}), .a ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, StateInMC[17]}), .c ({new_AGEMA_signal_4115, new_AGEMA_signal_4114, stateArray_outS20ser_MC[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS20_MC_mux_inst_2_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}), .a ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, StateInMC[18]}), .c ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, stateArray_outS20ser_MC[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS20_MC_mux_inst_3_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}), .a ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, StateInMC[19]}), .c ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, stateArray_outS20ser_MC[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS20_MC_mux_inst_4_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}), .a ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, StateInMC[20]}), .c ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, stateArray_outS20ser_MC[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS20_MC_mux_inst_5_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}), .a ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, StateInMC[21]}), .c ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, stateArray_outS20ser_MC[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS20_MC_mux_inst_6_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}), .a ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, StateInMC[22]}), .c ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, stateArray_outS20ser_MC[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS20_MC_mux_inst_7_U1 ( .s ({new_AGEMA_signal_4095, new_AGEMA_signal_4094, stateArray_n23}), .b ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .a ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, StateInMC[23]}), .c ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, stateArray_outS20ser_MC[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS13ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_4205, new_AGEMA_signal_4204, plaintext_s0[64]}), .a ({new_AGEMA_signal_4113, new_AGEMA_signal_4112, stateArray_outS20ser_MC[0]}), .c ({new_AGEMA_signal_4207, new_AGEMA_signal_4206, stateArray_inS13ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS13ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_4209, new_AGEMA_signal_4208, plaintext_s0[65]}), .a ({new_AGEMA_signal_4115, new_AGEMA_signal_4114, stateArray_outS20ser_MC[1]}), .c ({new_AGEMA_signal_4211, new_AGEMA_signal_4210, stateArray_inS13ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS13ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_4213, new_AGEMA_signal_4212, plaintext_s0[66]}), .a ({new_AGEMA_signal_4117, new_AGEMA_signal_4116, stateArray_outS20ser_MC[2]}), .c ({new_AGEMA_signal_4215, new_AGEMA_signal_4214, stateArray_inS13ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS13ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_4217, new_AGEMA_signal_4216, plaintext_s0[67]}), .a ({new_AGEMA_signal_4119, new_AGEMA_signal_4118, stateArray_outS20ser_MC[3]}), .c ({new_AGEMA_signal_4219, new_AGEMA_signal_4218, stateArray_inS13ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS13ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_4221, new_AGEMA_signal_4220, plaintext_s0[68]}), .a ({new_AGEMA_signal_4121, new_AGEMA_signal_4120, stateArray_outS20ser_MC[4]}), .c ({new_AGEMA_signal_4223, new_AGEMA_signal_4222, stateArray_inS13ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS13ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_4225, new_AGEMA_signal_4224, plaintext_s0[69]}), .a ({new_AGEMA_signal_4123, new_AGEMA_signal_4122, stateArray_outS20ser_MC[5]}), .c ({new_AGEMA_signal_4227, new_AGEMA_signal_4226, stateArray_inS13ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS13ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_4229, new_AGEMA_signal_4228, plaintext_s0[70]}), .a ({new_AGEMA_signal_4125, new_AGEMA_signal_4124, stateArray_outS20ser_MC[6]}), .c ({new_AGEMA_signal_4231, new_AGEMA_signal_4230, stateArray_inS13ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS13ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2577, new_AGEMA_signal_2576, stateArray_n29}), .b ({new_AGEMA_signal_4233, new_AGEMA_signal_4232, plaintext_s0[71]}), .a ({new_AGEMA_signal_4127, new_AGEMA_signal_4126, stateArray_outS20ser_MC[7]}), .c ({new_AGEMA_signal_4235, new_AGEMA_signal_4234, stateArray_inS13ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS20ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2629, new_AGEMA_signal_2628, plaintext_s0[56]}), .a ({new_AGEMA_signal_2631, ciphertext_s1[48], ciphertext_s0[48]}), .c ({new_AGEMA_signal_2633, new_AGEMA_signal_2632, stateArray_inS20ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS20ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2635, new_AGEMA_signal_2634, plaintext_s0[57]}), .a ({new_AGEMA_signal_2637, ciphertext_s1[49], ciphertext_s0[49]}), .c ({new_AGEMA_signal_2639, new_AGEMA_signal_2638, stateArray_inS20ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS20ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2641, new_AGEMA_signal_2640, plaintext_s0[58]}), .a ({new_AGEMA_signal_2643, ciphertext_s1[50], ciphertext_s0[50]}), .c ({new_AGEMA_signal_2645, new_AGEMA_signal_2644, stateArray_inS20ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS20ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2647, new_AGEMA_signal_2646, plaintext_s0[59]}), .a ({new_AGEMA_signal_2649, ciphertext_s1[51], ciphertext_s0[51]}), .c ({new_AGEMA_signal_2651, new_AGEMA_signal_2650, stateArray_inS20ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS20ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2653, new_AGEMA_signal_2652, plaintext_s0[60]}), .a ({new_AGEMA_signal_2655, ciphertext_s1[52], ciphertext_s0[52]}), .c ({new_AGEMA_signal_2657, new_AGEMA_signal_2656, stateArray_inS20ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS20ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2659, new_AGEMA_signal_2658, plaintext_s0[61]}), .a ({new_AGEMA_signal_2661, ciphertext_s1[53], ciphertext_s0[53]}), .c ({new_AGEMA_signal_2663, new_AGEMA_signal_2662, stateArray_inS20ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS20ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2665, new_AGEMA_signal_2664, plaintext_s0[62]}), .a ({new_AGEMA_signal_2667, ciphertext_s1[54], ciphertext_s0[54]}), .c ({new_AGEMA_signal_2669, new_AGEMA_signal_2668, stateArray_inS20ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS20ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2671, new_AGEMA_signal_2670, plaintext_s0[63]}), .a ({new_AGEMA_signal_2673, ciphertext_s1[55], ciphertext_s0[55]}), .c ({new_AGEMA_signal_2675, new_AGEMA_signal_2674, stateArray_inS20ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS21ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2677, new_AGEMA_signal_2676, plaintext_s0[48]}), .a ({new_AGEMA_signal_2679, ciphertext_s1[40], ciphertext_s0[40]}), .c ({new_AGEMA_signal_2681, new_AGEMA_signal_2680, stateArray_inS21ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS21ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2683, new_AGEMA_signal_2682, plaintext_s0[49]}), .a ({new_AGEMA_signal_2685, ciphertext_s1[41], ciphertext_s0[41]}), .c ({new_AGEMA_signal_2687, new_AGEMA_signal_2686, stateArray_inS21ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS21ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2689, new_AGEMA_signal_2688, plaintext_s0[50]}), .a ({new_AGEMA_signal_2691, ciphertext_s1[42], ciphertext_s0[42]}), .c ({new_AGEMA_signal_2693, new_AGEMA_signal_2692, stateArray_inS21ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS21ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2695, new_AGEMA_signal_2694, plaintext_s0[51]}), .a ({new_AGEMA_signal_2697, ciphertext_s1[43], ciphertext_s0[43]}), .c ({new_AGEMA_signal_2699, new_AGEMA_signal_2698, stateArray_inS21ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS21ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2701, new_AGEMA_signal_2700, plaintext_s0[52]}), .a ({new_AGEMA_signal_2703, ciphertext_s1[44], ciphertext_s0[44]}), .c ({new_AGEMA_signal_2705, new_AGEMA_signal_2704, stateArray_inS21ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS21ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2707, new_AGEMA_signal_2706, plaintext_s0[53]}), .a ({new_AGEMA_signal_2709, ciphertext_s1[45], ciphertext_s0[45]}), .c ({new_AGEMA_signal_2711, new_AGEMA_signal_2710, stateArray_inS21ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS21ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2713, new_AGEMA_signal_2712, plaintext_s0[54]}), .a ({new_AGEMA_signal_2715, ciphertext_s1[46], ciphertext_s0[46]}), .c ({new_AGEMA_signal_2717, new_AGEMA_signal_2716, stateArray_inS21ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS21ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2627, new_AGEMA_signal_2626, stateArray_n28}), .b ({new_AGEMA_signal_2719, new_AGEMA_signal_2718, plaintext_s0[55]}), .a ({new_AGEMA_signal_2721, ciphertext_s1[47], ciphertext_s0[47]}), .c ({new_AGEMA_signal_2723, new_AGEMA_signal_2722, stateArray_inS21ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS22ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_2727, new_AGEMA_signal_2726, plaintext_s0[40]}), .a ({new_AGEMA_signal_2729, ciphertext_s1[32], ciphertext_s0[32]}), .c ({new_AGEMA_signal_2731, new_AGEMA_signal_2730, stateArray_inS22ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS22ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_2733, new_AGEMA_signal_2732, plaintext_s0[41]}), .a ({new_AGEMA_signal_2735, ciphertext_s1[33], ciphertext_s0[33]}), .c ({new_AGEMA_signal_2737, new_AGEMA_signal_2736, stateArray_inS22ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS22ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_2739, new_AGEMA_signal_2738, plaintext_s0[42]}), .a ({new_AGEMA_signal_2741, ciphertext_s1[34], ciphertext_s0[34]}), .c ({new_AGEMA_signal_2743, new_AGEMA_signal_2742, stateArray_inS22ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS22ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_2745, new_AGEMA_signal_2744, plaintext_s0[43]}), .a ({new_AGEMA_signal_2747, ciphertext_s1[35], ciphertext_s0[35]}), .c ({new_AGEMA_signal_2749, new_AGEMA_signal_2748, stateArray_inS22ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS22ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_2751, new_AGEMA_signal_2750, plaintext_s0[44]}), .a ({new_AGEMA_signal_2753, ciphertext_s1[36], ciphertext_s0[36]}), .c ({new_AGEMA_signal_2755, new_AGEMA_signal_2754, stateArray_inS22ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS22ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_2757, new_AGEMA_signal_2756, plaintext_s0[45]}), .a ({new_AGEMA_signal_2759, ciphertext_s1[37], ciphertext_s0[37]}), .c ({new_AGEMA_signal_2761, new_AGEMA_signal_2760, stateArray_inS22ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS22ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_2763, new_AGEMA_signal_2762, plaintext_s0[46]}), .a ({new_AGEMA_signal_2765, ciphertext_s1[38], ciphertext_s0[38]}), .c ({new_AGEMA_signal_2767, new_AGEMA_signal_2766, stateArray_inS22ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS22ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_2769, new_AGEMA_signal_2768, plaintext_s0[47]}), .a ({new_AGEMA_signal_2771, ciphertext_s1[39], ciphertext_s0[39]}), .c ({new_AGEMA_signal_2773, new_AGEMA_signal_2772, stateArray_inS22ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS30_MC_mux_inst_0_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}), .a ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, StateInMC[8]}), .c ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, stateArray_outS30ser_MC[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS30_MC_mux_inst_1_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}), .a ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, StateInMC[9]}), .c ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, stateArray_outS30ser_MC[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS30_MC_mux_inst_2_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}), .a ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, StateInMC[10]}), .c ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, stateArray_outS30ser_MC[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS30_MC_mux_inst_3_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}), .a ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, StateInMC[11]}), .c ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, stateArray_outS30ser_MC[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS30_MC_mux_inst_4_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}), .a ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, StateInMC[12]}), .c ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, stateArray_outS30ser_MC[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS30_MC_mux_inst_5_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}), .a ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, StateInMC[13]}), .c ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, stateArray_outS30ser_MC[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS30_MC_mux_inst_6_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}), .a ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, StateInMC[14]}), .c ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, stateArray_outS30ser_MC[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_outS30_MC_mux_inst_7_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .a ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, StateInMC[15]}), .c ({new_AGEMA_signal_4145, new_AGEMA_signal_4144, stateArray_outS30ser_MC[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS23ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_4237, new_AGEMA_signal_4236, plaintext_s0[32]}), .a ({new_AGEMA_signal_4131, new_AGEMA_signal_4130, stateArray_outS30ser_MC[0]}), .c ({new_AGEMA_signal_4239, new_AGEMA_signal_4238, stateArray_inS23ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS23ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_4241, new_AGEMA_signal_4240, plaintext_s0[33]}), .a ({new_AGEMA_signal_4133, new_AGEMA_signal_4132, stateArray_outS30ser_MC[1]}), .c ({new_AGEMA_signal_4243, new_AGEMA_signal_4242, stateArray_inS23ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS23ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_4245, new_AGEMA_signal_4244, plaintext_s0[34]}), .a ({new_AGEMA_signal_4135, new_AGEMA_signal_4134, stateArray_outS30ser_MC[2]}), .c ({new_AGEMA_signal_4247, new_AGEMA_signal_4246, stateArray_inS23ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS23ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_4249, new_AGEMA_signal_4248, plaintext_s0[35]}), .a ({new_AGEMA_signal_4137, new_AGEMA_signal_4136, stateArray_outS30ser_MC[3]}), .c ({new_AGEMA_signal_4251, new_AGEMA_signal_4250, stateArray_inS23ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS23ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_4253, new_AGEMA_signal_4252, plaintext_s0[36]}), .a ({new_AGEMA_signal_4139, new_AGEMA_signal_4138, stateArray_outS30ser_MC[4]}), .c ({new_AGEMA_signal_4255, new_AGEMA_signal_4254, stateArray_inS23ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS23ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_4257, new_AGEMA_signal_4256, plaintext_s0[37]}), .a ({new_AGEMA_signal_4141, new_AGEMA_signal_4140, stateArray_outS30ser_MC[5]}), .c ({new_AGEMA_signal_4259, new_AGEMA_signal_4258, stateArray_inS23ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS23ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_4261, new_AGEMA_signal_4260, plaintext_s0[38]}), .a ({new_AGEMA_signal_4143, new_AGEMA_signal_4142, stateArray_outS30ser_MC[6]}), .c ({new_AGEMA_signal_4263, new_AGEMA_signal_4262, stateArray_inS23ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS23ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2725, new_AGEMA_signal_2724, stateArray_n27}), .b ({new_AGEMA_signal_4265, new_AGEMA_signal_4264, plaintext_s0[39]}), .a ({new_AGEMA_signal_4145, new_AGEMA_signal_4144, stateArray_outS30ser_MC[7]}), .c ({new_AGEMA_signal_4267, new_AGEMA_signal_4266, stateArray_inS23ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS30ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2777, new_AGEMA_signal_2776, plaintext_s0[24]}), .a ({new_AGEMA_signal_2779, ciphertext_s1[16], ciphertext_s0[16]}), .c ({new_AGEMA_signal_2781, new_AGEMA_signal_2780, stateArray_inS30ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS30ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2783, new_AGEMA_signal_2782, plaintext_s0[25]}), .a ({new_AGEMA_signal_2785, ciphertext_s1[17], ciphertext_s0[17]}), .c ({new_AGEMA_signal_2787, new_AGEMA_signal_2786, stateArray_inS30ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS30ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2789, new_AGEMA_signal_2788, plaintext_s0[26]}), .a ({new_AGEMA_signal_2791, ciphertext_s1[18], ciphertext_s0[18]}), .c ({new_AGEMA_signal_2793, new_AGEMA_signal_2792, stateArray_inS30ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS30ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2795, new_AGEMA_signal_2794, plaintext_s0[27]}), .a ({new_AGEMA_signal_2797, ciphertext_s1[19], ciphertext_s0[19]}), .c ({new_AGEMA_signal_2799, new_AGEMA_signal_2798, stateArray_inS30ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS30ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2801, new_AGEMA_signal_2800, plaintext_s0[28]}), .a ({new_AGEMA_signal_2803, ciphertext_s1[20], ciphertext_s0[20]}), .c ({new_AGEMA_signal_2805, new_AGEMA_signal_2804, stateArray_inS30ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS30ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2807, new_AGEMA_signal_2806, plaintext_s0[29]}), .a ({new_AGEMA_signal_2809, ciphertext_s1[21], ciphertext_s0[21]}), .c ({new_AGEMA_signal_2811, new_AGEMA_signal_2810, stateArray_inS30ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS30ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2813, new_AGEMA_signal_2812, plaintext_s0[30]}), .a ({new_AGEMA_signal_2815, ciphertext_s1[22], ciphertext_s0[22]}), .c ({new_AGEMA_signal_2817, new_AGEMA_signal_2816, stateArray_inS30ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS30ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2819, new_AGEMA_signal_2818, plaintext_s0[31]}), .a ({new_AGEMA_signal_2821, ciphertext_s1[23], ciphertext_s0[23]}), .c ({new_AGEMA_signal_2823, new_AGEMA_signal_2822, stateArray_inS30ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS31ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2825, new_AGEMA_signal_2824, plaintext_s0[16]}), .a ({new_AGEMA_signal_2827, ciphertext_s1[8], ciphertext_s0[8]}), .c ({new_AGEMA_signal_2829, new_AGEMA_signal_2828, stateArray_inS31ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS31ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2831, new_AGEMA_signal_2830, plaintext_s0[17]}), .a ({new_AGEMA_signal_2833, ciphertext_s1[9], ciphertext_s0[9]}), .c ({new_AGEMA_signal_2835, new_AGEMA_signal_2834, stateArray_inS31ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS31ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2837, new_AGEMA_signal_2836, plaintext_s0[18]}), .a ({new_AGEMA_signal_2839, ciphertext_s1[10], ciphertext_s0[10]}), .c ({new_AGEMA_signal_2841, new_AGEMA_signal_2840, stateArray_inS31ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS31ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2843, new_AGEMA_signal_2842, plaintext_s0[19]}), .a ({new_AGEMA_signal_2845, ciphertext_s1[11], ciphertext_s0[11]}), .c ({new_AGEMA_signal_2847, new_AGEMA_signal_2846, stateArray_inS31ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS31ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2849, new_AGEMA_signal_2848, plaintext_s0[20]}), .a ({new_AGEMA_signal_2851, ciphertext_s1[12], ciphertext_s0[12]}), .c ({new_AGEMA_signal_2853, new_AGEMA_signal_2852, stateArray_inS31ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS31ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2855, new_AGEMA_signal_2854, plaintext_s0[21]}), .a ({new_AGEMA_signal_2857, ciphertext_s1[13], ciphertext_s0[13]}), .c ({new_AGEMA_signal_2859, new_AGEMA_signal_2858, stateArray_inS31ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS31ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2861, new_AGEMA_signal_2860, plaintext_s0[22]}), .a ({new_AGEMA_signal_2863, ciphertext_s1[14], ciphertext_s0[14]}), .c ({new_AGEMA_signal_2865, new_AGEMA_signal_2864, stateArray_inS31ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS31ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2775, new_AGEMA_signal_2774, stateArray_n26}), .b ({new_AGEMA_signal_2867, new_AGEMA_signal_2866, plaintext_s0[23]}), .a ({new_AGEMA_signal_2869, ciphertext_s1[15], ciphertext_s0[15]}), .c ({new_AGEMA_signal_2871, new_AGEMA_signal_2870, stateArray_inS31ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS32ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_2875, new_AGEMA_signal_2874, plaintext_s0[8]}), .a ({new_AGEMA_signal_2877, ciphertext_s1[0], ciphertext_s0[0]}), .c ({new_AGEMA_signal_2879, new_AGEMA_signal_2878, stateArray_inS32ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS32ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_2881, new_AGEMA_signal_2880, plaintext_s0[9]}), .a ({new_AGEMA_signal_2883, ciphertext_s1[1], ciphertext_s0[1]}), .c ({new_AGEMA_signal_2885, new_AGEMA_signal_2884, stateArray_inS32ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS32ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_2887, new_AGEMA_signal_2886, plaintext_s0[10]}), .a ({new_AGEMA_signal_2889, ciphertext_s1[2], ciphertext_s0[2]}), .c ({new_AGEMA_signal_2891, new_AGEMA_signal_2890, stateArray_inS32ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS32ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_2893, new_AGEMA_signal_2892, plaintext_s0[11]}), .a ({new_AGEMA_signal_2895, ciphertext_s1[3], ciphertext_s0[3]}), .c ({new_AGEMA_signal_2897, new_AGEMA_signal_2896, stateArray_inS32ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS32ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_2899, new_AGEMA_signal_2898, plaintext_s0[12]}), .a ({new_AGEMA_signal_2901, ciphertext_s1[4], ciphertext_s0[4]}), .c ({new_AGEMA_signal_2903, new_AGEMA_signal_2902, stateArray_inS32ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS32ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_2905, new_AGEMA_signal_2904, plaintext_s0[13]}), .a ({new_AGEMA_signal_2907, ciphertext_s1[5], ciphertext_s0[5]}), .c ({new_AGEMA_signal_2909, new_AGEMA_signal_2908, stateArray_inS32ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS32ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_2911, new_AGEMA_signal_2910, plaintext_s0[14]}), .a ({new_AGEMA_signal_2913, ciphertext_s1[6], ciphertext_s0[6]}), .c ({new_AGEMA_signal_2915, new_AGEMA_signal_2914, stateArray_inS32ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS32ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_2917, new_AGEMA_signal_2916, plaintext_s0[15]}), .a ({new_AGEMA_signal_2919, ciphertext_s1[7], ciphertext_s0[7]}), .c ({new_AGEMA_signal_2921, new_AGEMA_signal_2920, stateArray_inS32ser[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_input_MC_mux_inst_0_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_5027, new_AGEMA_signal_5026, StateIn[0]}), .a ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, StateInMC[0]}), .c ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, stateArray_input_MC[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_input_MC_mux_inst_1_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_5045, new_AGEMA_signal_5044, StateIn[1]}), .a ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, StateInMC[1]}), .c ({new_AGEMA_signal_5077, new_AGEMA_signal_5076, stateArray_input_MC[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_input_MC_mux_inst_2_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_5047, new_AGEMA_signal_5046, StateIn[2]}), .a ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, StateInMC[2]}), .c ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, stateArray_input_MC[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_input_MC_mux_inst_3_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_5049, new_AGEMA_signal_5048, StateIn[3]}), .a ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, StateInMC[3]}), .c ({new_AGEMA_signal_5081, new_AGEMA_signal_5080, stateArray_input_MC[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_input_MC_mux_inst_4_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_5051, new_AGEMA_signal_5050, StateIn[4]}), .a ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, StateInMC[4]}), .c ({new_AGEMA_signal_5083, new_AGEMA_signal_5082, stateArray_input_MC[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_input_MC_mux_inst_5_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_5053, new_AGEMA_signal_5052, StateIn[5]}), .a ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, StateInMC[5]}), .c ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, stateArray_input_MC[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_input_MC_mux_inst_6_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_5055, new_AGEMA_signal_5054, StateIn[6]}), .a ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, StateInMC[6]}), .c ({new_AGEMA_signal_5087, new_AGEMA_signal_5086, stateArray_input_MC[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_input_MC_mux_inst_7_U1 ( .s ({new_AGEMA_signal_4129, new_AGEMA_signal_4128, stateArray_n22}), .b ({new_AGEMA_signal_5057, new_AGEMA_signal_5056, StateIn[7]}), .a ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, StateInMC[7]}), .c ({new_AGEMA_signal_5089, new_AGEMA_signal_5088, stateArray_input_MC[7]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS33ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_5091, new_AGEMA_signal_5090, plaintext_s0[0]}), .a ({new_AGEMA_signal_5059, new_AGEMA_signal_5058, stateArray_input_MC[0]}), .c ({new_AGEMA_signal_5093, new_AGEMA_signal_5092, stateArray_inS33ser[0]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS33ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_5113, new_AGEMA_signal_5112, plaintext_s0[1]}), .a ({new_AGEMA_signal_5077, new_AGEMA_signal_5076, stateArray_input_MC[1]}), .c ({new_AGEMA_signal_5115, new_AGEMA_signal_5114, stateArray_inS33ser[1]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS33ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_5117, new_AGEMA_signal_5116, plaintext_s0[2]}), .a ({new_AGEMA_signal_5079, new_AGEMA_signal_5078, stateArray_input_MC[2]}), .c ({new_AGEMA_signal_5119, new_AGEMA_signal_5118, stateArray_inS33ser[2]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS33ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_5121, new_AGEMA_signal_5120, plaintext_s0[3]}), .a ({new_AGEMA_signal_5081, new_AGEMA_signal_5080, stateArray_input_MC[3]}), .c ({new_AGEMA_signal_5123, new_AGEMA_signal_5122, stateArray_inS33ser[3]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS33ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_5125, new_AGEMA_signal_5124, plaintext_s0[4]}), .a ({new_AGEMA_signal_5083, new_AGEMA_signal_5082, stateArray_input_MC[4]}), .c ({new_AGEMA_signal_5127, new_AGEMA_signal_5126, stateArray_inS33ser[4]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS33ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_5129, new_AGEMA_signal_5128, plaintext_s0[5]}), .a ({new_AGEMA_signal_5085, new_AGEMA_signal_5084, stateArray_input_MC[5]}), .c ({new_AGEMA_signal_5131, new_AGEMA_signal_5130, stateArray_inS33ser[5]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS33ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_5133, new_AGEMA_signal_5132, plaintext_s0[6]}), .a ({new_AGEMA_signal_5087, new_AGEMA_signal_5086, stateArray_input_MC[6]}), .c ({new_AGEMA_signal_5135, new_AGEMA_signal_5134, stateArray_inS33ser[6]}) ) ;
    mux2_masked_LMDPL stateArray_MUX_inS33ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2873, new_AGEMA_signal_2872, stateArray_n25}), .b ({new_AGEMA_signal_5137, new_AGEMA_signal_5136, plaintext_s0[7]}), .a ({new_AGEMA_signal_5089, new_AGEMA_signal_5088, stateArray_input_MC[7]}), .c ({new_AGEMA_signal_5139, new_AGEMA_signal_5138, stateArray_inS33ser[7]}) ) ;
    INV_X1 MUX_StateInMC_U3 ( .A (intFinal), .ZN (MUX_StateInMC_n7) ) ;
    INV_X1 MUX_StateInMC_U2 ( .A (MUX_StateInMC_n7), .ZN (MUX_StateInMC_n6) ) ;
    INV_X1 MUX_StateInMC_U1 ( .A (MUX_StateInMC_n7), .ZN (MUX_StateInMC_n5) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, MCout[0]}), .a ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_3781, new_AGEMA_signal_3780, StateInMC[0]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, MCout[1]}), .a ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_3785, new_AGEMA_signal_3784, StateInMC[1]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, MCout[2]}), .a ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_3727, new_AGEMA_signal_3726, StateInMC[2]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, MCout[3]}), .a ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_3787, new_AGEMA_signal_3786, StateInMC[3]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, MCout[4]}), .a ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_3789, new_AGEMA_signal_3788, StateInMC[4]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, MCout[5]}), .a ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_3729, new_AGEMA_signal_3728, StateInMC[5]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, MCout[6]}), .a ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_3731, new_AGEMA_signal_3730, StateInMC[6]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3725, new_AGEMA_signal_3724, intFinal}), .b ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, MCout[7]}), .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_3733, new_AGEMA_signal_3732, StateInMC[7]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_8_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, MCout[8]}), .a ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_3791, new_AGEMA_signal_3790, StateInMC[8]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_9_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, MCout[9]}), .a ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_3793, new_AGEMA_signal_3792, StateInMC[9]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_10_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, MCout[10]}), .a ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_3795, new_AGEMA_signal_3794, StateInMC[10]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_11_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, MCout[11]}), .a ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_3797, new_AGEMA_signal_3796, StateInMC[11]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_12_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, MCout[12]}), .a ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_3799, new_AGEMA_signal_3798, StateInMC[12]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_13_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, MCout[13]}), .a ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_3801, new_AGEMA_signal_3800, StateInMC[13]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_14_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, MCout[14]}), .a ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_3803, new_AGEMA_signal_3802, StateInMC[14]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_15_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, MCout[15]}), .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_3805, new_AGEMA_signal_3804, StateInMC[15]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_16_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, MCout[16]}), .a ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_3807, new_AGEMA_signal_3806, StateInMC[16]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_17_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, MCout[17]}), .a ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_3809, new_AGEMA_signal_3808, StateInMC[17]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_18_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, MCout[18]}), .a ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_3811, new_AGEMA_signal_3810, StateInMC[18]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_19_U1 ( .s ({new_AGEMA_signal_3783, new_AGEMA_signal_3782, MUX_StateInMC_n6}), .b ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, MCout[19]}), .a ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_3813, new_AGEMA_signal_3812, StateInMC[19]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_20_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, MCout[20]}), .a ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_3815, new_AGEMA_signal_3814, StateInMC[20]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_21_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, MCout[21]}), .a ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_3817, new_AGEMA_signal_3816, StateInMC[21]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_22_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, MCout[22]}), .a ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_3819, new_AGEMA_signal_3818, StateInMC[22]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_23_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, MCout[23]}), .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_3821, new_AGEMA_signal_3820, StateInMC[23]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_24_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, MCout[24]}), .a ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_3823, new_AGEMA_signal_3822, StateInMC[24]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_25_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3739, new_AGEMA_signal_3738, MCout[25]}), .a ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_3825, new_AGEMA_signal_3824, StateInMC[25]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_26_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, MCout[26]}), .a ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_3827, new_AGEMA_signal_3826, StateInMC[26]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_27_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, MCout[27]}), .a ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_3829, new_AGEMA_signal_3828, StateInMC[27]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_28_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, MCout[28]}), .a ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_3831, new_AGEMA_signal_3830, StateInMC[28]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_29_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, MCout[29]}), .a ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_3833, new_AGEMA_signal_3832, StateInMC[29]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_30_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, MCout[30]}), .a ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_3835, new_AGEMA_signal_3834, StateInMC[30]}) ) ;
    mux2_masked_LMDPL MUX_StateInMC_mux_inst_31_U1 ( .s ({new_AGEMA_signal_3779, new_AGEMA_signal_3778, MUX_StateInMC_n5}), .b ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, MCout[31]}), .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_3837, new_AGEMA_signal_3836, StateInMC[31]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) KeyArray_U50 ( .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, KeyArray_outS01ser_7_}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[7]}), .c ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, KeyArray_outS01ser_XOR_00[7]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) KeyArray_U49 ( .a ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, KeyArray_outS01ser_6_}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, keyStateIn[6]}), .c ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, KeyArray_outS01ser_XOR_00[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) KeyArray_U48 ( .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, KeyArray_outS01ser_5_}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, keyStateIn[5]}), .c ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, KeyArray_outS01ser_XOR_00[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) KeyArray_U47 ( .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, KeyArray_outS01ser_4_}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[4]}), .c ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, KeyArray_outS01ser_XOR_00[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) KeyArray_U46 ( .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, KeyArray_outS01ser_3_}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, keyStateIn[3]}), .c ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, KeyArray_outS01ser_XOR_00[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) KeyArray_U45 ( .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_2_}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, keyStateIn[2]}), .c ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, KeyArray_outS01ser_XOR_00[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) KeyArray_U44 ( .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, KeyArray_outS01ser_1_}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .c ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, KeyArray_outS01ser_XOR_00[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) KeyArray_U43 ( .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, KeyArray_outS01ser_0_}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, keyStateIn[0]}), .c ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, KeyArray_outS01ser_XOR_00[0]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U42 ( .a ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, KeyArray_n55}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[7]}), .c ({new_AGEMA_signal_5095, new_AGEMA_signal_5094, KeyArray_inS30par[7]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U41 ( .a ({LMDPL_pre1, 1'b0, roundConstant[7]}), .b ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, SboxOut[7]}), .c ({new_AGEMA_signal_5061, new_AGEMA_signal_5060, KeyArray_n55}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U40 ( .a ({new_AGEMA_signal_5063, new_AGEMA_signal_5062, KeyArray_n54}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, keyStateIn[6]}), .c ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, KeyArray_inS30par[6]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U39 ( .a ({LMDPL_pre1, 1'b0, roundConstant[6]}), .b ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, SboxOut[6]}), .c ({new_AGEMA_signal_5063, new_AGEMA_signal_5062, KeyArray_n54}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U38 ( .a ({new_AGEMA_signal_5065, new_AGEMA_signal_5064, KeyArray_n53}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, keyStateIn[5]}), .c ({new_AGEMA_signal_5099, new_AGEMA_signal_5098, KeyArray_inS30par[5]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U37 ( .a ({LMDPL_pre1, 1'b0, roundConstant[5]}), .b ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, SboxOut[5]}), .c ({new_AGEMA_signal_5065, new_AGEMA_signal_5064, KeyArray_n53}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U36 ( .a ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, KeyArray_n52}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[4]}), .c ({new_AGEMA_signal_5101, new_AGEMA_signal_5100, KeyArray_inS30par[4]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U35 ( .a ({LMDPL_pre1, 1'b0, roundConstant[4]}), .b ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, SboxOut[4]}), .c ({new_AGEMA_signal_5067, new_AGEMA_signal_5066, KeyArray_n52}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U34 ( .a ({new_AGEMA_signal_5069, new_AGEMA_signal_5068, KeyArray_n51}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, keyStateIn[3]}), .c ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, KeyArray_inS30par[3]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U33 ( .a ({LMDPL_pre1, 1'b0, roundConstant[3]}), .b ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, SboxOut[3]}), .c ({new_AGEMA_signal_5069, new_AGEMA_signal_5068, KeyArray_n51}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U32 ( .a ({new_AGEMA_signal_5071, new_AGEMA_signal_5070, KeyArray_n50}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, keyStateIn[2]}), .c ({new_AGEMA_signal_5105, new_AGEMA_signal_5104, KeyArray_inS30par[2]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U31 ( .a ({LMDPL_pre1, 1'b0, roundConstant[2]}), .b ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, SboxOut[2]}), .c ({new_AGEMA_signal_5071, new_AGEMA_signal_5070, KeyArray_n50}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U30 ( .a ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, KeyArray_n49}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .c ({new_AGEMA_signal_5107, new_AGEMA_signal_5106, KeyArray_inS30par[1]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U29 ( .a ({LMDPL_pre1, 1'b0, roundConstant[1]}), .b ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, SboxOut[1]}), .c ({new_AGEMA_signal_5073, new_AGEMA_signal_5072, KeyArray_n49}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U28 ( .a ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, KeyArray_n48}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, keyStateIn[0]}), .c ({new_AGEMA_signal_5075, new_AGEMA_signal_5074, KeyArray_inS30par[0]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) KeyArray_U27 ( .a ({LMDPL_pre1, 1'b0, roundConstant[0]}), .b ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, SboxOut[0]}), .c ({new_AGEMA_signal_5029, new_AGEMA_signal_5028, KeyArray_n48}) ) ;
    INV_X1 KeyArray_U26 ( .A (KeyArray_n47), .ZN (KeyArray_n46) ) ;
    INV_X1 KeyArray_U25 ( .A (KeyArray_n47), .ZN (KeyArray_n45) ) ;
    INV_X1 KeyArray_U24 ( .A (KeyArray_n47), .ZN (KeyArray_n44) ) ;
    INV_X1 KeyArray_U23 ( .A (KeyArray_n47), .ZN (KeyArray_n43) ) ;
    INV_X1 KeyArray_U22 ( .A (KeyArray_n47), .ZN (KeyArray_n42) ) ;
    INV_X1 KeyArray_U21 ( .A (KeyArray_n47), .ZN (KeyArray_n41) ) ;
    INV_X1 KeyArray_U20 ( .A (KeyArray_n47), .ZN (KeyArray_n40) ) ;
    INV_X1 KeyArray_U19 ( .A (KeyArray_n47), .ZN (KeyArray_n39) ) ;
    INV_X1 KeyArray_U18 ( .A (nReset), .ZN (KeyArray_n47) ) ;
    INV_X1 KeyArray_U17 ( .A (KeyArray_n38), .ZN (KeyArray_n31) ) ;
    INV_X1 KeyArray_U16 ( .A (KeyArray_n29), .ZN (KeyArray_n23) ) ;
    INV_X1 KeyArray_U15 ( .A (KeyArray_n38), .ZN (KeyArray_n37) ) ;
    INV_X1 KeyArray_U14 ( .A (KeyArray_n29), .ZN (KeyArray_n28) ) ;
    INV_X1 KeyArray_U13 ( .A (KeyArray_n38), .ZN (KeyArray_n36) ) ;
    INV_X1 KeyArray_U12 ( .A (KeyArray_n29), .ZN (KeyArray_n27) ) ;
    INV_X1 KeyArray_U11 ( .A (KeyArray_n38), .ZN (KeyArray_n35) ) ;
    INV_X1 KeyArray_U10 ( .A (KeyArray_n29), .ZN (KeyArray_n26) ) ;
    INV_X1 KeyArray_U9 ( .A (KeyArray_n38), .ZN (KeyArray_n32) ) ;
    INV_X1 KeyArray_U8 ( .A (KeyArray_n29), .ZN (KeyArray_n24) ) ;
    INV_X1 KeyArray_U7 ( .A (KeyArray_n38), .ZN (KeyArray_n33) ) ;
    INV_X1 KeyArray_U6 ( .A (KeyArray_n29), .ZN (KeyArray_n25) ) ;
    INV_X1 KeyArray_U5 ( .A (KeyArray_n38), .ZN (KeyArray_n30) ) ;
    INV_X1 KeyArray_U4 ( .A (KeyArray_n29), .ZN (KeyArray_n22) ) ;
    INV_X1 KeyArray_U3 ( .A (KeyArray_n38), .ZN (KeyArray_n34) ) ;
    INV_X1 KeyArray_U2 ( .A (selMC), .ZN (KeyArray_n38) ) ;
    INV_X1 KeyArray_U1 ( .A (n12), .ZN (KeyArray_n29) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, keyStateIn[0]}), .a ({new_AGEMA_signal_4637, new_AGEMA_signal_4636, KeyArray_S00reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, KeyArray_S00reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, KeyArray_inS00ser[0]}), .a ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, KeyArray_outS10ser[0]}), .c ({new_AGEMA_signal_4637, new_AGEMA_signal_4636, KeyArray_S00reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .a ({new_AGEMA_signal_4639, new_AGEMA_signal_4638, KeyArray_S00reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyArray_S00reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, KeyArray_inS00ser[1]}), .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, KeyArray_outS10ser[1]}), .c ({new_AGEMA_signal_4639, new_AGEMA_signal_4638, KeyArray_S00reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, keyStateIn[2]}), .a ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, KeyArray_S00reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4871, new_AGEMA_signal_4870, KeyArray_S00reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, KeyArray_inS00ser[2]}), .a ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KeyArray_outS10ser[2]}), .c ({new_AGEMA_signal_4641, new_AGEMA_signal_4640, KeyArray_S00reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, keyStateIn[3]}), .a ({new_AGEMA_signal_4643, new_AGEMA_signal_4642, KeyArray_S00reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, KeyArray_S00reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, KeyArray_inS00ser[3]}), .a ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, KeyArray_outS10ser[3]}), .c ({new_AGEMA_signal_4643, new_AGEMA_signal_4642, KeyArray_S00reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[4]}), .a ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, KeyArray_S00reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyArray_S00reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, KeyArray_inS00ser[4]}), .a ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, KeyArray_outS10ser[4]}), .c ({new_AGEMA_signal_4645, new_AGEMA_signal_4644, KeyArray_S00reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, keyStateIn[5]}), .a ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, KeyArray_S00reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4877, new_AGEMA_signal_4876, KeyArray_S00reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, KeyArray_inS00ser[5]}), .a ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, KeyArray_outS10ser[5]}), .c ({new_AGEMA_signal_4647, new_AGEMA_signal_4646, KeyArray_S00reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, keyStateIn[6]}), .a ({new_AGEMA_signal_4649, new_AGEMA_signal_4648, KeyArray_S00reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, KeyArray_S00reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, KeyArray_inS00ser[6]}), .a ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, KeyArray_outS10ser[6]}), .c ({new_AGEMA_signal_4649, new_AGEMA_signal_4648, KeyArray_S00reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[7]}), .a ({new_AGEMA_signal_4651, new_AGEMA_signal_4650, KeyArray_S00reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyArray_S00reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S00reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_4625, new_AGEMA_signal_4624, KeyArray_inS00ser[7]}), .a ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, KeyArray_outS10ser[7]}), .c ({new_AGEMA_signal_4651, new_AGEMA_signal_4650, KeyArray_S00reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, KeyArray_outS01ser_0_}), .a ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, KeyArray_S01reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4655, new_AGEMA_signal_4654, KeyArray_S01reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, KeyArray_inS01ser[0]}), .a ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, KeyArray_outS11ser[0]}), .c ({new_AGEMA_signal_3841, new_AGEMA_signal_3840, KeyArray_S01reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, KeyArray_outS01ser_1_}), .a ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, KeyArray_S01reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4657, new_AGEMA_signal_4656, KeyArray_S01reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, KeyArray_inS01ser[1]}), .a ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, KeyArray_outS11ser[1]}), .c ({new_AGEMA_signal_3843, new_AGEMA_signal_3842, KeyArray_S01reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_2_}), .a ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, KeyArray_S01reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, KeyArray_S01reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, KeyArray_inS01ser[2]}), .a ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, KeyArray_outS11ser[2]}), .c ({new_AGEMA_signal_3845, new_AGEMA_signal_3844, KeyArray_S01reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, KeyArray_outS01ser_3_}), .a ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, KeyArray_S01reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4661, new_AGEMA_signal_4660, KeyArray_S01reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, KeyArray_inS01ser[3]}), .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, KeyArray_outS11ser[3]}), .c ({new_AGEMA_signal_3847, new_AGEMA_signal_3846, KeyArray_S01reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, KeyArray_outS01ser_4_}), .a ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, KeyArray_S01reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4663, new_AGEMA_signal_4662, KeyArray_S01reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, KeyArray_inS01ser[4]}), .a ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, KeyArray_outS11ser[4]}), .c ({new_AGEMA_signal_3849, new_AGEMA_signal_3848, KeyArray_S01reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, KeyArray_outS01ser_5_}), .a ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, KeyArray_S01reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, KeyArray_S01reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, KeyArray_inS01ser[5]}), .a ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, KeyArray_outS11ser[5]}), .c ({new_AGEMA_signal_3851, new_AGEMA_signal_3850, KeyArray_S01reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, KeyArray_outS01ser_6_}), .a ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, KeyArray_S01reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4667, new_AGEMA_signal_4666, KeyArray_S01reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, KeyArray_inS01ser[6]}), .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, KeyArray_outS11ser[6]}), .c ({new_AGEMA_signal_3853, new_AGEMA_signal_3852, KeyArray_S01reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4653, new_AGEMA_signal_4652, KeyArray_n28}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, KeyArray_outS01ser_7_}), .a ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, KeyArray_S01reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyArray_S01reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S01reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3839, new_AGEMA_signal_3838, KeyArray_n37}), .b ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KeyArray_inS01ser[7]}), .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, KeyArray_outS11ser[7]}), .c ({new_AGEMA_signal_3855, new_AGEMA_signal_3854, KeyArray_S01reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, KeyArray_outS02ser[0]}), .a ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, KeyArray_S02reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4673, new_AGEMA_signal_4672, KeyArray_S02reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, KeyArray_inS02ser[0]}), .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, KeyArray_outS12ser[0]}), .c ({new_AGEMA_signal_3859, new_AGEMA_signal_3858, KeyArray_S02reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, KeyArray_outS02ser[1]}), .a ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, KeyArray_S02reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4675, new_AGEMA_signal_4674, KeyArray_S02reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, KeyArray_inS02ser[1]}), .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, KeyArray_outS12ser[1]}), .c ({new_AGEMA_signal_3861, new_AGEMA_signal_3860, KeyArray_S02reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, KeyArray_outS02ser[2]}), .a ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, KeyArray_S02reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, KeyArray_S02reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, KeyArray_inS02ser[2]}), .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, KeyArray_outS12ser[2]}), .c ({new_AGEMA_signal_3863, new_AGEMA_signal_3862, KeyArray_S02reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, KeyArray_outS02ser[3]}), .a ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, KeyArray_S02reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4679, new_AGEMA_signal_4678, KeyArray_S02reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, KeyArray_inS02ser[3]}), .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, KeyArray_outS12ser[3]}), .c ({new_AGEMA_signal_3865, new_AGEMA_signal_3864, KeyArray_S02reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, KeyArray_outS02ser[4]}), .a ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, KeyArray_S02reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4681, new_AGEMA_signal_4680, KeyArray_S02reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, KeyArray_inS02ser[4]}), .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, KeyArray_outS12ser[4]}), .c ({new_AGEMA_signal_3867, new_AGEMA_signal_3866, KeyArray_S02reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, KeyArray_outS02ser[5]}), .a ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, KeyArray_S02reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, KeyArray_S02reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, KeyArray_inS02ser[5]}), .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, KeyArray_outS12ser[5]}), .c ({new_AGEMA_signal_3869, new_AGEMA_signal_3868, KeyArray_S02reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, KeyArray_outS02ser[6]}), .a ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, KeyArray_S02reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4685, new_AGEMA_signal_4684, KeyArray_S02reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, KeyArray_inS02ser[6]}), .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, KeyArray_outS12ser[6]}), .c ({new_AGEMA_signal_3871, new_AGEMA_signal_3870, KeyArray_S02reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, KeyArray_outS02ser[7]}), .a ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, KeyArray_S02reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4687, new_AGEMA_signal_4686, KeyArray_S02reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S02reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, KeyArray_inS02ser[7]}), .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, KeyArray_outS12ser[7]}), .c ({new_AGEMA_signal_3873, new_AGEMA_signal_3872, KeyArray_S02reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, KeyArray_outS03ser[0]}), .a ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, KeyArray_S03reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, KeyArray_S03reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, KeyArray_inS03ser[0]}), .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, keySBIn[0]}), .c ({new_AGEMA_signal_3875, new_AGEMA_signal_3874, KeyArray_S03reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, KeyArray_outS03ser[1]}), .a ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, KeyArray_S03reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyArray_S03reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, KeyArray_inS03ser[1]}), .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, keySBIn[1]}), .c ({new_AGEMA_signal_3877, new_AGEMA_signal_3876, KeyArray_S03reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, KeyArray_outS03ser[2]}), .a ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, KeyArray_S03reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4693, new_AGEMA_signal_4692, KeyArray_S03reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, KeyArray_inS03ser[2]}), .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, keySBIn[2]}), .c ({new_AGEMA_signal_3879, new_AGEMA_signal_3878, KeyArray_S03reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, KeyArray_outS03ser[3]}), .a ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, KeyArray_S03reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, KeyArray_S03reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, KeyArray_inS03ser[3]}), .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, keySBIn[3]}), .c ({new_AGEMA_signal_3881, new_AGEMA_signal_3880, KeyArray_S03reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, KeyArray_outS03ser[4]}), .a ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, KeyArray_S03reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4697, new_AGEMA_signal_4696, KeyArray_S03reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, KeyArray_inS03ser[4]}), .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, keySBIn[4]}), .c ({new_AGEMA_signal_3883, new_AGEMA_signal_3882, KeyArray_S03reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, KeyArray_outS03ser[5]}), .a ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, KeyArray_S03reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4699, new_AGEMA_signal_4698, KeyArray_S03reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, KeyArray_inS03ser[5]}), .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, keySBIn[5]}), .c ({new_AGEMA_signal_3885, new_AGEMA_signal_3884, KeyArray_S03reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, KeyArray_outS03ser[6]}), .a ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, KeyArray_S03reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, KeyArray_S03reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, KeyArray_inS03ser[6]}), .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, keySBIn[6]}), .c ({new_AGEMA_signal_3887, new_AGEMA_signal_3886, KeyArray_S03reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4671, new_AGEMA_signal_4670, KeyArray_n27}), .b ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, KeyArray_outS03ser[7]}), .a ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, KeyArray_S03reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4703, new_AGEMA_signal_4702, KeyArray_S03reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S03reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3857, new_AGEMA_signal_3856, KeyArray_n36}), .b ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, KeyArray_inS03ser[7]}), .a ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, keySBIn[7]}), .c ({new_AGEMA_signal_3889, new_AGEMA_signal_3888, KeyArray_S03reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, KeyArray_outS10ser[0]}), .a ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, KeyArray_S10reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, KeyArray_S10reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, KeyArray_inS10ser[0]}), .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, KeyArray_outS20ser[0]}), .c ({new_AGEMA_signal_3893, new_AGEMA_signal_3892, KeyArray_S10reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, KeyArray_outS10ser[1]}), .a ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, KeyArray_S10reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4709, new_AGEMA_signal_4708, KeyArray_S10reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, KeyArray_inS10ser[1]}), .a ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, KeyArray_outS20ser[1]}), .c ({new_AGEMA_signal_3895, new_AGEMA_signal_3894, KeyArray_S10reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KeyArray_outS10ser[2]}), .a ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, KeyArray_S10reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4711, new_AGEMA_signal_4710, KeyArray_S10reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, KeyArray_inS10ser[2]}), .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, KeyArray_outS20ser[2]}), .c ({new_AGEMA_signal_3897, new_AGEMA_signal_3896, KeyArray_S10reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, KeyArray_outS10ser[3]}), .a ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, KeyArray_S10reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyArray_S10reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, KeyArray_inS10ser[3]}), .a ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, KeyArray_outS20ser[3]}), .c ({new_AGEMA_signal_3899, new_AGEMA_signal_3898, KeyArray_S10reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, KeyArray_outS10ser[4]}), .a ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, KeyArray_S10reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, KeyArray_S10reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, KeyArray_inS10ser[4]}), .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, KeyArray_outS20ser[4]}), .c ({new_AGEMA_signal_3901, new_AGEMA_signal_3900, KeyArray_S10reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, KeyArray_outS10ser[5]}), .a ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, KeyArray_S10reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, KeyArray_S10reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, KeyArray_inS10ser[5]}), .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, KeyArray_outS20ser[5]}), .c ({new_AGEMA_signal_3903, new_AGEMA_signal_3902, KeyArray_S10reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, KeyArray_outS10ser[6]}), .a ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, KeyArray_S10reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, KeyArray_S10reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, KeyArray_inS10ser[6]}), .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, KeyArray_outS20ser[6]}), .c ({new_AGEMA_signal_3905, new_AGEMA_signal_3904, KeyArray_S10reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, KeyArray_outS10ser[7]}), .a ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, KeyArray_S10reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, KeyArray_S10reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S10reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, KeyArray_inS10ser[7]}), .a ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, KeyArray_outS20ser[7]}), .c ({new_AGEMA_signal_3907, new_AGEMA_signal_3906, KeyArray_S10reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, KeyArray_outS11ser[0]}), .a ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, KeyArray_S11reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, KeyArray_S11reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, KeyArray_inS11ser[0]}), .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, KeyArray_outS21ser[0]}), .c ({new_AGEMA_signal_3909, new_AGEMA_signal_3908, KeyArray_S11reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, KeyArray_outS11ser[1]}), .a ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, KeyArray_S11reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, KeyArray_S11reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, KeyArray_inS11ser[1]}), .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, KeyArray_outS21ser[1]}), .c ({new_AGEMA_signal_3911, new_AGEMA_signal_3910, KeyArray_S11reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, KeyArray_outS11ser[2]}), .a ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, KeyArray_S11reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, KeyArray_S11reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, KeyArray_inS11ser[2]}), .a ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, KeyArray_outS21ser[2]}), .c ({new_AGEMA_signal_3913, new_AGEMA_signal_3912, KeyArray_S11reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, KeyArray_outS11ser[3]}), .a ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, KeyArray_S11reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyArray_S11reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, KeyArray_inS11ser[3]}), .a ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, KeyArray_outS21ser[3]}), .c ({new_AGEMA_signal_3915, new_AGEMA_signal_3914, KeyArray_S11reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, KeyArray_outS11ser[4]}), .a ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, KeyArray_S11reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyArray_S11reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, KeyArray_inS11ser[4]}), .a ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, KeyArray_outS21ser[4]}), .c ({new_AGEMA_signal_3917, new_AGEMA_signal_3916, KeyArray_S11reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, KeyArray_outS11ser[5]}), .a ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, KeyArray_S11reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyArray_S11reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, KeyArray_inS11ser[5]}), .a ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, KeyArray_outS21ser[5]}), .c ({new_AGEMA_signal_3919, new_AGEMA_signal_3918, KeyArray_S11reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, KeyArray_outS11ser[6]}), .a ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, KeyArray_S11reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyArray_S11reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, KeyArray_inS11ser[6]}), .a ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, KeyArray_outS21ser[6]}), .c ({new_AGEMA_signal_3921, new_AGEMA_signal_3920, KeyArray_S11reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4705, new_AGEMA_signal_4704, KeyArray_n26}), .b ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, KeyArray_outS11ser[7]}), .a ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, KeyArray_S11reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyArray_S11reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S11reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3891, new_AGEMA_signal_3890, KeyArray_n35}), .b ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, KeyArray_inS11ser[7]}), .a ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, KeyArray_outS21ser[7]}), .c ({new_AGEMA_signal_3923, new_AGEMA_signal_3922, KeyArray_S11reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, KeyArray_outS12ser[0]}), .a ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, KeyArray_S12reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, KeyArray_S12reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, KeyArray_inS12ser[0]}), .a ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, KeyArray_outS22ser[0]}), .c ({new_AGEMA_signal_3927, new_AGEMA_signal_3926, KeyArray_S12reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, KeyArray_outS12ser[1]}), .a ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, KeyArray_S12reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, KeyArray_S12reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, KeyArray_inS12ser[1]}), .a ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, KeyArray_outS22ser[1]}), .c ({new_AGEMA_signal_3929, new_AGEMA_signal_3928, KeyArray_S12reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, KeyArray_outS12ser[2]}), .a ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, KeyArray_S12reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, KeyArray_S12reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, KeyArray_inS12ser[2]}), .a ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, KeyArray_outS22ser[2]}), .c ({new_AGEMA_signal_3931, new_AGEMA_signal_3930, KeyArray_S12reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, KeyArray_outS12ser[3]}), .a ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, KeyArray_S12reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, KeyArray_S12reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, KeyArray_inS12ser[3]}), .a ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, KeyArray_outS22ser[3]}), .c ({new_AGEMA_signal_3933, new_AGEMA_signal_3932, KeyArray_S12reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, KeyArray_outS12ser[4]}), .a ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, KeyArray_S12reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, KeyArray_S12reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, KeyArray_inS12ser[4]}), .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, KeyArray_outS22ser[4]}), .c ({new_AGEMA_signal_3935, new_AGEMA_signal_3934, KeyArray_S12reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, KeyArray_outS12ser[5]}), .a ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, KeyArray_S12reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, KeyArray_S12reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, KeyArray_inS12ser[5]}), .a ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, KeyArray_outS22ser[5]}), .c ({new_AGEMA_signal_3937, new_AGEMA_signal_3936, KeyArray_S12reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, KeyArray_outS12ser[6]}), .a ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, KeyArray_S12reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, KeyArray_S12reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, KeyArray_inS12ser[6]}), .a ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, KeyArray_outS22ser[6]}), .c ({new_AGEMA_signal_3939, new_AGEMA_signal_3938, KeyArray_S12reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, KeyArray_outS12ser[7]}), .a ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, KeyArray_S12reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, KeyArray_S12reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S12reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, KeyArray_inS12ser[7]}), .a ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, KeyArray_outS22ser[7]}), .c ({new_AGEMA_signal_3941, new_AGEMA_signal_3940, KeyArray_S12reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, keySBIn[0]}), .a ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, KeyArray_S13reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, KeyArray_S13reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, KeyArray_inS13ser[0]}), .a ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, KeyArray_outS23ser[0]}), .c ({new_AGEMA_signal_3943, new_AGEMA_signal_3942, KeyArray_S13reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, keySBIn[1]}), .a ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, KeyArray_S13reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, KeyArray_S13reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, KeyArray_inS13ser[1]}), .a ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, KeyArray_outS23ser[1]}), .c ({new_AGEMA_signal_3945, new_AGEMA_signal_3944, KeyArray_S13reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, keySBIn[2]}), .a ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, KeyArray_S13reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4291, new_AGEMA_signal_4290, KeyArray_S13reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, KeyArray_inS13ser[2]}), .a ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, KeyArray_outS23ser[2]}), .c ({new_AGEMA_signal_3947, new_AGEMA_signal_3946, KeyArray_S13reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, keySBIn[3]}), .a ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, KeyArray_S13reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, KeyArray_S13reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, KeyArray_inS13ser[3]}), .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, KeyArray_outS23ser[3]}), .c ({new_AGEMA_signal_3949, new_AGEMA_signal_3948, KeyArray_S13reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, keySBIn[4]}), .a ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, KeyArray_S13reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4295, new_AGEMA_signal_4294, KeyArray_S13reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, KeyArray_inS13ser[4]}), .a ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, KeyArray_outS23ser[4]}), .c ({new_AGEMA_signal_3951, new_AGEMA_signal_3950, KeyArray_S13reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, keySBIn[5]}), .a ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, KeyArray_S13reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, KeyArray_S13reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, KeyArray_inS13ser[5]}), .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, KeyArray_outS23ser[5]}), .c ({new_AGEMA_signal_3953, new_AGEMA_signal_3952, KeyArray_S13reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, keySBIn[6]}), .a ({new_AGEMA_signal_3955, new_AGEMA_signal_3954, KeyArray_S13reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, KeyArray_S13reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, KeyArray_inS13ser[6]}), .a ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, KeyArray_outS23ser[6]}), .c ({new_AGEMA_signal_3955, new_AGEMA_signal_3954, KeyArray_S13reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4269, new_AGEMA_signal_4268, n12}), .b ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, keySBIn[7]}), .a ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, KeyArray_S13reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4301, new_AGEMA_signal_4300, KeyArray_S13reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S13reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3925, new_AGEMA_signal_3924, KeyArray_n34}), .b ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, KeyArray_inS13ser[7]}), .a ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, KeyArray_outS23ser[7]}), .c ({new_AGEMA_signal_3957, new_AGEMA_signal_3956, KeyArray_S13reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, KeyArray_outS20ser[0]}), .a ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, KeyArray_S20reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyArray_S20reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, KeyArray_inS20ser[0]}), .a ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, KeyArray_outS30ser[0]}), .c ({new_AGEMA_signal_3961, new_AGEMA_signal_3960, KeyArray_S20reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, KeyArray_outS20ser[1]}), .a ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, KeyArray_S20reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyArray_S20reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, KeyArray_inS20ser[1]}), .a ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, KeyArray_outS30ser[1]}), .c ({new_AGEMA_signal_3963, new_AGEMA_signal_3962, KeyArray_S20reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, KeyArray_outS20ser[2]}), .a ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, KeyArray_S20reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyArray_S20reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, KeyArray_inS20ser[2]}), .a ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, KeyArray_outS30ser[2]}), .c ({new_AGEMA_signal_3965, new_AGEMA_signal_3964, KeyArray_S20reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, KeyArray_outS20ser[3]}), .a ({new_AGEMA_signal_3967, new_AGEMA_signal_3966, KeyArray_S20reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyArray_S20reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, KeyArray_inS20ser[3]}), .a ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, KeyArray_outS30ser[3]}), .c ({new_AGEMA_signal_3967, new_AGEMA_signal_3966, KeyArray_S20reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, KeyArray_outS20ser[4]}), .a ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, KeyArray_S20reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyArray_S20reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, KeyArray_inS20ser[4]}), .a ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, KeyArray_outS30ser[4]}), .c ({new_AGEMA_signal_3969, new_AGEMA_signal_3968, KeyArray_S20reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, KeyArray_outS20ser[5]}), .a ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, KeyArray_S20reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyArray_S20reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, KeyArray_inS20ser[5]}), .a ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, KeyArray_outS30ser[5]}), .c ({new_AGEMA_signal_3971, new_AGEMA_signal_3970, KeyArray_S20reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, KeyArray_outS20ser[6]}), .a ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, KeyArray_S20reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyArray_S20reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, KeyArray_inS20ser[6]}), .a ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, KeyArray_outS30ser[6]}), .c ({new_AGEMA_signal_3973, new_AGEMA_signal_3972, KeyArray_S20reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, KeyArray_outS20ser[7]}), .a ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, KeyArray_S20reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyArray_S20reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S20reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, KeyArray_inS20ser[7]}), .a ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, KeyArray_outS30ser[7]}), .c ({new_AGEMA_signal_3975, new_AGEMA_signal_3974, KeyArray_S20reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, KeyArray_outS21ser[0]}), .a ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, KeyArray_S21reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyArray_S21reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, KeyArray_inS21ser[0]}), .a ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, KeyArray_outS31ser[0]}), .c ({new_AGEMA_signal_3977, new_AGEMA_signal_3976, KeyArray_S21reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, KeyArray_outS21ser[1]}), .a ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, KeyArray_S21reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyArray_S21reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, KeyArray_inS21ser[1]}), .a ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, KeyArray_outS31ser[1]}), .c ({new_AGEMA_signal_3979, new_AGEMA_signal_3978, KeyArray_S21reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, KeyArray_outS21ser[2]}), .a ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, KeyArray_S21reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyArray_S21reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, KeyArray_inS21ser[2]}), .a ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, KeyArray_outS31ser[2]}), .c ({new_AGEMA_signal_3981, new_AGEMA_signal_3980, KeyArray_S21reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, KeyArray_outS21ser[3]}), .a ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, KeyArray_S21reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyArray_S21reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, KeyArray_inS21ser[3]}), .a ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, KeyArray_outS31ser[3]}), .c ({new_AGEMA_signal_3983, new_AGEMA_signal_3982, KeyArray_S21reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, KeyArray_outS21ser[4]}), .a ({new_AGEMA_signal_3985, new_AGEMA_signal_3984, KeyArray_S21reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyArray_S21reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, KeyArray_inS21ser[4]}), .a ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, KeyArray_outS31ser[4]}), .c ({new_AGEMA_signal_3985, new_AGEMA_signal_3984, KeyArray_S21reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, KeyArray_outS21ser[5]}), .a ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, KeyArray_S21reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyArray_S21reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, KeyArray_inS21ser[5]}), .a ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, KeyArray_outS31ser[5]}), .c ({new_AGEMA_signal_3987, new_AGEMA_signal_3986, KeyArray_S21reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, KeyArray_outS21ser[6]}), .a ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, KeyArray_S21reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyArray_S21reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, KeyArray_inS21ser[6]}), .a ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, KeyArray_outS31ser[6]}), .c ({new_AGEMA_signal_3989, new_AGEMA_signal_3988, KeyArray_S21reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4739, new_AGEMA_signal_4738, KeyArray_n25}), .b ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, KeyArray_outS21ser[7]}), .a ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, KeyArray_S21reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, KeyArray_S21reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S21reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3959, new_AGEMA_signal_3958, KeyArray_n33}), .b ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, KeyArray_inS21ser[7]}), .a ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, KeyArray_outS31ser[7]}), .c ({new_AGEMA_signal_3991, new_AGEMA_signal_3990, KeyArray_S21reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, KeyArray_outS22ser[0]}), .a ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, KeyArray_S22reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4775, new_AGEMA_signal_4774, KeyArray_S22reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, KeyArray_inS22ser[0]}), .a ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, KeyArray_outS32ser[0]}), .c ({new_AGEMA_signal_3995, new_AGEMA_signal_3994, KeyArray_S22reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, KeyArray_outS22ser[1]}), .a ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, KeyArray_S22reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4777, new_AGEMA_signal_4776, KeyArray_S22reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, KeyArray_inS22ser[1]}), .a ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, KeyArray_outS32ser[1]}), .c ({new_AGEMA_signal_3997, new_AGEMA_signal_3996, KeyArray_S22reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, KeyArray_outS22ser[2]}), .a ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, KeyArray_S22reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, KeyArray_S22reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, KeyArray_inS22ser[2]}), .a ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, KeyArray_outS32ser[2]}), .c ({new_AGEMA_signal_3999, new_AGEMA_signal_3998, KeyArray_S22reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, KeyArray_outS22ser[3]}), .a ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, KeyArray_S22reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4781, new_AGEMA_signal_4780, KeyArray_S22reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, KeyArray_inS22ser[3]}), .a ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, KeyArray_outS32ser[3]}), .c ({new_AGEMA_signal_4001, new_AGEMA_signal_4000, KeyArray_S22reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, KeyArray_outS22ser[4]}), .a ({new_AGEMA_signal_4003, new_AGEMA_signal_4002, KeyArray_S22reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, KeyArray_S22reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, KeyArray_inS22ser[4]}), .a ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, KeyArray_outS32ser[4]}), .c ({new_AGEMA_signal_4003, new_AGEMA_signal_4002, KeyArray_S22reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, KeyArray_outS22ser[5]}), .a ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, KeyArray_S22reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, KeyArray_S22reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, KeyArray_inS22ser[5]}), .a ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, KeyArray_outS32ser[5]}), .c ({new_AGEMA_signal_4005, new_AGEMA_signal_4004, KeyArray_S22reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, KeyArray_outS22ser[6]}), .a ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, KeyArray_S22reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4787, new_AGEMA_signal_4786, KeyArray_S22reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, KeyArray_inS22ser[6]}), .a ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, KeyArray_outS32ser[6]}), .c ({new_AGEMA_signal_4007, new_AGEMA_signal_4006, KeyArray_S22reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, KeyArray_outS22ser[7]}), .a ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, KeyArray_S22reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, KeyArray_S22reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S22reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, KeyArray_inS22ser[7]}), .a ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, KeyArray_outS32ser[7]}), .c ({new_AGEMA_signal_4009, new_AGEMA_signal_4008, KeyArray_S22reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, KeyArray_outS23ser[0]}), .a ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, KeyArray_S23reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, KeyArray_S23reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, KeyArray_inS23ser[0]}), .a ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, KeyArray_outS33ser[0]}), .c ({new_AGEMA_signal_4011, new_AGEMA_signal_4010, KeyArray_S23reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, KeyArray_outS23ser[1]}), .a ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, KeyArray_S23reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4793, new_AGEMA_signal_4792, KeyArray_S23reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, KeyArray_inS23ser[1]}), .a ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, KeyArray_outS33ser[1]}), .c ({new_AGEMA_signal_4013, new_AGEMA_signal_4012, KeyArray_S23reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, KeyArray_outS23ser[2]}), .a ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, KeyArray_S23reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, KeyArray_S23reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, KeyArray_inS23ser[2]}), .a ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, KeyArray_outS33ser[2]}), .c ({new_AGEMA_signal_4015, new_AGEMA_signal_4014, KeyArray_S23reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, KeyArray_outS23ser[3]}), .a ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, KeyArray_S23reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, KeyArray_S23reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, KeyArray_inS23ser[3]}), .a ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, KeyArray_outS33ser[3]}), .c ({new_AGEMA_signal_4017, new_AGEMA_signal_4016, KeyArray_S23reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, KeyArray_outS23ser[4]}), .a ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, KeyArray_S23reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4799, new_AGEMA_signal_4798, KeyArray_S23reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, KeyArray_inS23ser[4]}), .a ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, KeyArray_outS33ser[4]}), .c ({new_AGEMA_signal_4019, new_AGEMA_signal_4018, KeyArray_S23reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, KeyArray_outS23ser[5]}), .a ({new_AGEMA_signal_4021, new_AGEMA_signal_4020, KeyArray_S23reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, KeyArray_S23reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, KeyArray_inS23ser[5]}), .a ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, KeyArray_outS33ser[5]}), .c ({new_AGEMA_signal_4021, new_AGEMA_signal_4020, KeyArray_S23reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, KeyArray_outS23ser[6]}), .a ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, KeyArray_S23reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, KeyArray_S23reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, KeyArray_inS23ser[6]}), .a ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, KeyArray_outS33ser[6]}), .c ({new_AGEMA_signal_4023, new_AGEMA_signal_4022, KeyArray_S23reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4773, new_AGEMA_signal_4772, KeyArray_n24}), .b ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, KeyArray_outS23ser[7]}), .a ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, KeyArray_S23reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4805, new_AGEMA_signal_4804, KeyArray_S23reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S23reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_3993, new_AGEMA_signal_3992, KeyArray_n32}), .b ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, KeyArray_inS23ser[7]}), .a ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, KeyArray_outS33ser[7]}), .c ({new_AGEMA_signal_4025, new_AGEMA_signal_4024, KeyArray_S23reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, KeyArray_outS30ser[0]}), .a ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, KeyArray_S30reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_5141, new_AGEMA_signal_5140, KeyArray_S30reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, KeyArray_inS30ser[0]}), .a ({new_AGEMA_signal_5075, new_AGEMA_signal_5074, KeyArray_inS30par[0]}), .c ({new_AGEMA_signal_5109, new_AGEMA_signal_5108, KeyArray_S30reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, KeyArray_outS30ser[1]}), .a ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, KeyArray_S30reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_5171, new_AGEMA_signal_5170, KeyArray_S30reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, KeyArray_inS30ser[1]}), .a ({new_AGEMA_signal_5107, new_AGEMA_signal_5106, KeyArray_inS30par[1]}), .c ({new_AGEMA_signal_5143, new_AGEMA_signal_5142, KeyArray_S30reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, KeyArray_outS30ser[2]}), .a ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, KeyArray_S30reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_5173, new_AGEMA_signal_5172, KeyArray_S30reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, KeyArray_inS30ser[2]}), .a ({new_AGEMA_signal_5105, new_AGEMA_signal_5104, KeyArray_inS30par[2]}), .c ({new_AGEMA_signal_5145, new_AGEMA_signal_5144, KeyArray_S30reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, KeyArray_outS30ser[3]}), .a ({new_AGEMA_signal_5147, new_AGEMA_signal_5146, KeyArray_S30reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, KeyArray_S30reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, KeyArray_inS30ser[3]}), .a ({new_AGEMA_signal_5103, new_AGEMA_signal_5102, KeyArray_inS30par[3]}), .c ({new_AGEMA_signal_5147, new_AGEMA_signal_5146, KeyArray_S30reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, KeyArray_outS30ser[4]}), .a ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, KeyArray_S30reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_5177, new_AGEMA_signal_5176, KeyArray_S30reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, KeyArray_inS30ser[4]}), .a ({new_AGEMA_signal_5101, new_AGEMA_signal_5100, KeyArray_inS30par[4]}), .c ({new_AGEMA_signal_5149, new_AGEMA_signal_5148, KeyArray_S30reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, KeyArray_outS30ser[5]}), .a ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, KeyArray_S30reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_5179, new_AGEMA_signal_5178, KeyArray_S30reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, KeyArray_inS30ser[5]}), .a ({new_AGEMA_signal_5099, new_AGEMA_signal_5098, KeyArray_inS30par[5]}), .c ({new_AGEMA_signal_5151, new_AGEMA_signal_5150, KeyArray_S30reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, KeyArray_outS30ser[6]}), .a ({new_AGEMA_signal_5153, new_AGEMA_signal_5152, KeyArray_S30reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, KeyArray_S30reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, KeyArray_inS30ser[6]}), .a ({new_AGEMA_signal_5097, new_AGEMA_signal_5096, KeyArray_inS30par[6]}), .c ({new_AGEMA_signal_5153, new_AGEMA_signal_5152, KeyArray_S30reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, KeyArray_outS30ser[7]}), .a ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, KeyArray_S30reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_5183, new_AGEMA_signal_5182, KeyArray_S30reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S30reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, KeyArray_inS30ser[7]}), .a ({new_AGEMA_signal_5095, new_AGEMA_signal_5094, KeyArray_inS30par[7]}), .c ({new_AGEMA_signal_5155, new_AGEMA_signal_5154, KeyArray_S30reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, KeyArray_outS31ser[0]}), .a ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, KeyArray_S31reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, KeyArray_S31reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, KeyArray_inS31ser[0]}), .a ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, KeyArray_outS01ser_0_}), .c ({new_AGEMA_signal_4029, new_AGEMA_signal_4028, KeyArray_S31reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, KeyArray_outS31ser[1]}), .a ({new_AGEMA_signal_4031, new_AGEMA_signal_4030, KeyArray_S31reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4811, new_AGEMA_signal_4810, KeyArray_S31reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, KeyArray_inS31ser[1]}), .a ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, KeyArray_outS01ser_1_}), .c ({new_AGEMA_signal_4031, new_AGEMA_signal_4030, KeyArray_S31reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, KeyArray_outS31ser[2]}), .a ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, KeyArray_S31reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, KeyArray_S31reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, KeyArray_inS31ser[2]}), .a ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_2_}), .c ({new_AGEMA_signal_4033, new_AGEMA_signal_4032, KeyArray_S31reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, KeyArray_outS31ser[3]}), .a ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, KeyArray_S31reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, KeyArray_S31reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, KeyArray_inS31ser[3]}), .a ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, KeyArray_outS01ser_3_}), .c ({new_AGEMA_signal_4035, new_AGEMA_signal_4034, KeyArray_S31reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, KeyArray_outS31ser[4]}), .a ({new_AGEMA_signal_4037, new_AGEMA_signal_4036, KeyArray_S31reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4817, new_AGEMA_signal_4816, KeyArray_S31reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, KeyArray_inS31ser[4]}), .a ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, KeyArray_outS01ser_4_}), .c ({new_AGEMA_signal_4037, new_AGEMA_signal_4036, KeyArray_S31reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, KeyArray_outS31ser[5]}), .a ({new_AGEMA_signal_4039, new_AGEMA_signal_4038, KeyArray_S31reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4819, new_AGEMA_signal_4818, KeyArray_S31reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, KeyArray_inS31ser[5]}), .a ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, KeyArray_outS01ser_5_}), .c ({new_AGEMA_signal_4039, new_AGEMA_signal_4038, KeyArray_S31reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, KeyArray_outS31ser[6]}), .a ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, KeyArray_S31reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, KeyArray_S31reg_gff_1_SFF_6_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, KeyArray_inS31ser[6]}), .a ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, KeyArray_outS01ser_6_}), .c ({new_AGEMA_signal_4041, new_AGEMA_signal_4040, KeyArray_S31reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4807, new_AGEMA_signal_4806, KeyArray_n23}), .b ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, KeyArray_outS31ser[7]}), .a ({new_AGEMA_signal_4043, new_AGEMA_signal_4042, KeyArray_S31reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4823, new_AGEMA_signal_4822, KeyArray_S31reg_gff_1_SFF_7_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S31reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4027, new_AGEMA_signal_4026, KeyArray_n31}), .b ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, KeyArray_inS31ser[7]}), .a ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, KeyArray_outS01ser_7_}), .c ({new_AGEMA_signal_4043, new_AGEMA_signal_4042, KeyArray_S31reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, KeyArray_outS32ser[0]}), .a ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, KeyArray_S32reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, KeyArray_S32reg_gff_1_SFF_0_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, KeyArray_inS32ser[0]}), .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, KeyArray_outS02ser[0]}), .c ({new_AGEMA_signal_4047, new_AGEMA_signal_4046, KeyArray_S32reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, KeyArray_outS32ser[1]}), .a ({new_AGEMA_signal_4049, new_AGEMA_signal_4048, KeyArray_S32reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4829, new_AGEMA_signal_4828, KeyArray_S32reg_gff_1_SFF_1_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, KeyArray_inS32ser[1]}), .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, KeyArray_outS02ser[1]}), .c ({new_AGEMA_signal_4049, new_AGEMA_signal_4048, KeyArray_S32reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, KeyArray_outS32ser[2]}), .a ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, KeyArray_S32reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4831, new_AGEMA_signal_4830, KeyArray_S32reg_gff_1_SFF_2_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, KeyArray_inS32ser[2]}), .a ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, KeyArray_outS02ser[2]}), .c ({new_AGEMA_signal_4051, new_AGEMA_signal_4050, KeyArray_S32reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, KeyArray_outS32ser[3]}), .a ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, KeyArray_S32reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, KeyArray_S32reg_gff_1_SFF_3_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, KeyArray_inS32ser[3]}), .a ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, KeyArray_outS02ser[3]}), .c ({new_AGEMA_signal_4053, new_AGEMA_signal_4052, KeyArray_S32reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, KeyArray_outS32ser[4]}), .a ({new_AGEMA_signal_4055, new_AGEMA_signal_4054, KeyArray_S32reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4835, new_AGEMA_signal_4834, KeyArray_S32reg_gff_1_SFF_4_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, KeyArray_inS32ser[4]}), .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, KeyArray_outS02ser[4]}), .c ({new_AGEMA_signal_4055, new_AGEMA_signal_4054, KeyArray_S32reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, KeyArray_outS32ser[5]}), .a ({new_AGEMA_signal_4057, new_AGEMA_signal_4056, KeyArray_S32reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4837, new_AGEMA_signal_4836, KeyArray_S32reg_gff_1_SFF_5_n6}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, KeyArray_inS32ser[5]}), .a ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, KeyArray_outS02ser[5]}), .c ({new_AGEMA_signal_4057, new_AGEMA_signal_4056, KeyArray_S32reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, KeyArray_outS32ser[6]}), .a ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, KeyArray_S32reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, KeyArray_S32reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, KeyArray_inS32ser[6]}), .a ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, KeyArray_outS02ser[6]}), .c ({new_AGEMA_signal_4059, new_AGEMA_signal_4058, KeyArray_S32reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, KeyArray_outS32ser[7]}), .a ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, KeyArray_S32reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4841, new_AGEMA_signal_4840, KeyArray_S32reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S32reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, KeyArray_inS32ser[7]}), .a ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, KeyArray_outS02ser[7]}), .c ({new_AGEMA_signal_4061, new_AGEMA_signal_4060, KeyArray_S32reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_0_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, KeyArray_outS33ser[0]}), .a ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, KeyArray_S33reg_gff_1_SFF_0_QD}), .c ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, KeyArray_S33reg_gff_1_SFF_0_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_0_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, KeyArray_inS33ser[0]}), .a ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, KeyArray_outS03ser[0]}), .c ({new_AGEMA_signal_4063, new_AGEMA_signal_4062, KeyArray_S33reg_gff_1_SFF_0_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_1_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, KeyArray_outS33ser[1]}), .a ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, KeyArray_S33reg_gff_1_SFF_1_QD}), .c ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyArray_S33reg_gff_1_SFF_1_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_1_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, KeyArray_inS33ser[1]}), .a ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, KeyArray_outS03ser[1]}), .c ({new_AGEMA_signal_4065, new_AGEMA_signal_4064, KeyArray_S33reg_gff_1_SFF_1_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_2_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, KeyArray_outS33ser[2]}), .a ({new_AGEMA_signal_4067, new_AGEMA_signal_4066, KeyArray_S33reg_gff_1_SFF_2_QD}), .c ({new_AGEMA_signal_4847, new_AGEMA_signal_4846, KeyArray_S33reg_gff_1_SFF_2_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_2_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, KeyArray_inS33ser[2]}), .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, KeyArray_outS03ser[2]}), .c ({new_AGEMA_signal_4067, new_AGEMA_signal_4066, KeyArray_S33reg_gff_1_SFF_2_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_3_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, KeyArray_outS33ser[3]}), .a ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, KeyArray_S33reg_gff_1_SFF_3_QD}), .c ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, KeyArray_S33reg_gff_1_SFF_3_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_3_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, KeyArray_inS33ser[3]}), .a ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, KeyArray_outS03ser[3]}), .c ({new_AGEMA_signal_4069, new_AGEMA_signal_4068, KeyArray_S33reg_gff_1_SFF_3_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_4_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, KeyArray_outS33ser[4]}), .a ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, KeyArray_S33reg_gff_1_SFF_4_QD}), .c ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyArray_S33reg_gff_1_SFF_4_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_4_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, KeyArray_inS33ser[4]}), .a ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, KeyArray_outS03ser[4]}), .c ({new_AGEMA_signal_4071, new_AGEMA_signal_4070, KeyArray_S33reg_gff_1_SFF_4_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_5_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, KeyArray_outS33ser[5]}), .a ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, KeyArray_S33reg_gff_1_SFF_5_QD}), .c ({new_AGEMA_signal_4853, new_AGEMA_signal_4852, KeyArray_S33reg_gff_1_SFF_5_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_5_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, KeyArray_inS33ser[5]}), .a ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, KeyArray_outS03ser[5]}), .c ({new_AGEMA_signal_4073, new_AGEMA_signal_4072, KeyArray_S33reg_gff_1_SFF_5_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_6_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, KeyArray_outS33ser[6]}), .a ({new_AGEMA_signal_4075, new_AGEMA_signal_4074, KeyArray_S33reg_gff_1_SFF_6_QD}), .c ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, KeyArray_S33reg_gff_1_SFF_6_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_6_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, KeyArray_inS33ser[6]}), .a ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, KeyArray_outS03ser[6]}), .c ({new_AGEMA_signal_4075, new_AGEMA_signal_4074, KeyArray_S33reg_gff_1_SFF_6_QD}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_7_U1 ( .s ({new_AGEMA_signal_4825, new_AGEMA_signal_4824, KeyArray_n22}), .b ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, KeyArray_outS33ser[7]}), .a ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, KeyArray_S33reg_gff_1_SFF_7_QD}), .c ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyArray_S33reg_gff_1_SFF_7_n5}) ) ;
    mux2_masked_LMDPL KeyArray_S33reg_gff_1_SFF_7_MUXInst_U1 ( .s ({new_AGEMA_signal_4045, new_AGEMA_signal_4044, KeyArray_n30}), .b ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, KeyArray_inS33ser[7]}), .a ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, KeyArray_outS03ser[7]}), .c ({new_AGEMA_signal_4077, new_AGEMA_signal_4076, KeyArray_S33reg_gff_1_SFF_7_QD}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_selXOR_mux_inst_0_U1 ( .s ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, intselXOR}), .b ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, KeyArray_outS01ser_0_}), .a ({new_AGEMA_signal_2065, new_AGEMA_signal_2064, KeyArray_outS01ser_XOR_00[0]}), .c ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, KeyArray_outS01ser_p[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_selXOR_mux_inst_1_U1 ( .s ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, intselXOR}), .b ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, KeyArray_outS01ser_1_}), .a ({new_AGEMA_signal_2061, new_AGEMA_signal_2060, KeyArray_outS01ser_XOR_00[1]}), .c ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, KeyArray_outS01ser_p[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_selXOR_mux_inst_2_U1 ( .s ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, intselXOR}), .b ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_2_}), .a ({new_AGEMA_signal_2057, new_AGEMA_signal_2056, KeyArray_outS01ser_XOR_00[2]}), .c ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, KeyArray_outS01ser_p[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_selXOR_mux_inst_3_U1 ( .s ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, intselXOR}), .b ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, KeyArray_outS01ser_3_}), .a ({new_AGEMA_signal_2053, new_AGEMA_signal_2052, KeyArray_outS01ser_XOR_00[3]}), .c ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, KeyArray_outS01ser_p[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_selXOR_mux_inst_4_U1 ( .s ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, intselXOR}), .b ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, KeyArray_outS01ser_4_}), .a ({new_AGEMA_signal_2049, new_AGEMA_signal_2048, KeyArray_outS01ser_XOR_00[4]}), .c ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, KeyArray_outS01ser_p[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_selXOR_mux_inst_5_U1 ( .s ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, intselXOR}), .b ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, KeyArray_outS01ser_5_}), .a ({new_AGEMA_signal_2045, new_AGEMA_signal_2044, KeyArray_outS01ser_XOR_00[5]}), .c ({new_AGEMA_signal_4315, new_AGEMA_signal_4314, KeyArray_outS01ser_p[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_selXOR_mux_inst_6_U1 ( .s ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, intselXOR}), .b ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, KeyArray_outS01ser_6_}), .a ({new_AGEMA_signal_2041, new_AGEMA_signal_2040, KeyArray_outS01ser_XOR_00[6]}), .c ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, KeyArray_outS01ser_p[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_selXOR_mux_inst_7_U1 ( .s ({new_AGEMA_signal_4303, new_AGEMA_signal_4302, intselXOR}), .b ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, KeyArray_outS01ser_7_}), .a ({new_AGEMA_signal_2037, new_AGEMA_signal_2036, KeyArray_outS01ser_XOR_00[7]}), .c ({new_AGEMA_signal_4319, new_AGEMA_signal_4318, KeyArray_outS01ser_p[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS00ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_4595, new_AGEMA_signal_4594, key_s0[120]}), .a ({new_AGEMA_signal_4305, new_AGEMA_signal_4304, KeyArray_outS01ser_p[0]}), .c ({new_AGEMA_signal_4597, new_AGEMA_signal_4596, KeyArray_inS00ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS00ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_4599, new_AGEMA_signal_4598, key_s0[121]}), .a ({new_AGEMA_signal_4307, new_AGEMA_signal_4306, KeyArray_outS01ser_p[1]}), .c ({new_AGEMA_signal_4601, new_AGEMA_signal_4600, KeyArray_inS00ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS00ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_4603, new_AGEMA_signal_4602, key_s0[122]}), .a ({new_AGEMA_signal_4309, new_AGEMA_signal_4308, KeyArray_outS01ser_p[2]}), .c ({new_AGEMA_signal_4605, new_AGEMA_signal_4604, KeyArray_inS00ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS00ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_4607, new_AGEMA_signal_4606, key_s0[123]}), .a ({new_AGEMA_signal_4311, new_AGEMA_signal_4310, KeyArray_outS01ser_p[3]}), .c ({new_AGEMA_signal_4609, new_AGEMA_signal_4608, KeyArray_inS00ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS00ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_4611, new_AGEMA_signal_4610, key_s0[124]}), .a ({new_AGEMA_signal_4313, new_AGEMA_signal_4312, KeyArray_outS01ser_p[4]}), .c ({new_AGEMA_signal_4613, new_AGEMA_signal_4612, KeyArray_inS00ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS00ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_4615, new_AGEMA_signal_4614, key_s0[125]}), .a ({new_AGEMA_signal_4315, new_AGEMA_signal_4314, KeyArray_outS01ser_p[5]}), .c ({new_AGEMA_signal_4617, new_AGEMA_signal_4616, KeyArray_inS00ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS00ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_4619, new_AGEMA_signal_4618, key_s0[126]}), .a ({new_AGEMA_signal_4317, new_AGEMA_signal_4316, KeyArray_outS01ser_p[6]}), .c ({new_AGEMA_signal_4621, new_AGEMA_signal_4620, KeyArray_inS00ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS00ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_4623, new_AGEMA_signal_4622, key_s0[127]}), .a ({new_AGEMA_signal_4319, new_AGEMA_signal_4318, KeyArray_outS01ser_p[7]}), .c ({new_AGEMA_signal_4625, new_AGEMA_signal_4624, KeyArray_inS00ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS01ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_2925, new_AGEMA_signal_2924, key_s0[112]}), .a ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, KeyArray_outS02ser[0]}), .c ({new_AGEMA_signal_2929, new_AGEMA_signal_2928, KeyArray_inS01ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS01ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_2931, new_AGEMA_signal_2930, key_s0[113]}), .a ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, KeyArray_outS02ser[1]}), .c ({new_AGEMA_signal_2935, new_AGEMA_signal_2934, KeyArray_inS01ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS01ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_2937, new_AGEMA_signal_2936, key_s0[114]}), .a ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, KeyArray_outS02ser[2]}), .c ({new_AGEMA_signal_2941, new_AGEMA_signal_2940, KeyArray_inS01ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS01ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_2943, new_AGEMA_signal_2942, key_s0[115]}), .a ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, KeyArray_outS02ser[3]}), .c ({new_AGEMA_signal_2947, new_AGEMA_signal_2946, KeyArray_inS01ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS01ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_2949, new_AGEMA_signal_2948, key_s0[116]}), .a ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, KeyArray_outS02ser[4]}), .c ({new_AGEMA_signal_2953, new_AGEMA_signal_2952, KeyArray_inS01ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS01ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_2955, new_AGEMA_signal_2954, key_s0[117]}), .a ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, KeyArray_outS02ser[5]}), .c ({new_AGEMA_signal_2959, new_AGEMA_signal_2958, KeyArray_inS01ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS01ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_2961, new_AGEMA_signal_2960, key_s0[118]}), .a ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, KeyArray_outS02ser[6]}), .c ({new_AGEMA_signal_2965, new_AGEMA_signal_2964, KeyArray_inS01ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS01ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2923, new_AGEMA_signal_2922, KeyArray_n46}), .b ({new_AGEMA_signal_2967, new_AGEMA_signal_2966, key_s0[119]}), .a ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, KeyArray_outS02ser[7]}), .c ({new_AGEMA_signal_2971, new_AGEMA_signal_2970, KeyArray_inS01ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS02ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_2975, new_AGEMA_signal_2974, key_s0[104]}), .a ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, KeyArray_outS03ser[0]}), .c ({new_AGEMA_signal_2979, new_AGEMA_signal_2978, KeyArray_inS02ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS02ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_2981, new_AGEMA_signal_2980, key_s0[105]}), .a ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, KeyArray_outS03ser[1]}), .c ({new_AGEMA_signal_2985, new_AGEMA_signal_2984, KeyArray_inS02ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS02ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_2987, new_AGEMA_signal_2986, key_s0[106]}), .a ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, KeyArray_outS03ser[2]}), .c ({new_AGEMA_signal_2991, new_AGEMA_signal_2990, KeyArray_inS02ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS02ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_2993, new_AGEMA_signal_2992, key_s0[107]}), .a ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, KeyArray_outS03ser[3]}), .c ({new_AGEMA_signal_2997, new_AGEMA_signal_2996, KeyArray_inS02ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS02ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_2999, new_AGEMA_signal_2998, key_s0[108]}), .a ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, KeyArray_outS03ser[4]}), .c ({new_AGEMA_signal_3003, new_AGEMA_signal_3002, KeyArray_inS02ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS02ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3005, new_AGEMA_signal_3004, key_s0[109]}), .a ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, KeyArray_outS03ser[5]}), .c ({new_AGEMA_signal_3009, new_AGEMA_signal_3008, KeyArray_inS02ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS02ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3011, new_AGEMA_signal_3010, key_s0[110]}), .a ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, KeyArray_outS03ser[6]}), .c ({new_AGEMA_signal_3015, new_AGEMA_signal_3014, KeyArray_inS02ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS02ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3017, new_AGEMA_signal_3016, key_s0[111]}), .a ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, KeyArray_outS03ser[7]}), .c ({new_AGEMA_signal_3021, new_AGEMA_signal_3020, KeyArray_inS02ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS03ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3023, new_AGEMA_signal_3022, key_s0[96]}), .a ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, KeyArray_outS10ser[0]}), .c ({new_AGEMA_signal_3027, new_AGEMA_signal_3026, KeyArray_inS03ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS03ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3029, new_AGEMA_signal_3028, key_s0[97]}), .a ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, KeyArray_outS10ser[1]}), .c ({new_AGEMA_signal_3033, new_AGEMA_signal_3032, KeyArray_inS03ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS03ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3035, new_AGEMA_signal_3034, key_s0[98]}), .a ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KeyArray_outS10ser[2]}), .c ({new_AGEMA_signal_3039, new_AGEMA_signal_3038, KeyArray_inS03ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS03ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3041, new_AGEMA_signal_3040, key_s0[99]}), .a ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, KeyArray_outS10ser[3]}), .c ({new_AGEMA_signal_3045, new_AGEMA_signal_3044, KeyArray_inS03ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS03ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3047, new_AGEMA_signal_3046, key_s0[100]}), .a ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, KeyArray_outS10ser[4]}), .c ({new_AGEMA_signal_3051, new_AGEMA_signal_3050, KeyArray_inS03ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS03ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3053, new_AGEMA_signal_3052, key_s0[101]}), .a ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, KeyArray_outS10ser[5]}), .c ({new_AGEMA_signal_3057, new_AGEMA_signal_3056, KeyArray_inS03ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS03ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3059, new_AGEMA_signal_3058, key_s0[102]}), .a ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, KeyArray_outS10ser[6]}), .c ({new_AGEMA_signal_3063, new_AGEMA_signal_3062, KeyArray_inS03ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS03ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_2973, new_AGEMA_signal_2972, KeyArray_n45}), .b ({new_AGEMA_signal_3065, new_AGEMA_signal_3064, key_s0[103]}), .a ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, KeyArray_outS10ser[7]}), .c ({new_AGEMA_signal_3069, new_AGEMA_signal_3068, KeyArray_inS03ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS10ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3073, new_AGEMA_signal_3072, key_s0[88]}), .a ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, KeyArray_outS11ser[0]}), .c ({new_AGEMA_signal_3077, new_AGEMA_signal_3076, KeyArray_inS10ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS10ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3079, new_AGEMA_signal_3078, key_s0[89]}), .a ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, KeyArray_outS11ser[1]}), .c ({new_AGEMA_signal_3083, new_AGEMA_signal_3082, KeyArray_inS10ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS10ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3085, new_AGEMA_signal_3084, key_s0[90]}), .a ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, KeyArray_outS11ser[2]}), .c ({new_AGEMA_signal_3089, new_AGEMA_signal_3088, KeyArray_inS10ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS10ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3091, new_AGEMA_signal_3090, key_s0[91]}), .a ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, KeyArray_outS11ser[3]}), .c ({new_AGEMA_signal_3095, new_AGEMA_signal_3094, KeyArray_inS10ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS10ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3097, new_AGEMA_signal_3096, key_s0[92]}), .a ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, KeyArray_outS11ser[4]}), .c ({new_AGEMA_signal_3101, new_AGEMA_signal_3100, KeyArray_inS10ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS10ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3103, new_AGEMA_signal_3102, key_s0[93]}), .a ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, KeyArray_outS11ser[5]}), .c ({new_AGEMA_signal_3107, new_AGEMA_signal_3106, KeyArray_inS10ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS10ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3109, new_AGEMA_signal_3108, key_s0[94]}), .a ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, KeyArray_outS11ser[6]}), .c ({new_AGEMA_signal_3113, new_AGEMA_signal_3112, KeyArray_inS10ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS10ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3115, new_AGEMA_signal_3114, key_s0[95]}), .a ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, KeyArray_outS11ser[7]}), .c ({new_AGEMA_signal_3119, new_AGEMA_signal_3118, KeyArray_inS10ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS11ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3121, new_AGEMA_signal_3120, key_s0[80]}), .a ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, KeyArray_outS12ser[0]}), .c ({new_AGEMA_signal_3125, new_AGEMA_signal_3124, KeyArray_inS11ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS11ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3127, new_AGEMA_signal_3126, key_s0[81]}), .a ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, KeyArray_outS12ser[1]}), .c ({new_AGEMA_signal_3131, new_AGEMA_signal_3130, KeyArray_inS11ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS11ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3133, new_AGEMA_signal_3132, key_s0[82]}), .a ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, KeyArray_outS12ser[2]}), .c ({new_AGEMA_signal_3137, new_AGEMA_signal_3136, KeyArray_inS11ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS11ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3139, new_AGEMA_signal_3138, key_s0[83]}), .a ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, KeyArray_outS12ser[3]}), .c ({new_AGEMA_signal_3143, new_AGEMA_signal_3142, KeyArray_inS11ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS11ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3145, new_AGEMA_signal_3144, key_s0[84]}), .a ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, KeyArray_outS12ser[4]}), .c ({new_AGEMA_signal_3149, new_AGEMA_signal_3148, KeyArray_inS11ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS11ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3151, new_AGEMA_signal_3150, key_s0[85]}), .a ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, KeyArray_outS12ser[5]}), .c ({new_AGEMA_signal_3155, new_AGEMA_signal_3154, KeyArray_inS11ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS11ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3157, new_AGEMA_signal_3156, key_s0[86]}), .a ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, KeyArray_outS12ser[6]}), .c ({new_AGEMA_signal_3161, new_AGEMA_signal_3160, KeyArray_inS11ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS11ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3071, new_AGEMA_signal_3070, KeyArray_n44}), .b ({new_AGEMA_signal_3163, new_AGEMA_signal_3162, key_s0[87]}), .a ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, KeyArray_outS12ser[7]}), .c ({new_AGEMA_signal_3167, new_AGEMA_signal_3166, KeyArray_inS11ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS12ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3171, new_AGEMA_signal_3170, key_s0[72]}), .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, keySBIn[0]}), .c ({new_AGEMA_signal_3175, new_AGEMA_signal_3174, KeyArray_inS12ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS12ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3177, new_AGEMA_signal_3176, key_s0[73]}), .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, keySBIn[1]}), .c ({new_AGEMA_signal_3181, new_AGEMA_signal_3180, KeyArray_inS12ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS12ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3183, new_AGEMA_signal_3182, key_s0[74]}), .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, keySBIn[2]}), .c ({new_AGEMA_signal_3187, new_AGEMA_signal_3186, KeyArray_inS12ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS12ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3189, new_AGEMA_signal_3188, key_s0[75]}), .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, keySBIn[3]}), .c ({new_AGEMA_signal_3193, new_AGEMA_signal_3192, KeyArray_inS12ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS12ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3195, new_AGEMA_signal_3194, key_s0[76]}), .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, keySBIn[4]}), .c ({new_AGEMA_signal_3199, new_AGEMA_signal_3198, KeyArray_inS12ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS12ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3201, new_AGEMA_signal_3200, key_s0[77]}), .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, keySBIn[5]}), .c ({new_AGEMA_signal_3205, new_AGEMA_signal_3204, KeyArray_inS12ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS12ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3207, new_AGEMA_signal_3206, key_s0[78]}), .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, keySBIn[6]}), .c ({new_AGEMA_signal_3211, new_AGEMA_signal_3210, KeyArray_inS12ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS12ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3213, new_AGEMA_signal_3212, key_s0[79]}), .a ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, keySBIn[7]}), .c ({new_AGEMA_signal_3217, new_AGEMA_signal_3216, KeyArray_inS12ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS13ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3219, new_AGEMA_signal_3218, key_s0[64]}), .a ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, KeyArray_outS20ser[0]}), .c ({new_AGEMA_signal_3223, new_AGEMA_signal_3222, KeyArray_inS13ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS13ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3225, new_AGEMA_signal_3224, key_s0[65]}), .a ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, KeyArray_outS20ser[1]}), .c ({new_AGEMA_signal_3229, new_AGEMA_signal_3228, KeyArray_inS13ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS13ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3231, new_AGEMA_signal_3230, key_s0[66]}), .a ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, KeyArray_outS20ser[2]}), .c ({new_AGEMA_signal_3235, new_AGEMA_signal_3234, KeyArray_inS13ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS13ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3237, new_AGEMA_signal_3236, key_s0[67]}), .a ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, KeyArray_outS20ser[3]}), .c ({new_AGEMA_signal_3241, new_AGEMA_signal_3240, KeyArray_inS13ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS13ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3243, new_AGEMA_signal_3242, key_s0[68]}), .a ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, KeyArray_outS20ser[4]}), .c ({new_AGEMA_signal_3247, new_AGEMA_signal_3246, KeyArray_inS13ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS13ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3249, new_AGEMA_signal_3248, key_s0[69]}), .a ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, KeyArray_outS20ser[5]}), .c ({new_AGEMA_signal_3253, new_AGEMA_signal_3252, KeyArray_inS13ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS13ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3255, new_AGEMA_signal_3254, key_s0[70]}), .a ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, KeyArray_outS20ser[6]}), .c ({new_AGEMA_signal_3259, new_AGEMA_signal_3258, KeyArray_inS13ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS13ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3169, new_AGEMA_signal_3168, KeyArray_n43}), .b ({new_AGEMA_signal_3261, new_AGEMA_signal_3260, key_s0[71]}), .a ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, KeyArray_outS20ser[7]}), .c ({new_AGEMA_signal_3265, new_AGEMA_signal_3264, KeyArray_inS13ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS20ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3269, new_AGEMA_signal_3268, key_s0[56]}), .a ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, KeyArray_outS21ser[0]}), .c ({new_AGEMA_signal_3273, new_AGEMA_signal_3272, KeyArray_inS20ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS20ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3275, new_AGEMA_signal_3274, key_s0[57]}), .a ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, KeyArray_outS21ser[1]}), .c ({new_AGEMA_signal_3279, new_AGEMA_signal_3278, KeyArray_inS20ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS20ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3281, new_AGEMA_signal_3280, key_s0[58]}), .a ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, KeyArray_outS21ser[2]}), .c ({new_AGEMA_signal_3285, new_AGEMA_signal_3284, KeyArray_inS20ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS20ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3287, new_AGEMA_signal_3286, key_s0[59]}), .a ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, KeyArray_outS21ser[3]}), .c ({new_AGEMA_signal_3291, new_AGEMA_signal_3290, KeyArray_inS20ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS20ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3293, new_AGEMA_signal_3292, key_s0[60]}), .a ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, KeyArray_outS21ser[4]}), .c ({new_AGEMA_signal_3297, new_AGEMA_signal_3296, KeyArray_inS20ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS20ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3299, new_AGEMA_signal_3298, key_s0[61]}), .a ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, KeyArray_outS21ser[5]}), .c ({new_AGEMA_signal_3303, new_AGEMA_signal_3302, KeyArray_inS20ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS20ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3305, new_AGEMA_signal_3304, key_s0[62]}), .a ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, KeyArray_outS21ser[6]}), .c ({new_AGEMA_signal_3309, new_AGEMA_signal_3308, KeyArray_inS20ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS20ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3311, new_AGEMA_signal_3310, key_s0[63]}), .a ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, KeyArray_outS21ser[7]}), .c ({new_AGEMA_signal_3315, new_AGEMA_signal_3314, KeyArray_inS20ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS21ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3317, new_AGEMA_signal_3316, key_s0[48]}), .a ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, KeyArray_outS22ser[0]}), .c ({new_AGEMA_signal_3321, new_AGEMA_signal_3320, KeyArray_inS21ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS21ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3323, new_AGEMA_signal_3322, key_s0[49]}), .a ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, KeyArray_outS22ser[1]}), .c ({new_AGEMA_signal_3327, new_AGEMA_signal_3326, KeyArray_inS21ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS21ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3329, new_AGEMA_signal_3328, key_s0[50]}), .a ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, KeyArray_outS22ser[2]}), .c ({new_AGEMA_signal_3333, new_AGEMA_signal_3332, KeyArray_inS21ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS21ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3335, new_AGEMA_signal_3334, key_s0[51]}), .a ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, KeyArray_outS22ser[3]}), .c ({new_AGEMA_signal_3339, new_AGEMA_signal_3338, KeyArray_inS21ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS21ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3341, new_AGEMA_signal_3340, key_s0[52]}), .a ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, KeyArray_outS22ser[4]}), .c ({new_AGEMA_signal_3345, new_AGEMA_signal_3344, KeyArray_inS21ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS21ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3347, new_AGEMA_signal_3346, key_s0[53]}), .a ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, KeyArray_outS22ser[5]}), .c ({new_AGEMA_signal_3351, new_AGEMA_signal_3350, KeyArray_inS21ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS21ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3353, new_AGEMA_signal_3352, key_s0[54]}), .a ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, KeyArray_outS22ser[6]}), .c ({new_AGEMA_signal_3357, new_AGEMA_signal_3356, KeyArray_inS21ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS21ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3267, new_AGEMA_signal_3266, KeyArray_n42}), .b ({new_AGEMA_signal_3359, new_AGEMA_signal_3358, key_s0[55]}), .a ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, KeyArray_outS22ser[7]}), .c ({new_AGEMA_signal_3363, new_AGEMA_signal_3362, KeyArray_inS21ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS22ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3367, new_AGEMA_signal_3366, key_s0[40]}), .a ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, KeyArray_outS23ser[0]}), .c ({new_AGEMA_signal_3371, new_AGEMA_signal_3370, KeyArray_inS22ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS22ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3373, new_AGEMA_signal_3372, key_s0[41]}), .a ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, KeyArray_outS23ser[1]}), .c ({new_AGEMA_signal_3377, new_AGEMA_signal_3376, KeyArray_inS22ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS22ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3379, new_AGEMA_signal_3378, key_s0[42]}), .a ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, KeyArray_outS23ser[2]}), .c ({new_AGEMA_signal_3383, new_AGEMA_signal_3382, KeyArray_inS22ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS22ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3385, new_AGEMA_signal_3384, key_s0[43]}), .a ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, KeyArray_outS23ser[3]}), .c ({new_AGEMA_signal_3389, new_AGEMA_signal_3388, KeyArray_inS22ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS22ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3391, new_AGEMA_signal_3390, key_s0[44]}), .a ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, KeyArray_outS23ser[4]}), .c ({new_AGEMA_signal_3395, new_AGEMA_signal_3394, KeyArray_inS22ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS22ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3397, new_AGEMA_signal_3396, key_s0[45]}), .a ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, KeyArray_outS23ser[5]}), .c ({new_AGEMA_signal_3401, new_AGEMA_signal_3400, KeyArray_inS22ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS22ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3403, new_AGEMA_signal_3402, key_s0[46]}), .a ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, KeyArray_outS23ser[6]}), .c ({new_AGEMA_signal_3407, new_AGEMA_signal_3406, KeyArray_inS22ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS22ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3409, new_AGEMA_signal_3408, key_s0[47]}), .a ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, KeyArray_outS23ser[7]}), .c ({new_AGEMA_signal_3413, new_AGEMA_signal_3412, KeyArray_inS22ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS23ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3415, new_AGEMA_signal_3414, key_s0[32]}), .a ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, KeyArray_outS30ser[0]}), .c ({new_AGEMA_signal_3419, new_AGEMA_signal_3418, KeyArray_inS23ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS23ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3421, new_AGEMA_signal_3420, key_s0[33]}), .a ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, KeyArray_outS30ser[1]}), .c ({new_AGEMA_signal_3425, new_AGEMA_signal_3424, KeyArray_inS23ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS23ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3427, new_AGEMA_signal_3426, key_s0[34]}), .a ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, KeyArray_outS30ser[2]}), .c ({new_AGEMA_signal_3431, new_AGEMA_signal_3430, KeyArray_inS23ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS23ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3433, new_AGEMA_signal_3432, key_s0[35]}), .a ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, KeyArray_outS30ser[3]}), .c ({new_AGEMA_signal_3437, new_AGEMA_signal_3436, KeyArray_inS23ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS23ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3439, new_AGEMA_signal_3438, key_s0[36]}), .a ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, KeyArray_outS30ser[4]}), .c ({new_AGEMA_signal_3443, new_AGEMA_signal_3442, KeyArray_inS23ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS23ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3445, new_AGEMA_signal_3444, key_s0[37]}), .a ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, KeyArray_outS30ser[5]}), .c ({new_AGEMA_signal_3449, new_AGEMA_signal_3448, KeyArray_inS23ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS23ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3451, new_AGEMA_signal_3450, key_s0[38]}), .a ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, KeyArray_outS30ser[6]}), .c ({new_AGEMA_signal_3455, new_AGEMA_signal_3454, KeyArray_inS23ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS23ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3365, new_AGEMA_signal_3364, KeyArray_n41}), .b ({new_AGEMA_signal_3457, new_AGEMA_signal_3456, key_s0[39]}), .a ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, KeyArray_outS30ser[7]}), .c ({new_AGEMA_signal_3461, new_AGEMA_signal_3460, KeyArray_inS23ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS30ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3465, new_AGEMA_signal_3464, key_s0[24]}), .a ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, KeyArray_outS31ser[0]}), .c ({new_AGEMA_signal_3469, new_AGEMA_signal_3468, KeyArray_inS30ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS30ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3471, new_AGEMA_signal_3470, key_s0[25]}), .a ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, KeyArray_outS31ser[1]}), .c ({new_AGEMA_signal_3475, new_AGEMA_signal_3474, KeyArray_inS30ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS30ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3477, new_AGEMA_signal_3476, key_s0[26]}), .a ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, KeyArray_outS31ser[2]}), .c ({new_AGEMA_signal_3481, new_AGEMA_signal_3480, KeyArray_inS30ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS30ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3483, new_AGEMA_signal_3482, key_s0[27]}), .a ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, KeyArray_outS31ser[3]}), .c ({new_AGEMA_signal_3487, new_AGEMA_signal_3486, KeyArray_inS30ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS30ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3489, new_AGEMA_signal_3488, key_s0[28]}), .a ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, KeyArray_outS31ser[4]}), .c ({new_AGEMA_signal_3493, new_AGEMA_signal_3492, KeyArray_inS30ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS30ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3495, new_AGEMA_signal_3494, key_s0[29]}), .a ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, KeyArray_outS31ser[5]}), .c ({new_AGEMA_signal_3499, new_AGEMA_signal_3498, KeyArray_inS30ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS30ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3501, new_AGEMA_signal_3500, key_s0[30]}), .a ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, KeyArray_outS31ser[6]}), .c ({new_AGEMA_signal_3505, new_AGEMA_signal_3504, KeyArray_inS30ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS30ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3507, new_AGEMA_signal_3506, key_s0[31]}), .a ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, KeyArray_outS31ser[7]}), .c ({new_AGEMA_signal_3511, new_AGEMA_signal_3510, KeyArray_inS30ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS31ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3513, new_AGEMA_signal_3512, key_s0[16]}), .a ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, KeyArray_outS32ser[0]}), .c ({new_AGEMA_signal_3517, new_AGEMA_signal_3516, KeyArray_inS31ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS31ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3519, new_AGEMA_signal_3518, key_s0[17]}), .a ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, KeyArray_outS32ser[1]}), .c ({new_AGEMA_signal_3523, new_AGEMA_signal_3522, KeyArray_inS31ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS31ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3525, new_AGEMA_signal_3524, key_s0[18]}), .a ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, KeyArray_outS32ser[2]}), .c ({new_AGEMA_signal_3529, new_AGEMA_signal_3528, KeyArray_inS31ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS31ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3531, new_AGEMA_signal_3530, key_s0[19]}), .a ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, KeyArray_outS32ser[3]}), .c ({new_AGEMA_signal_3535, new_AGEMA_signal_3534, KeyArray_inS31ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS31ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3537, new_AGEMA_signal_3536, key_s0[20]}), .a ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, KeyArray_outS32ser[4]}), .c ({new_AGEMA_signal_3541, new_AGEMA_signal_3540, KeyArray_inS31ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS31ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3543, new_AGEMA_signal_3542, key_s0[21]}), .a ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, KeyArray_outS32ser[5]}), .c ({new_AGEMA_signal_3547, new_AGEMA_signal_3546, KeyArray_inS31ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS31ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3549, new_AGEMA_signal_3548, key_s0[22]}), .a ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, KeyArray_outS32ser[6]}), .c ({new_AGEMA_signal_3553, new_AGEMA_signal_3552, KeyArray_inS31ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS31ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3463, new_AGEMA_signal_3462, KeyArray_n40}), .b ({new_AGEMA_signal_3555, new_AGEMA_signal_3554, key_s0[23]}), .a ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, KeyArray_outS32ser[7]}), .c ({new_AGEMA_signal_3559, new_AGEMA_signal_3558, KeyArray_inS31ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS32ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3563, new_AGEMA_signal_3562, key_s0[8]}), .a ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, KeyArray_outS33ser[0]}), .c ({new_AGEMA_signal_3567, new_AGEMA_signal_3566, KeyArray_inS32ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS32ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3569, new_AGEMA_signal_3568, key_s0[9]}), .a ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, KeyArray_outS33ser[1]}), .c ({new_AGEMA_signal_3573, new_AGEMA_signal_3572, KeyArray_inS32ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS32ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3575, new_AGEMA_signal_3574, key_s0[10]}), .a ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, KeyArray_outS33ser[2]}), .c ({new_AGEMA_signal_3579, new_AGEMA_signal_3578, KeyArray_inS32ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS32ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3581, new_AGEMA_signal_3580, key_s0[11]}), .a ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, KeyArray_outS33ser[3]}), .c ({new_AGEMA_signal_3585, new_AGEMA_signal_3584, KeyArray_inS32ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS32ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3587, new_AGEMA_signal_3586, key_s0[12]}), .a ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, KeyArray_outS33ser[4]}), .c ({new_AGEMA_signal_3591, new_AGEMA_signal_3590, KeyArray_inS32ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS32ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3593, new_AGEMA_signal_3592, key_s0[13]}), .a ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, KeyArray_outS33ser[5]}), .c ({new_AGEMA_signal_3597, new_AGEMA_signal_3596, KeyArray_inS32ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS32ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3599, new_AGEMA_signal_3598, key_s0[14]}), .a ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, KeyArray_outS33ser[6]}), .c ({new_AGEMA_signal_3603, new_AGEMA_signal_3602, KeyArray_inS32ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS32ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3605, new_AGEMA_signal_3604, key_s0[15]}), .a ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, KeyArray_outS33ser[7]}), .c ({new_AGEMA_signal_3609, new_AGEMA_signal_3608, KeyArray_inS32ser[7]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS33ser_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3611, new_AGEMA_signal_3610, key_s0[0]}), .a ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, keyStateIn[0]}), .c ({new_AGEMA_signal_3613, new_AGEMA_signal_3612, KeyArray_inS33ser[0]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS33ser_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3615, new_AGEMA_signal_3614, key_s0[1]}), .a ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}), .c ({new_AGEMA_signal_3617, new_AGEMA_signal_3616, KeyArray_inS33ser[1]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS33ser_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3619, new_AGEMA_signal_3618, key_s0[2]}), .a ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, keyStateIn[2]}), .c ({new_AGEMA_signal_3621, new_AGEMA_signal_3620, KeyArray_inS33ser[2]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS33ser_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3623, new_AGEMA_signal_3622, key_s0[3]}), .a ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, keyStateIn[3]}), .c ({new_AGEMA_signal_3625, new_AGEMA_signal_3624, KeyArray_inS33ser[3]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS33ser_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3627, new_AGEMA_signal_3626, key_s0[4]}), .a ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[4]}), .c ({new_AGEMA_signal_3629, new_AGEMA_signal_3628, KeyArray_inS33ser[4]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS33ser_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3631, new_AGEMA_signal_3630, key_s0[5]}), .a ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, keyStateIn[5]}), .c ({new_AGEMA_signal_3633, new_AGEMA_signal_3632, KeyArray_inS33ser[5]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS33ser_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3635, new_AGEMA_signal_3634, key_s0[6]}), .a ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, keyStateIn[6]}), .c ({new_AGEMA_signal_3637, new_AGEMA_signal_3636, KeyArray_inS33ser[6]}) ) ;
    mux2_masked_LMDPL KeyArray_MUX_inS33ser_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3561, new_AGEMA_signal_3560, KeyArray_n39}), .b ({new_AGEMA_signal_3639, new_AGEMA_signal_3638, key_s0[7]}), .a ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[7]}), .c ({new_AGEMA_signal_3641, new_AGEMA_signal_3640, KeyArray_inS33ser[7]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U24 ( .a ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, MixColumns_line0_n16}), .b ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, MixColumns_line0_n15}), .c ({new_AGEMA_signal_3643, new_AGEMA_signal_3642, MCout[31]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U23 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2071, new_AGEMA_signal_2070, MixColumns_line0_n15}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_U22 ( .a ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, MixColumns_line0_S13[7]}), .c ({new_AGEMA_signal_2267, new_AGEMA_signal_2266, MixColumns_line0_n16}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U21 ( .a ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, MixColumns_line0_n14}), .b ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, MixColumns_line0_n13}), .c ({new_AGEMA_signal_3645, new_AGEMA_signal_3644, MCout[30]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U20 ( .a ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2077, new_AGEMA_signal_2076, MixColumns_line0_n13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_U19 ( .a ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, MixColumns_line0_S13[6]}), .c ({new_AGEMA_signal_2269, new_AGEMA_signal_2268, MixColumns_line0_n14}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U18 ( .a ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, MixColumns_line0_n12}), .b ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, MixColumns_line0_n11}), .c ({new_AGEMA_signal_3647, new_AGEMA_signal_3646, MCout[29]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U17 ( .a ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2083, new_AGEMA_signal_2082, MixColumns_line0_n11}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_U16 ( .a ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, MixColumns_line0_S13[5]}), .c ({new_AGEMA_signal_2271, new_AGEMA_signal_2270, MixColumns_line0_n12}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U15 ( .a ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, MixColumns_line0_n10}), .b ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, MixColumns_line0_n9}), .c ({new_AGEMA_signal_3735, new_AGEMA_signal_3734, MCout[28]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U14 ( .a ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2089, new_AGEMA_signal_2088, MixColumns_line0_n9}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_U13 ( .a ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, MixColumns_line0_S02[4]}), .b ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, MixColumns_line0_S13[4]}), .c ({new_AGEMA_signal_3649, new_AGEMA_signal_3648, MixColumns_line0_n10}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U12 ( .a ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, MixColumns_line0_n8}), .b ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, MixColumns_line0_n7}), .c ({new_AGEMA_signal_3737, new_AGEMA_signal_3736, MCout[27]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U11 ( .a ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2095, new_AGEMA_signal_2094, MixColumns_line0_n7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_U10 ( .a ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, MixColumns_line0_S02[3]}), .b ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, MixColumns_line0_S13[3]}), .c ({new_AGEMA_signal_3651, new_AGEMA_signal_3650, MixColumns_line0_n8}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U9 ( .a ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, MixColumns_line0_n6}), .b ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, MixColumns_line0_n5}), .c ({new_AGEMA_signal_3653, new_AGEMA_signal_3652, MCout[26]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U8 ( .a ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2101, new_AGEMA_signal_2100, MixColumns_line0_n5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_U7 ( .a ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, MixColumns_line0_S13[2]}), .c ({new_AGEMA_signal_2273, new_AGEMA_signal_2272, MixColumns_line0_n6}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U6 ( .a ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, MixColumns_line0_n4}), .b ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, MixColumns_line0_n3}), .c ({new_AGEMA_signal_3739, new_AGEMA_signal_3738, MCout[25]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U5 ( .a ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2107, new_AGEMA_signal_2106, MixColumns_line0_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_U4 ( .a ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, MixColumns_line0_S02[1]}), .b ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, MixColumns_line0_S13[1]}), .c ({new_AGEMA_signal_3655, new_AGEMA_signal_3654, MixColumns_line0_n4}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U3 ( .a ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, MixColumns_line0_n2}), .b ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, MixColumns_line0_n1}), .c ({new_AGEMA_signal_3657, new_AGEMA_signal_3656, MCout[24]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line0_U2 ( .a ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2113, new_AGEMA_signal_2112, MixColumns_line0_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_U1 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, MixColumns_line0_S13[0]}), .c ({new_AGEMA_signal_2275, new_AGEMA_signal_2274, MixColumns_line0_n2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTWO_U3 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2115, new_AGEMA_signal_2114, MixColumns_line0_S02[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTWO_U2 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2117, new_AGEMA_signal_2116, MixColumns_line0_S02[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTWO_U1 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2119, new_AGEMA_signal_2118, MixColumns_line0_S02[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_U8 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2125, new_AGEMA_signal_2124, MixColumns_line0_S13[7]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_U7 ( .a ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2129, new_AGEMA_signal_2128, MixColumns_line0_S13[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_U6 ( .a ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2133, new_AGEMA_signal_2132, MixColumns_line0_S13[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_U5 ( .a ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, MixColumns_line0_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2277, new_AGEMA_signal_2276, MixColumns_line0_S13[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_U4 ( .a ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, MixColumns_line0_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2279, new_AGEMA_signal_2278, MixColumns_line0_S13[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_U3 ( .a ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}), .b ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2139, new_AGEMA_signal_2138, MixColumns_line0_S13[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_U2 ( .a ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, MixColumns_line0_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2281, new_AGEMA_signal_2280, MixColumns_line0_S13[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_U1 ( .a ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2143, new_AGEMA_signal_2142, MixColumns_line0_S13[0]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U3 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2147, new_AGEMA_signal_2146, MixColumns_line0_timesTHREE_input2[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U2 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2149, new_AGEMA_signal_2148, MixColumns_line0_timesTHREE_input2[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line0_timesTHREE_timesTWO_U1 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2151, new_AGEMA_signal_2150, MixColumns_line0_timesTHREE_input2[1]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U24 ( .a ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, MixColumns_line1_n16}), .b ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, MixColumns_line1_n15}), .c ({new_AGEMA_signal_3659, new_AGEMA_signal_3658, MCout[23]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U23 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2153, new_AGEMA_signal_2152, MixColumns_line1_n15}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_U22 ( .a ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, MixColumns_line1_S13[7]}), .c ({new_AGEMA_signal_2283, new_AGEMA_signal_2282, MixColumns_line1_n16}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U21 ( .a ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, MixColumns_line1_n14}), .b ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, MixColumns_line1_n13}), .c ({new_AGEMA_signal_3661, new_AGEMA_signal_3660, MCout[22]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U20 ( .a ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2155, new_AGEMA_signal_2154, MixColumns_line1_n13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_U19 ( .a ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, MixColumns_line1_S13[6]}), .c ({new_AGEMA_signal_2285, new_AGEMA_signal_2284, MixColumns_line1_n14}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U18 ( .a ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, MixColumns_line1_n12}), .b ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, MixColumns_line1_n11}), .c ({new_AGEMA_signal_3663, new_AGEMA_signal_3662, MCout[21]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U17 ( .a ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2157, new_AGEMA_signal_2156, MixColumns_line1_n11}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_U16 ( .a ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, MixColumns_line1_S13[5]}), .c ({new_AGEMA_signal_2287, new_AGEMA_signal_2286, MixColumns_line1_n12}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U15 ( .a ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, MixColumns_line1_n10}), .b ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, MixColumns_line1_n9}), .c ({new_AGEMA_signal_3741, new_AGEMA_signal_3740, MCout[20]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U14 ( .a ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2159, new_AGEMA_signal_2158, MixColumns_line1_n9}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_U13 ( .a ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, MixColumns_line1_S02_4_}), .b ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, MixColumns_line1_S13[4]}), .c ({new_AGEMA_signal_3665, new_AGEMA_signal_3664, MixColumns_line1_n10}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U12 ( .a ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, MixColumns_line1_n8}), .b ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, MixColumns_line1_n7}), .c ({new_AGEMA_signal_3743, new_AGEMA_signal_3742, MCout[19]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U11 ( .a ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2161, new_AGEMA_signal_2160, MixColumns_line1_n7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_U10 ( .a ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, MixColumns_line1_S02_3_}), .b ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, MixColumns_line1_S13[3]}), .c ({new_AGEMA_signal_3667, new_AGEMA_signal_3666, MixColumns_line1_n8}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U9 ( .a ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, MixColumns_line1_n6}), .b ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, MixColumns_line1_n5}), .c ({new_AGEMA_signal_3669, new_AGEMA_signal_3668, MCout[18]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U8 ( .a ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2163, new_AGEMA_signal_2162, MixColumns_line1_n5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_U7 ( .a ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, MixColumns_line1_S13[2]}), .c ({new_AGEMA_signal_2289, new_AGEMA_signal_2288, MixColumns_line1_n6}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U6 ( .a ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, MixColumns_line1_n4}), .b ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, MixColumns_line1_n3}), .c ({new_AGEMA_signal_3745, new_AGEMA_signal_3744, MCout[17]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U5 ( .a ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2165, new_AGEMA_signal_2164, MixColumns_line1_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_U4 ( .a ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, MixColumns_line1_S02_1_}), .b ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, MixColumns_line1_S13[1]}), .c ({new_AGEMA_signal_3671, new_AGEMA_signal_3670, MixColumns_line1_n4}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U3 ( .a ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, MixColumns_line1_n2}), .b ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, MixColumns_line1_n1}), .c ({new_AGEMA_signal_3673, new_AGEMA_signal_3672, MCout[16]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line1_U2 ( .a ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2167, new_AGEMA_signal_2166, MixColumns_line1_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_U1 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, MixColumns_line1_S13[0]}), .c ({new_AGEMA_signal_2291, new_AGEMA_signal_2290, MixColumns_line1_n2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTWO_U3 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2169, new_AGEMA_signal_2168, MixColumns_line1_S02_4_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTWO_U2 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2171, new_AGEMA_signal_2170, MixColumns_line1_S02_3_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTWO_U1 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2173, new_AGEMA_signal_2172, MixColumns_line1_S02_1_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_U8 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2175, new_AGEMA_signal_2174, MixColumns_line1_S13[7]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_U7 ( .a ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2177, new_AGEMA_signal_2176, MixColumns_line1_S13[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_U6 ( .a ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2179, new_AGEMA_signal_2178, MixColumns_line1_S13[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_U5 ( .a ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, MixColumns_line1_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2293, new_AGEMA_signal_2292, MixColumns_line1_S13[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_U4 ( .a ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}), .b ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, MixColumns_line1_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2295, new_AGEMA_signal_2294, MixColumns_line1_S13[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_U3 ( .a ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}), .b ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}), .c ({new_AGEMA_signal_2181, new_AGEMA_signal_2180, MixColumns_line1_S13[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_U2 ( .a ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, MixColumns_line1_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2297, new_AGEMA_signal_2296, MixColumns_line1_S13[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_U1 ( .a ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2183, new_AGEMA_signal_2182, MixColumns_line1_S13[0]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U3 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2185, new_AGEMA_signal_2184, MixColumns_line1_timesTHREE_input2[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U2 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2187, new_AGEMA_signal_2186, MixColumns_line1_timesTHREE_input2[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line1_timesTHREE_timesTWO_U1 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2189, new_AGEMA_signal_2188, MixColumns_line1_timesTHREE_input2[1]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U24 ( .a ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, MixColumns_line2_n16}), .b ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, MixColumns_line2_n15}), .c ({new_AGEMA_signal_3675, new_AGEMA_signal_3674, MCout[15]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U23 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .c ({new_AGEMA_signal_2191, new_AGEMA_signal_2190, MixColumns_line2_n15}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_U22 ( .a ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}), .b ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, MixColumns_line2_S13[7]}), .c ({new_AGEMA_signal_2299, new_AGEMA_signal_2298, MixColumns_line2_n16}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U21 ( .a ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, MixColumns_line2_n14}), .b ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, MixColumns_line2_n13}), .c ({new_AGEMA_signal_3677, new_AGEMA_signal_3676, MCout[14]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U20 ( .a ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}), .c ({new_AGEMA_signal_2193, new_AGEMA_signal_2192, MixColumns_line2_n13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_U19 ( .a ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}), .b ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, MixColumns_line2_S13[6]}), .c ({new_AGEMA_signal_2301, new_AGEMA_signal_2300, MixColumns_line2_n14}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U18 ( .a ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, MixColumns_line2_n12}), .b ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, MixColumns_line2_n11}), .c ({new_AGEMA_signal_3679, new_AGEMA_signal_3678, MCout[13]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U17 ( .a ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}), .c ({new_AGEMA_signal_2195, new_AGEMA_signal_2194, MixColumns_line2_n11}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_U16 ( .a ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}), .b ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, MixColumns_line2_S13[5]}), .c ({new_AGEMA_signal_2303, new_AGEMA_signal_2302, MixColumns_line2_n12}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U15 ( .a ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, MixColumns_line2_n10}), .b ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, MixColumns_line2_n9}), .c ({new_AGEMA_signal_3747, new_AGEMA_signal_3746, MCout[12]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U14 ( .a ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}), .c ({new_AGEMA_signal_2197, new_AGEMA_signal_2196, MixColumns_line2_n9}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_U13 ( .a ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, MixColumns_line2_S02_4_}), .b ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, MixColumns_line2_S13[4]}), .c ({new_AGEMA_signal_3681, new_AGEMA_signal_3680, MixColumns_line2_n10}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U12 ( .a ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, MixColumns_line2_n8}), .b ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, MixColumns_line2_n7}), .c ({new_AGEMA_signal_3749, new_AGEMA_signal_3748, MCout[11]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U11 ( .a ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}), .c ({new_AGEMA_signal_2199, new_AGEMA_signal_2198, MixColumns_line2_n7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_U10 ( .a ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, MixColumns_line2_S02_3_}), .b ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, MixColumns_line2_S13[3]}), .c ({new_AGEMA_signal_3683, new_AGEMA_signal_3682, MixColumns_line2_n8}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U9 ( .a ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, MixColumns_line2_n6}), .b ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, MixColumns_line2_n5}), .c ({new_AGEMA_signal_3685, new_AGEMA_signal_3684, MCout[10]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U8 ( .a ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}), .c ({new_AGEMA_signal_2201, new_AGEMA_signal_2200, MixColumns_line2_n5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_U7 ( .a ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, MixColumns_line2_S13[2]}), .c ({new_AGEMA_signal_2305, new_AGEMA_signal_2304, MixColumns_line2_n6}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U6 ( .a ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, MixColumns_line2_n4}), .b ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, MixColumns_line2_n3}), .c ({new_AGEMA_signal_3751, new_AGEMA_signal_3750, MCout[9]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U5 ( .a ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}), .b ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2203, new_AGEMA_signal_2202, MixColumns_line2_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_U4 ( .a ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, MixColumns_line2_S02_1_}), .b ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, MixColumns_line2_S13[1]}), .c ({new_AGEMA_signal_3687, new_AGEMA_signal_3686, MixColumns_line2_n4}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U3 ( .a ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, MixColumns_line2_n2}), .b ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, MixColumns_line2_n1}), .c ({new_AGEMA_signal_3689, new_AGEMA_signal_3688, MCout[8]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line2_U2 ( .a ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}), .b ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2205, new_AGEMA_signal_2204, MixColumns_line2_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_U1 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, MixColumns_line2_S13[0]}), .c ({new_AGEMA_signal_2307, new_AGEMA_signal_2306, MixColumns_line2_n2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTWO_U3 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2207, new_AGEMA_signal_2206, MixColumns_line2_S02_4_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTWO_U2 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2209, new_AGEMA_signal_2208, MixColumns_line2_S02_3_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTWO_U1 ( .a ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .b ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}), .c ({new_AGEMA_signal_2211, new_AGEMA_signal_2210, MixColumns_line2_S02_1_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_U8 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}), .c ({new_AGEMA_signal_2213, new_AGEMA_signal_2212, MixColumns_line2_S13[7]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_U7 ( .a ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}), .c ({new_AGEMA_signal_2215, new_AGEMA_signal_2214, MixColumns_line2_S13[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_U6 ( .a ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}), .c ({new_AGEMA_signal_2217, new_AGEMA_signal_2216, MixColumns_line2_S13[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_U5 ( .a ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, MixColumns_line2_timesTHREE_input2[4]}), .c ({new_AGEMA_signal_2309, new_AGEMA_signal_2308, MixColumns_line2_S13[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_U4 ( .a ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}), .b ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, MixColumns_line2_timesTHREE_input2[3]}), .c ({new_AGEMA_signal_2311, new_AGEMA_signal_2310, MixColumns_line2_S13[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_U3 ( .a ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}), .b ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}), .c ({new_AGEMA_signal_2219, new_AGEMA_signal_2218, MixColumns_line2_S13[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_U2 ( .a ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, MixColumns_line2_timesTHREE_input2[1]}), .c ({new_AGEMA_signal_2313, new_AGEMA_signal_2312, MixColumns_line2_S13[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_U1 ( .a ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}), .b ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .c ({new_AGEMA_signal_2221, new_AGEMA_signal_2220, MixColumns_line2_S13[0]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U3 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2223, new_AGEMA_signal_2222, MixColumns_line2_timesTHREE_input2[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U2 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2225, new_AGEMA_signal_2224, MixColumns_line2_timesTHREE_input2[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line2_timesTHREE_timesTWO_U1 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2227, new_AGEMA_signal_2226, MixColumns_line2_timesTHREE_input2[1]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U24 ( .a ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, MixColumns_line3_n16}), .b ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, MixColumns_line3_n15}), .c ({new_AGEMA_signal_3691, new_AGEMA_signal_3690, MCout[7]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U23 ( .a ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}), .b ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}), .c ({new_AGEMA_signal_2229, new_AGEMA_signal_2228, MixColumns_line3_n15}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_U22 ( .a ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}), .b ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, MixColumns_line3_S13[7]}), .c ({new_AGEMA_signal_2315, new_AGEMA_signal_2314, MixColumns_line3_n16}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U21 ( .a ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, MixColumns_line3_n14}), .b ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, MixColumns_line3_n13}), .c ({new_AGEMA_signal_3693, new_AGEMA_signal_3692, MCout[6]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U20 ( .a ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}), .b ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}), .c ({new_AGEMA_signal_2231, new_AGEMA_signal_2230, MixColumns_line3_n13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_U19 ( .a ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}), .b ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, MixColumns_line3_S13[6]}), .c ({new_AGEMA_signal_2317, new_AGEMA_signal_2316, MixColumns_line3_n14}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U18 ( .a ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, MixColumns_line3_n12}), .b ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, MixColumns_line3_n11}), .c ({new_AGEMA_signal_3695, new_AGEMA_signal_3694, MCout[5]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U17 ( .a ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}), .b ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}), .c ({new_AGEMA_signal_2233, new_AGEMA_signal_2232, MixColumns_line3_n11}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_U16 ( .a ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}), .b ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, MixColumns_line3_S13[5]}), .c ({new_AGEMA_signal_2319, new_AGEMA_signal_2318, MixColumns_line3_n12}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U15 ( .a ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, MixColumns_line3_n10}), .b ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, MixColumns_line3_n9}), .c ({new_AGEMA_signal_3753, new_AGEMA_signal_3752, MCout[4]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U14 ( .a ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}), .b ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}), .c ({new_AGEMA_signal_2235, new_AGEMA_signal_2234, MixColumns_line3_n9}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_U13 ( .a ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, MixColumns_line3_S02_4_}), .b ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, MixColumns_line3_S13[4]}), .c ({new_AGEMA_signal_3697, new_AGEMA_signal_3696, MixColumns_line3_n10}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U12 ( .a ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, MixColumns_line3_n8}), .b ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, MixColumns_line3_n7}), .c ({new_AGEMA_signal_3755, new_AGEMA_signal_3754, MCout[3]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U11 ( .a ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}), .b ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}), .c ({new_AGEMA_signal_2237, new_AGEMA_signal_2236, MixColumns_line3_n7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_U10 ( .a ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, MixColumns_line3_S02_3_}), .b ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, MixColumns_line3_S13[3]}), .c ({new_AGEMA_signal_3699, new_AGEMA_signal_3698, MixColumns_line3_n8}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U9 ( .a ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, MixColumns_line3_n6}), .b ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, MixColumns_line3_n5}), .c ({new_AGEMA_signal_3701, new_AGEMA_signal_3700, MCout[2]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U8 ( .a ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}), .b ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}), .c ({new_AGEMA_signal_2239, new_AGEMA_signal_2238, MixColumns_line3_n5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_U7 ( .a ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}), .b ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, MixColumns_line3_S13[2]}), .c ({new_AGEMA_signal_2321, new_AGEMA_signal_2320, MixColumns_line3_n6}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U6 ( .a ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, MixColumns_line3_n4}), .b ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, MixColumns_line3_n3}), .c ({new_AGEMA_signal_3757, new_AGEMA_signal_3756, MCout[1]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U5 ( .a ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}), .b ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}), .c ({new_AGEMA_signal_2241, new_AGEMA_signal_2240, MixColumns_line3_n3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_U4 ( .a ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, MixColumns_line3_S02_1_}), .b ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, MixColumns_line3_S13[1]}), .c ({new_AGEMA_signal_3703, new_AGEMA_signal_3702, MixColumns_line3_n4}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U3 ( .a ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, MixColumns_line3_n2}), .b ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, MixColumns_line3_n1}), .c ({new_AGEMA_signal_3705, new_AGEMA_signal_3704, MCout[0]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) MixColumns_line3_U2 ( .a ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}), .b ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}), .c ({new_AGEMA_signal_2243, new_AGEMA_signal_2242, MixColumns_line3_n1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_U1 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, MixColumns_line3_S13[0]}), .c ({new_AGEMA_signal_2323, new_AGEMA_signal_2322, MixColumns_line3_n2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTWO_U3 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}), .c ({new_AGEMA_signal_2245, new_AGEMA_signal_2244, MixColumns_line3_S02_4_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTWO_U2 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}), .c ({new_AGEMA_signal_2247, new_AGEMA_signal_2246, MixColumns_line3_S02_3_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTWO_U1 ( .a ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}), .b ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}), .c ({new_AGEMA_signal_2249, new_AGEMA_signal_2248, MixColumns_line3_S02_1_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_U8 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}), .c ({new_AGEMA_signal_2251, new_AGEMA_signal_2250, MixColumns_line3_S13[7]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_U7 ( .a ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}), .b ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}), .c ({new_AGEMA_signal_2253, new_AGEMA_signal_2252, MixColumns_line3_S13[6]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_U6 ( .a ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}), .b ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}), .c ({new_AGEMA_signal_2255, new_AGEMA_signal_2254, MixColumns_line3_S13[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_U5 ( .a ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}), .b ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, MixColumns_line3_timesTHREE_input2_4_}), .c ({new_AGEMA_signal_2325, new_AGEMA_signal_2324, MixColumns_line3_S13[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_U4 ( .a ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}), .b ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, MixColumns_line3_timesTHREE_input2_3_}), .c ({new_AGEMA_signal_2327, new_AGEMA_signal_2326, MixColumns_line3_S13[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_U3 ( .a ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}), .b ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}), .c ({new_AGEMA_signal_2257, new_AGEMA_signal_2256, MixColumns_line3_S13[2]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_U2 ( .a ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}), .b ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, MixColumns_line3_timesTHREE_input2_1_}), .c ({new_AGEMA_signal_2329, new_AGEMA_signal_2328, MixColumns_line3_S13[1]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_U1 ( .a ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}), .b ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .c ({new_AGEMA_signal_2259, new_AGEMA_signal_2258, MixColumns_line3_S13[0]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U3 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}), .c ({new_AGEMA_signal_2261, new_AGEMA_signal_2260, MixColumns_line3_timesTHREE_input2_4_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U2 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}), .c ({new_AGEMA_signal_2263, new_AGEMA_signal_2262, MixColumns_line3_timesTHREE_input2_3_}) ) ;
    linear_LMDPL #(.CONF(1'b0)) MixColumns_line3_timesTHREE_timesTWO_U1 ( .a ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}), .b ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}), .c ({new_AGEMA_signal_2265, new_AGEMA_signal_2264, MixColumns_line3_timesTHREE_input2_1_}) ) ;
    NOR2_X1 calcRCon_U46 ( .A1 (calcRCon_n11), .A2 (calcRCon_n38), .ZN (roundConstant[7]) ) ;
    NOR2_X1 calcRCon_U45 ( .A1 (calcRCon_n16), .A2 (calcRCon_n38), .ZN (roundConstant[6]) ) ;
    AND2_X1 calcRCon_U44 ( .A1 (calcRCon_s_current_state_5_), .A2 (enRCon), .ZN (roundConstant[5]) ) ;
    AND2_X1 calcRCon_U43 ( .A1 (calcRCon_s_current_state_4_), .A2 (enRCon), .ZN (roundConstant[4]) ) ;
    NOR2_X1 calcRCon_U42 ( .A1 (calcRCon_n15), .A2 (calcRCon_n38), .ZN (roundConstant[3]) ) ;
    NOR2_X1 calcRCon_U41 ( .A1 (calcRCon_n12), .A2 (calcRCon_n38), .ZN (roundConstant[2]) ) ;
    NOR2_X1 calcRCon_U40 ( .A1 (calcRCon_n14), .A2 (calcRCon_n38), .ZN (roundConstant[1]) ) ;
    NOR2_X1 calcRCon_U39 ( .A1 (calcRCon_n13), .A2 (calcRCon_n38), .ZN (roundConstant[0]) ) ;
    INV_X1 calcRCon_U38 ( .A (enRCon), .ZN (calcRCon_n38) ) ;
    NAND2_X1 calcRCon_U37 ( .A1 (calcRCon_n37), .A2 (calcRCon_n36), .ZN (notFirst) ) ;
    NOR2_X1 calcRCon_U36 ( .A1 (calcRCon_n35), .A2 (calcRCon_n34), .ZN (calcRCon_n36) ) ;
    NAND2_X1 calcRCon_U35 ( .A1 (calcRCon_n33), .A2 (calcRCon_n32), .ZN (calcRCon_n34) ) ;
    NOR2_X1 calcRCon_U34 ( .A1 (calcRCon_s_current_state_1_), .A2 (calcRCon_n15), .ZN (calcRCon_n32) ) ;
    NOR2_X1 calcRCon_U33 ( .A1 (calcRCon_s_current_state_6_), .A2 (calcRCon_n13), .ZN (calcRCon_n33) ) ;
    NAND2_X1 calcRCon_U32 ( .A1 (calcRCon_s_current_state_2_), .A2 (calcRCon_n3), .ZN (calcRCon_n35) ) ;
    NOR2_X1 calcRCon_U31 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_s_current_state_5_), .ZN (calcRCon_n37) ) ;
    NAND2_X1 calcRCon_U30 ( .A1 (nReset), .A2 (calcRCon_n31), .ZN (calcRCon_n51) ) ;
    MUX2_X1 calcRCon_U29 ( .S (calcRCon_n5), .A (calcRCon_n11), .B (calcRCon_n13), .Z (calcRCon_n31) ) ;
    NAND2_X1 calcRCon_U28 ( .A1 (calcRCon_n30), .A2 (calcRCon_n29), .ZN (calcRCon_n50) ) ;
    NAND2_X1 calcRCon_U27 ( .A1 (calcRCon_n28), .A2 (calcRCon_s_current_state_1_), .ZN (calcRCon_n29) ) ;
    NAND2_X1 calcRCon_U26 ( .A1 (calcRCon_n27), .A2 (calcRCon_n26), .ZN (calcRCon_n30) ) ;
    XOR2_X1 calcRCon_U25 ( .A (calcRCon_s_current_state_0_), .B (calcRCon_n3), .Z (calcRCon_n27) ) ;
    NAND2_X1 calcRCon_U24 ( .A1 (nReset), .A2 (calcRCon_n25), .ZN (calcRCon_n49) ) ;
    MUX2_X1 calcRCon_U23 ( .S (calcRCon_n5), .A (calcRCon_n14), .B (calcRCon_n12), .Z (calcRCon_n25) ) ;
    NAND2_X1 calcRCon_U22 ( .A1 (nReset), .A2 (calcRCon_n24), .ZN (calcRCon_n48) ) ;
    MUX2_X1 calcRCon_U21 ( .S (calcRCon_n5), .A (calcRCon_n23), .B (calcRCon_n15), .Z (calcRCon_n24) ) ;
    XNOR2_X1 calcRCon_U20 ( .A (calcRCon_n3), .B (calcRCon_s_current_state_2_), .ZN (calcRCon_n23) ) ;
    NAND2_X1 calcRCon_U19 ( .A1 (calcRCon_n22), .A2 (calcRCon_n21), .ZN (calcRCon_n47) ) ;
    NAND2_X1 calcRCon_U18 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_n28), .ZN (calcRCon_n21) ) ;
    NAND2_X1 calcRCon_U17 ( .A1 (calcRCon_n20), .A2 (calcRCon_n26), .ZN (calcRCon_n22) ) ;
    XOR2_X1 calcRCon_U16 ( .A (calcRCon_n15), .B (calcRCon_n11), .Z (calcRCon_n20) ) ;
    NAND2_X1 calcRCon_U15 ( .A1 (calcRCon_n19), .A2 (calcRCon_n18), .ZN (calcRCon_n46) ) ;
    NAND2_X1 calcRCon_U14 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_n26), .ZN (calcRCon_n18) ) ;
    NAND2_X1 calcRCon_U13 ( .A1 (calcRCon_s_current_state_5_), .A2 (calcRCon_n28), .ZN (calcRCon_n19) ) ;
    NAND2_X1 calcRCon_U12 ( .A1 (calcRCon_n17), .A2 (calcRCon_n10), .ZN (calcRCon_n45) ) ;
    NAND2_X1 calcRCon_U11 ( .A1 (calcRCon_s_current_state_5_), .A2 (calcRCon_n26), .ZN (calcRCon_n10) ) ;
    NOR2_X1 calcRCon_U10 ( .A1 (calcRCon_n5), .A2 (calcRCon_n6), .ZN (calcRCon_n26) ) ;
    NAND2_X1 calcRCon_U9 ( .A1 (calcRCon_s_current_state_6_), .A2 (calcRCon_n28), .ZN (calcRCon_n17) ) ;
    NOR2_X1 calcRCon_U8 ( .A1 (selSR), .A2 (calcRCon_n6), .ZN (calcRCon_n28) ) ;
    NAND2_X1 calcRCon_U7 ( .A1 (nReset), .A2 (calcRCon_n9), .ZN (calcRCon_n44) ) ;
    MUX2_X1 calcRCon_U6 ( .S (calcRCon_n5), .A (calcRCon_n16), .B (calcRCon_n11), .Z (calcRCon_n9) ) ;
    NAND2_X1 calcRCon_U5 ( .A1 (calcRCon_s_current_state_4_), .A2 (calcRCon_s_current_state_2_), .ZN (calcRCon_n7) ) ;
    NAND2_X1 calcRCon_U4 ( .A1 (calcRCon_s_current_state_1_), .A2 (calcRCon_s_current_state_5_), .ZN (calcRCon_n8) ) ;
    INV_X1 calcRCon_U3 ( .A (nReset), .ZN (calcRCon_n6) ) ;
    INV_X1 calcRCon_U2 ( .A (selSR), .ZN (calcRCon_n5) ) ;
    NOR2_X1 calcRCon_U1 ( .A1 (calcRCon_n8), .A2 (calcRCon_n7), .ZN (intFinal) ) ;
    INV_X1 calcRCon_s_current_state_reg_0__U1 ( .A (calcRCon_s_current_state_0_), .ZN (calcRCon_n13) ) ;
    INV_X1 calcRCon_s_current_state_reg_1__U1 ( .A (calcRCon_s_current_state_1_), .ZN (calcRCon_n14) ) ;
    INV_X1 calcRCon_s_current_state_reg_2__U1 ( .A (calcRCon_s_current_state_2_), .ZN (calcRCon_n12) ) ;
    INV_X1 calcRCon_s_current_state_reg_3__U1 ( .A (calcRCon_s_current_state_3_), .ZN (calcRCon_n15) ) ;
    INV_X1 calcRCon_s_current_state_reg_6__U1 ( .A (calcRCon_s_current_state_6_), .ZN (calcRCon_n16) ) ;
    INV_X1 calcRCon_s_current_state_reg_7__U1 ( .A (calcRCon_n3), .ZN (calcRCon_n11) ) ;
    mux2_masked_LMDPL MUX_SboxIn_mux_inst_0_U1 ( .s ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, selMC}), .b ({new_AGEMA_signal_1991, new_AGEMA_signal_1990, StateOutXORroundKey[0]}), .a ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, keySBIn[0]}), .c ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, SboxIn[0]}) ) ;
    mux2_masked_LMDPL MUX_SboxIn_mux_inst_1_U1 ( .s ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, selMC}), .b ({new_AGEMA_signal_1997, new_AGEMA_signal_1996, StateOutXORroundKey[1]}), .a ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, keySBIn[1]}), .c ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, SboxIn[1]}) ) ;
    mux2_masked_LMDPL MUX_SboxIn_mux_inst_2_U1 ( .s ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, selMC}), .b ({new_AGEMA_signal_2003, new_AGEMA_signal_2002, StateOutXORroundKey[2]}), .a ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, keySBIn[2]}), .c ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, SboxIn[2]}) ) ;
    mux2_masked_LMDPL MUX_SboxIn_mux_inst_3_U1 ( .s ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, selMC}), .b ({new_AGEMA_signal_2009, new_AGEMA_signal_2008, StateOutXORroundKey[3]}), .a ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, keySBIn[3]}), .c ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, SboxIn[3]}) ) ;
    mux2_masked_LMDPL MUX_SboxIn_mux_inst_4_U1 ( .s ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, selMC}), .b ({new_AGEMA_signal_2015, new_AGEMA_signal_2014, StateOutXORroundKey[4]}), .a ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, keySBIn[4]}), .c ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, SboxIn[4]}) ) ;
    mux2_masked_LMDPL MUX_SboxIn_mux_inst_5_U1 ( .s ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, selMC}), .b ({new_AGEMA_signal_2021, new_AGEMA_signal_2020, StateOutXORroundKey[5]}), .a ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, keySBIn[5]}), .c ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, SboxIn[5]}) ) ;
    mux2_masked_LMDPL MUX_SboxIn_mux_inst_6_U1 ( .s ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, selMC}), .b ({new_AGEMA_signal_2027, new_AGEMA_signal_2026, StateOutXORroundKey[6]}), .a ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, keySBIn[6]}), .c ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, SboxIn[6]}) ) ;
    mux2_masked_LMDPL MUX_SboxIn_mux_inst_7_U1 ( .s ({new_AGEMA_signal_3707, new_AGEMA_signal_3706, selMC}), .b ({new_AGEMA_signal_2033, new_AGEMA_signal_2032, StateOutXORroundKey[7]}), .a ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, keySBIn[7]}), .c ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, SboxIn[7]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T1_U1 ( .a ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, SboxIn[7]}), .b ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, SboxIn[4]}), .c ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Inst_bSbox_T1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T2_U1 ( .a ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, SboxIn[7]}), .b ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, SboxIn[2]}), .c ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Inst_bSbox_T2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T3_U1 ( .a ({new_AGEMA_signal_3723, new_AGEMA_signal_3722, SboxIn[7]}), .b ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, SboxIn[1]}), .c ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Inst_bSbox_T3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T4_U1 ( .a ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, SboxIn[4]}), .b ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, SboxIn[2]}), .c ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, Inst_bSbox_T4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T5_U1 ( .a ({new_AGEMA_signal_3715, new_AGEMA_signal_3714, SboxIn[3]}), .b ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, SboxIn[1]}), .c ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Inst_bSbox_T5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T6_U1 ( .a ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Inst_bSbox_T1}), .b ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Inst_bSbox_T5}), .c ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, Inst_bSbox_T6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T7_U1 ( .a ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, SboxIn[6]}), .b ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, SboxIn[5]}), .c ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Inst_bSbox_T7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T8_U1 ( .a ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, SboxIn[0]}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, Inst_bSbox_T6}), .c ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, Inst_bSbox_T8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T9_U1 ( .a ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, SboxIn[0]}), .b ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Inst_bSbox_T7}), .c ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, Inst_bSbox_T9}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T10_U1 ( .a ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, Inst_bSbox_T6}), .b ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Inst_bSbox_T7}), .c ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, Inst_bSbox_T10}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T11_U1 ( .a ({new_AGEMA_signal_3721, new_AGEMA_signal_3720, SboxIn[6]}), .b ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, SboxIn[2]}), .c ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Inst_bSbox_T11}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T12_U1 ( .a ({new_AGEMA_signal_3719, new_AGEMA_signal_3718, SboxIn[5]}), .b ({new_AGEMA_signal_3713, new_AGEMA_signal_3712, SboxIn[2]}), .c ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Inst_bSbox_T12}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T13_U1 ( .a ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Inst_bSbox_T3}), .b ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, Inst_bSbox_T4}), .c ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, Inst_bSbox_T13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T14_U1 ( .a ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, Inst_bSbox_T6}), .b ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Inst_bSbox_T11}), .c ({new_AGEMA_signal_4151, new_AGEMA_signal_4150, Inst_bSbox_T14}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T15_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Inst_bSbox_T5}), .b ({new_AGEMA_signal_3771, new_AGEMA_signal_3770, Inst_bSbox_T11}), .c ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, Inst_bSbox_T15}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T16_U1 ( .a ({new_AGEMA_signal_3767, new_AGEMA_signal_3766, Inst_bSbox_T5}), .b ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Inst_bSbox_T12}), .c ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, Inst_bSbox_T16}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T17_U1 ( .a ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, Inst_bSbox_T9}), .b ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, Inst_bSbox_T16}), .c ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, Inst_bSbox_T17}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T18_U1 ( .a ({new_AGEMA_signal_3717, new_AGEMA_signal_3716, SboxIn[4]}), .b ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, SboxIn[0]}), .c ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Inst_bSbox_T18}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T19_U1 ( .a ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Inst_bSbox_T7}), .b ({new_AGEMA_signal_3775, new_AGEMA_signal_3774, Inst_bSbox_T18}), .c ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, Inst_bSbox_T19}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T20_U1 ( .a ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Inst_bSbox_T1}), .b ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, Inst_bSbox_T19}), .c ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, Inst_bSbox_T20}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T21_U1 ( .a ({new_AGEMA_signal_3711, new_AGEMA_signal_3710, SboxIn[1]}), .b ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, SboxIn[0]}), .c ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Inst_bSbox_T21}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T22_U1 ( .a ({new_AGEMA_signal_3769, new_AGEMA_signal_3768, Inst_bSbox_T7}), .b ({new_AGEMA_signal_3777, new_AGEMA_signal_3776, Inst_bSbox_T21}), .c ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, Inst_bSbox_T22}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T23_U1 ( .a ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Inst_bSbox_T2}), .b ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, Inst_bSbox_T22}), .c ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, Inst_bSbox_T23}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T24_U1 ( .a ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Inst_bSbox_T2}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, Inst_bSbox_T10}), .c ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, Inst_bSbox_T24}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T25_U1 ( .a ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, Inst_bSbox_T20}), .b ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, Inst_bSbox_T17}), .c ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, Inst_bSbox_T25}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T26_U1 ( .a ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Inst_bSbox_T3}), .b ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, Inst_bSbox_T16}), .c ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, Inst_bSbox_T26}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_T27_U1 ( .a ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Inst_bSbox_T1}), .b ({new_AGEMA_signal_3773, new_AGEMA_signal_3772, Inst_bSbox_T12}), .c ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, Inst_bSbox_T27}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M1_U1 ( .a ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, Inst_bSbox_T13}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, Inst_bSbox_T6}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[0]), .c ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, Inst_bSbox_M1}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M2_U1 ( .a ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, Inst_bSbox_T23}), .b ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, Inst_bSbox_T8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[1]), .c ({new_AGEMA_signal_4325, new_AGEMA_signal_4324, Inst_bSbox_M2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M3_U1 ( .a ({new_AGEMA_signal_4151, new_AGEMA_signal_4150, Inst_bSbox_T14}), .b ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, Inst_bSbox_M1}), .c ({new_AGEMA_signal_4327, new_AGEMA_signal_4326, Inst_bSbox_M3}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M4_U1 ( .a ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, Inst_bSbox_T19}), .b ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, SboxIn[0]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[2]), .c ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, Inst_bSbox_M4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M5_U1 ( .a ({new_AGEMA_signal_4163, new_AGEMA_signal_4162, Inst_bSbox_M4}), .b ({new_AGEMA_signal_4161, new_AGEMA_signal_4160, Inst_bSbox_M1}), .c ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, Inst_bSbox_M5}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M6_U1 ( .a ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Inst_bSbox_T3}), .b ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, Inst_bSbox_T16}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[3]), .c ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, Inst_bSbox_M6}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M7_U1 ( .a ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, Inst_bSbox_T22}), .b ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, Inst_bSbox_T9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[4]), .c ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, Inst_bSbox_M7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M8_U1 ( .a ({new_AGEMA_signal_4159, new_AGEMA_signal_4158, Inst_bSbox_T26}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, Inst_bSbox_M6}), .c ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, Inst_bSbox_M8}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M9_U1 ( .a ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, Inst_bSbox_T20}), .b ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, Inst_bSbox_T17}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[5]), .c ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, Inst_bSbox_M9}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M10_U1 ( .a ({new_AGEMA_signal_4333, new_AGEMA_signal_4332, Inst_bSbox_M9}), .b ({new_AGEMA_signal_4165, new_AGEMA_signal_4164, Inst_bSbox_M6}), .c ({new_AGEMA_signal_4627, new_AGEMA_signal_4626, Inst_bSbox_M10}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M11_U1 ( .a ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Inst_bSbox_T1}), .b ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, Inst_bSbox_T15}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[6]), .c ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, Inst_bSbox_M11}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M12_U1 ( .a ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, Inst_bSbox_T4}), .b ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, Inst_bSbox_T27}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[7]), .c ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, Inst_bSbox_M12}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M13_U1 ( .a ({new_AGEMA_signal_4171, new_AGEMA_signal_4170, Inst_bSbox_M12}), .b ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, Inst_bSbox_M11}), .c ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, Inst_bSbox_M13}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M14_U1 ( .a ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Inst_bSbox_T2}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, Inst_bSbox_T10}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[8]), .c ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, Inst_bSbox_M14}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M15_U1 ( .a ({new_AGEMA_signal_4337, new_AGEMA_signal_4336, Inst_bSbox_M14}), .b ({new_AGEMA_signal_4169, new_AGEMA_signal_4168, Inst_bSbox_M11}), .c ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, Inst_bSbox_M15}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M16_U1 ( .a ({new_AGEMA_signal_4327, new_AGEMA_signal_4326, Inst_bSbox_M3}), .b ({new_AGEMA_signal_4325, new_AGEMA_signal_4324, Inst_bSbox_M2}), .c ({new_AGEMA_signal_4631, new_AGEMA_signal_4630, Inst_bSbox_M16}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M17_U1 ( .a ({new_AGEMA_signal_4329, new_AGEMA_signal_4328, Inst_bSbox_M5}), .b ({new_AGEMA_signal_4321, new_AGEMA_signal_4320, Inst_bSbox_T24}), .c ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, Inst_bSbox_M17}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M18_U1 ( .a ({new_AGEMA_signal_4331, new_AGEMA_signal_4330, Inst_bSbox_M8}), .b ({new_AGEMA_signal_4167, new_AGEMA_signal_4166, Inst_bSbox_M7}), .c ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, Inst_bSbox_M18}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M19_U1 ( .a ({new_AGEMA_signal_4627, new_AGEMA_signal_4626, Inst_bSbox_M10}), .b ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, Inst_bSbox_M15}), .c ({new_AGEMA_signal_4859, new_AGEMA_signal_4858, Inst_bSbox_M19}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M20_U1 ( .a ({new_AGEMA_signal_4631, new_AGEMA_signal_4630, Inst_bSbox_M16}), .b ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, Inst_bSbox_M13}), .c ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, Inst_bSbox_M20}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M21_U1 ( .a ({new_AGEMA_signal_4633, new_AGEMA_signal_4632, Inst_bSbox_M17}), .b ({new_AGEMA_signal_4629, new_AGEMA_signal_4628, Inst_bSbox_M15}), .c ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, Inst_bSbox_M21}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M22_U1 ( .a ({new_AGEMA_signal_4635, new_AGEMA_signal_4634, Inst_bSbox_M18}), .b ({new_AGEMA_signal_4335, new_AGEMA_signal_4334, Inst_bSbox_M13}), .c ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, Inst_bSbox_M22}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M23_U1 ( .a ({new_AGEMA_signal_4859, new_AGEMA_signal_4858, Inst_bSbox_M19}), .b ({new_AGEMA_signal_4323, new_AGEMA_signal_4322, Inst_bSbox_T25}), .c ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, Inst_bSbox_M23}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M24_U1 ( .a ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, Inst_bSbox_M22}), .b ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, Inst_bSbox_M23}), .c ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, Inst_bSbox_M24}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M25_U1 ( .a ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, Inst_bSbox_M22}), .b ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, Inst_bSbox_M20}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[9]), .c ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, Inst_bSbox_M25}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M26_U1 ( .a ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, Inst_bSbox_M21}), .b ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, Inst_bSbox_M25}), .c ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, Inst_bSbox_M26}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M27_U1 ( .a ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, Inst_bSbox_M20}), .b ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, Inst_bSbox_M21}), .c ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, Inst_bSbox_M27}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M28_U1 ( .a ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, Inst_bSbox_M23}), .b ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, Inst_bSbox_M25}), .c ({new_AGEMA_signal_4895, new_AGEMA_signal_4894, Inst_bSbox_M28}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M29_U1 ( .a ({new_AGEMA_signal_4895, new_AGEMA_signal_4894, Inst_bSbox_M28}), .b ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, Inst_bSbox_M27}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[10]), .c ({new_AGEMA_signal_4901, new_AGEMA_signal_4900, Inst_bSbox_M29}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M30_U1 ( .a ({new_AGEMA_signal_4893, new_AGEMA_signal_4892, Inst_bSbox_M26}), .b ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, Inst_bSbox_M24}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[11]), .c ({new_AGEMA_signal_4903, new_AGEMA_signal_4902, Inst_bSbox_M30}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M31_U1 ( .a ({new_AGEMA_signal_4861, new_AGEMA_signal_4860, Inst_bSbox_M20}), .b ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, Inst_bSbox_M23}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[12]), .c ({new_AGEMA_signal_4897, new_AGEMA_signal_4896, Inst_bSbox_M31}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M32_U1 ( .a ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, Inst_bSbox_M27}), .b ({new_AGEMA_signal_4897, new_AGEMA_signal_4896, Inst_bSbox_M31}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[13]), .c ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, Inst_bSbox_M32}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M33_U1 ( .a ({new_AGEMA_signal_4887, new_AGEMA_signal_4886, Inst_bSbox_M27}), .b ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, Inst_bSbox_M25}), .c ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, Inst_bSbox_M33}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M34_U1 ( .a ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, Inst_bSbox_M21}), .b ({new_AGEMA_signal_4865, new_AGEMA_signal_4864, Inst_bSbox_M22}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[14]), .c ({new_AGEMA_signal_4889, new_AGEMA_signal_4888, Inst_bSbox_M34}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M35_U1 ( .a ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, Inst_bSbox_M24}), .b ({new_AGEMA_signal_4889, new_AGEMA_signal_4888, Inst_bSbox_M34}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[15]), .c ({new_AGEMA_signal_4907, new_AGEMA_signal_4906, Inst_bSbox_M35}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M36_U1 ( .a ({new_AGEMA_signal_4891, new_AGEMA_signal_4890, Inst_bSbox_M24}), .b ({new_AGEMA_signal_4885, new_AGEMA_signal_4884, Inst_bSbox_M25}), .c ({new_AGEMA_signal_4909, new_AGEMA_signal_4908, Inst_bSbox_M36}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M37_U1 ( .a ({new_AGEMA_signal_4863, new_AGEMA_signal_4862, Inst_bSbox_M21}), .b ({new_AGEMA_signal_4901, new_AGEMA_signal_4900, Inst_bSbox_M29}), .c ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, Inst_bSbox_M37}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M38_U1 ( .a ({new_AGEMA_signal_4905, new_AGEMA_signal_4904, Inst_bSbox_M32}), .b ({new_AGEMA_signal_4899, new_AGEMA_signal_4898, Inst_bSbox_M33}), .c ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, Inst_bSbox_M38}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M39_U1 ( .a ({new_AGEMA_signal_4883, new_AGEMA_signal_4882, Inst_bSbox_M23}), .b ({new_AGEMA_signal_4903, new_AGEMA_signal_4902, Inst_bSbox_M30}), .c ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, Inst_bSbox_M39}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M40_U1 ( .a ({new_AGEMA_signal_4907, new_AGEMA_signal_4906, Inst_bSbox_M35}), .b ({new_AGEMA_signal_4909, new_AGEMA_signal_4908, Inst_bSbox_M36}), .c ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, Inst_bSbox_M40}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M41_U1 ( .a ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, Inst_bSbox_M38}), .b ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, Inst_bSbox_M40}), .c ({new_AGEMA_signal_4919, new_AGEMA_signal_4918, Inst_bSbox_M41}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M42_U1 ( .a ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, Inst_bSbox_M37}), .b ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, Inst_bSbox_M39}), .c ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, Inst_bSbox_M42}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M43_U1 ( .a ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, Inst_bSbox_M37}), .b ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, Inst_bSbox_M38}), .c ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, Inst_bSbox_M43}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M44_U1 ( .a ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, Inst_bSbox_M39}), .b ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, Inst_bSbox_M40}), .c ({new_AGEMA_signal_4925, new_AGEMA_signal_4924, Inst_bSbox_M44}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_M45_U1 ( .a ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, Inst_bSbox_M42}), .b ({new_AGEMA_signal_4919, new_AGEMA_signal_4918, Inst_bSbox_M41}), .c ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, Inst_bSbox_M45}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M46_U1 ( .a ({new_AGEMA_signal_4925, new_AGEMA_signal_4924, Inst_bSbox_M44}), .b ({new_AGEMA_signal_4079, new_AGEMA_signal_4078, Inst_bSbox_T6}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[16]), .c ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, Inst_bSbox_M46}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M47_U1 ( .a ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, Inst_bSbox_M40}), .b ({new_AGEMA_signal_4147, new_AGEMA_signal_4146, Inst_bSbox_T8}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[17]), .c ({new_AGEMA_signal_4927, new_AGEMA_signal_4926, Inst_bSbox_M47}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M48_U1 ( .a ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, Inst_bSbox_M39}), .b ({new_AGEMA_signal_3709, new_AGEMA_signal_3708, SboxIn[0]}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[18]), .c ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, Inst_bSbox_M48}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M49_U1 ( .a ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, Inst_bSbox_M43}), .b ({new_AGEMA_signal_4087, new_AGEMA_signal_4086, Inst_bSbox_T16}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[19]), .c ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, Inst_bSbox_M49}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M50_U1 ( .a ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, Inst_bSbox_M38}), .b ({new_AGEMA_signal_4081, new_AGEMA_signal_4080, Inst_bSbox_T9}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[20]), .c ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, Inst_bSbox_M50}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M51_U1 ( .a ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, Inst_bSbox_M37}), .b ({new_AGEMA_signal_4153, new_AGEMA_signal_4152, Inst_bSbox_T17}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[21]), .c ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, Inst_bSbox_M51}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M52_U1 ( .a ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, Inst_bSbox_M42}), .b ({new_AGEMA_signal_4085, new_AGEMA_signal_4084, Inst_bSbox_T15}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[22]), .c ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, Inst_bSbox_M52}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M53_U1 ( .a ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, Inst_bSbox_M45}), .b ({new_AGEMA_signal_4093, new_AGEMA_signal_4092, Inst_bSbox_T27}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[23]), .c ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, Inst_bSbox_M53}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M54_U1 ( .a ({new_AGEMA_signal_4919, new_AGEMA_signal_4918, Inst_bSbox_M41}), .b ({new_AGEMA_signal_4149, new_AGEMA_signal_4148, Inst_bSbox_T10}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[24]), .c ({new_AGEMA_signal_4951, new_AGEMA_signal_4950, Inst_bSbox_M54}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M55_U1 ( .a ({new_AGEMA_signal_4925, new_AGEMA_signal_4924, Inst_bSbox_M44}), .b ({new_AGEMA_signal_4083, new_AGEMA_signal_4082, Inst_bSbox_T13}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[25]), .c ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, Inst_bSbox_M55}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M56_U1 ( .a ({new_AGEMA_signal_4917, new_AGEMA_signal_4916, Inst_bSbox_M40}), .b ({new_AGEMA_signal_4157, new_AGEMA_signal_4156, Inst_bSbox_T23}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[26]), .c ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, Inst_bSbox_M56}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M57_U1 ( .a ({new_AGEMA_signal_4915, new_AGEMA_signal_4914, Inst_bSbox_M39}), .b ({new_AGEMA_signal_4089, new_AGEMA_signal_4088, Inst_bSbox_T19}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[27]), .c ({new_AGEMA_signal_4937, new_AGEMA_signal_4936, Inst_bSbox_M57}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M58_U1 ( .a ({new_AGEMA_signal_4923, new_AGEMA_signal_4922, Inst_bSbox_M43}), .b ({new_AGEMA_signal_3763, new_AGEMA_signal_3762, Inst_bSbox_T3}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[28]), .c ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, Inst_bSbox_M58}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M59_U1 ( .a ({new_AGEMA_signal_4913, new_AGEMA_signal_4912, Inst_bSbox_M38}), .b ({new_AGEMA_signal_4091, new_AGEMA_signal_4090, Inst_bSbox_T22}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[29]), .c ({new_AGEMA_signal_4939, new_AGEMA_signal_4938, Inst_bSbox_M59}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M60_U1 ( .a ({new_AGEMA_signal_4911, new_AGEMA_signal_4910, Inst_bSbox_M37}), .b ({new_AGEMA_signal_4155, new_AGEMA_signal_4154, Inst_bSbox_T20}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[30]), .c ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, Inst_bSbox_M60}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M61_U1 ( .a ({new_AGEMA_signal_4921, new_AGEMA_signal_4920, Inst_bSbox_M42}), .b ({new_AGEMA_signal_3759, new_AGEMA_signal_3758, Inst_bSbox_T1}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[31]), .c ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, Inst_bSbox_M61}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M62_U1 ( .a ({new_AGEMA_signal_4943, new_AGEMA_signal_4942, Inst_bSbox_M45}), .b ({new_AGEMA_signal_3765, new_AGEMA_signal_3764, Inst_bSbox_T4}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[32]), .c ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, Inst_bSbox_M62}) ) ;
    nonlinear_LMDPL #(.CONF(2'b00)) Inst_bSbox_AND_M63_U1 ( .a ({new_AGEMA_signal_4919, new_AGEMA_signal_4918, Inst_bSbox_M41}), .b ({new_AGEMA_signal_3761, new_AGEMA_signal_3760, Inst_bSbox_T2}), .mid_rst (mid_rst), .clk (clk), .r (Fresh[33]), .c ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, Inst_bSbox_M63}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L0_U1 ( .a ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, Inst_bSbox_M61}), .b ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, Inst_bSbox_M62}), .c ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, Inst_bSbox_L0}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L1_U1 ( .a ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, Inst_bSbox_M50}), .b ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, Inst_bSbox_M56}), .c ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, Inst_bSbox_L1}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L2_U1 ( .a ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, Inst_bSbox_M46}), .b ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, Inst_bSbox_M48}), .c ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, Inst_bSbox_L2}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L3_U1 ( .a ({new_AGEMA_signal_4927, new_AGEMA_signal_4926, Inst_bSbox_M47}), .b ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, Inst_bSbox_M55}), .c ({new_AGEMA_signal_4973, new_AGEMA_signal_4972, Inst_bSbox_L3}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L4_U1 ( .a ({new_AGEMA_signal_4951, new_AGEMA_signal_4950, Inst_bSbox_M54}), .b ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, Inst_bSbox_M58}), .c ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, Inst_bSbox_L4}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L5_U1 ( .a ({new_AGEMA_signal_4947, new_AGEMA_signal_4946, Inst_bSbox_M49}), .b ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, Inst_bSbox_M61}), .c ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, Inst_bSbox_L5}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L6_U1 ( .a ({new_AGEMA_signal_4969, new_AGEMA_signal_4968, Inst_bSbox_M62}), .b ({new_AGEMA_signal_4977, new_AGEMA_signal_4976, Inst_bSbox_L5}), .c ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, Inst_bSbox_L6}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L7_U1 ( .a ({new_AGEMA_signal_4945, new_AGEMA_signal_4944, Inst_bSbox_M46}), .b ({new_AGEMA_signal_4973, new_AGEMA_signal_4972, Inst_bSbox_L3}), .c ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, Inst_bSbox_L7}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L8_U1 ( .a ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, Inst_bSbox_M51}), .b ({new_AGEMA_signal_4939, new_AGEMA_signal_4938, Inst_bSbox_M59}), .c ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, Inst_bSbox_L8}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L9_U1 ( .a ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, Inst_bSbox_M52}), .b ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, Inst_bSbox_M53}), .c ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, Inst_bSbox_L9}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L10_U1 ( .a ({new_AGEMA_signal_4967, new_AGEMA_signal_4966, Inst_bSbox_M53}), .b ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, Inst_bSbox_L4}), .c ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, Inst_bSbox_L10}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L11_U1 ( .a ({new_AGEMA_signal_4941, new_AGEMA_signal_4940, Inst_bSbox_M60}), .b ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, Inst_bSbox_L2}), .c ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, Inst_bSbox_L11}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L12_U1 ( .a ({new_AGEMA_signal_4929, new_AGEMA_signal_4928, Inst_bSbox_M48}), .b ({new_AGEMA_signal_4933, new_AGEMA_signal_4932, Inst_bSbox_M51}), .c ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, Inst_bSbox_L12}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L13_U1 ( .a ({new_AGEMA_signal_4931, new_AGEMA_signal_4930, Inst_bSbox_M50}), .b ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, Inst_bSbox_L0}), .c ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, Inst_bSbox_L13}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L14_U1 ( .a ({new_AGEMA_signal_4949, new_AGEMA_signal_4948, Inst_bSbox_M52}), .b ({new_AGEMA_signal_4957, new_AGEMA_signal_4956, Inst_bSbox_M61}), .c ({new_AGEMA_signal_4979, new_AGEMA_signal_4978, Inst_bSbox_L14}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L15_U1 ( .a ({new_AGEMA_signal_4953, new_AGEMA_signal_4952, Inst_bSbox_M55}), .b ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, Inst_bSbox_L1}), .c ({new_AGEMA_signal_4981, new_AGEMA_signal_4980, Inst_bSbox_L15}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L16_U1 ( .a ({new_AGEMA_signal_4935, new_AGEMA_signal_4934, Inst_bSbox_M56}), .b ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, Inst_bSbox_L0}), .c ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, Inst_bSbox_L16}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L17_U1 ( .a ({new_AGEMA_signal_4937, new_AGEMA_signal_4936, Inst_bSbox_M57}), .b ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, Inst_bSbox_L1}), .c ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, Inst_bSbox_L17}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L18_U1 ( .a ({new_AGEMA_signal_4955, new_AGEMA_signal_4954, Inst_bSbox_M58}), .b ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, Inst_bSbox_L8}), .c ({new_AGEMA_signal_4985, new_AGEMA_signal_4984, Inst_bSbox_L18}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L19_U1 ( .a ({new_AGEMA_signal_4959, new_AGEMA_signal_4958, Inst_bSbox_M63}), .b ({new_AGEMA_signal_4975, new_AGEMA_signal_4974, Inst_bSbox_L4}), .c ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, Inst_bSbox_L19}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L20_U1 ( .a ({new_AGEMA_signal_4987, new_AGEMA_signal_4986, Inst_bSbox_L0}), .b ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, Inst_bSbox_L1}), .c ({new_AGEMA_signal_5009, new_AGEMA_signal_5008, Inst_bSbox_L20}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L21_U1 ( .a ({new_AGEMA_signal_4961, new_AGEMA_signal_4960, Inst_bSbox_L1}), .b ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, Inst_bSbox_L7}), .c ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, Inst_bSbox_L21}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L22_U1 ( .a ({new_AGEMA_signal_4973, new_AGEMA_signal_4972, Inst_bSbox_L3}), .b ({new_AGEMA_signal_4965, new_AGEMA_signal_4964, Inst_bSbox_L12}), .c ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, Inst_bSbox_L22}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L23_U1 ( .a ({new_AGEMA_signal_4985, new_AGEMA_signal_4984, Inst_bSbox_L18}), .b ({new_AGEMA_signal_4971, new_AGEMA_signal_4970, Inst_bSbox_L2}), .c ({new_AGEMA_signal_5003, new_AGEMA_signal_5002, Inst_bSbox_L23}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L24_U1 ( .a ({new_AGEMA_signal_4981, new_AGEMA_signal_4980, Inst_bSbox_L15}), .b ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, Inst_bSbox_L9}), .c ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, Inst_bSbox_L24}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L25_U1 ( .a ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, Inst_bSbox_L6}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, Inst_bSbox_L10}), .c ({new_AGEMA_signal_5015, new_AGEMA_signal_5014, Inst_bSbox_L25}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L26_U1 ( .a ({new_AGEMA_signal_4991, new_AGEMA_signal_4990, Inst_bSbox_L7}), .b ({new_AGEMA_signal_4993, new_AGEMA_signal_4992, Inst_bSbox_L9}), .c ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, Inst_bSbox_L26}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L27_U1 ( .a ({new_AGEMA_signal_4963, new_AGEMA_signal_4962, Inst_bSbox_L8}), .b ({new_AGEMA_signal_4995, new_AGEMA_signal_4994, Inst_bSbox_L10}), .c ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, Inst_bSbox_L27}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L28_U1 ( .a ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, Inst_bSbox_L11}), .b ({new_AGEMA_signal_4979, new_AGEMA_signal_4978, Inst_bSbox_L14}), .c ({new_AGEMA_signal_5021, new_AGEMA_signal_5020, Inst_bSbox_L28}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_L29_U1 ( .a ({new_AGEMA_signal_4997, new_AGEMA_signal_4996, Inst_bSbox_L11}), .b ({new_AGEMA_signal_4983, new_AGEMA_signal_4982, Inst_bSbox_L17}), .c ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, Inst_bSbox_L29}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_S0_U1 ( .a ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, Inst_bSbox_L6}), .b ({new_AGEMA_signal_5013, new_AGEMA_signal_5012, Inst_bSbox_L24}), .c ({new_AGEMA_signal_5031, new_AGEMA_signal_5030, SboxOut[7]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) Inst_bSbox_XOR_S1_U1 ( .a ({new_AGEMA_signal_5007, new_AGEMA_signal_5006, Inst_bSbox_L16}), .b ({new_AGEMA_signal_5017, new_AGEMA_signal_5016, Inst_bSbox_L26}), .c ({new_AGEMA_signal_5033, new_AGEMA_signal_5032, SboxOut[6]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) Inst_bSbox_XOR_S2_U1 ( .a ({new_AGEMA_signal_4999, new_AGEMA_signal_4998, Inst_bSbox_L19}), .b ({new_AGEMA_signal_5021, new_AGEMA_signal_5020, Inst_bSbox_L28}), .c ({new_AGEMA_signal_5035, new_AGEMA_signal_5034, SboxOut[5]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_S3_U1 ( .a ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, Inst_bSbox_L6}), .b ({new_AGEMA_signal_5011, new_AGEMA_signal_5010, Inst_bSbox_L21}), .c ({new_AGEMA_signal_5037, new_AGEMA_signal_5036, SboxOut[4]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_S4_U1 ( .a ({new_AGEMA_signal_5009, new_AGEMA_signal_5008, Inst_bSbox_L20}), .b ({new_AGEMA_signal_5001, new_AGEMA_signal_5000, Inst_bSbox_L22}), .c ({new_AGEMA_signal_5039, new_AGEMA_signal_5038, SboxOut[3]}) ) ;
    linear_LMDPL #(.CONF(1'b0)) Inst_bSbox_XOR_S5_U1 ( .a ({new_AGEMA_signal_5015, new_AGEMA_signal_5014, Inst_bSbox_L25}), .b ({new_AGEMA_signal_5023, new_AGEMA_signal_5022, Inst_bSbox_L29}), .c ({new_AGEMA_signal_5041, new_AGEMA_signal_5040, SboxOut[2]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) Inst_bSbox_XOR_S6_U1 ( .a ({new_AGEMA_signal_5005, new_AGEMA_signal_5004, Inst_bSbox_L13}), .b ({new_AGEMA_signal_5019, new_AGEMA_signal_5018, Inst_bSbox_L27}), .c ({new_AGEMA_signal_5043, new_AGEMA_signal_5042, SboxOut[1]}) ) ;
    linear_LMDPL #(.CONF(1'b1)) Inst_bSbox_XOR_S7_U1 ( .a ({new_AGEMA_signal_4989, new_AGEMA_signal_4988, Inst_bSbox_L6}), .b ({new_AGEMA_signal_5003, new_AGEMA_signal_5002, Inst_bSbox_L23}), .c ({new_AGEMA_signal_5025, new_AGEMA_signal_5024, SboxOut[0]}) ) ;
    INV_X1 nReset_reg_U1 ( .A (nReset), .ZN (n10) ) ;
    Precharger_reg new_AGEMA_gate_1714 ( .D (stateArray_n32), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2331, new_AGEMA_signal_2330}) ) ;
    Precharger_reg new_AGEMA_gate_1715 ( .D (stateArray_n31), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2429, new_AGEMA_signal_2428}) ) ;
    Precharger_reg new_AGEMA_gate_1716 ( .D (stateArray_n30), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2479, new_AGEMA_signal_2478}) ) ;
    Precharger_reg new_AGEMA_gate_1717 ( .D (stateArray_n29), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2577, new_AGEMA_signal_2576}) ) ;
    Precharger_reg new_AGEMA_gate_1718 ( .D (stateArray_n28), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2627, new_AGEMA_signal_2626}) ) ;
    Precharger_reg new_AGEMA_gate_1719 ( .D (stateArray_n27), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2725, new_AGEMA_signal_2724}) ) ;
    Precharger_reg new_AGEMA_gate_1720 ( .D (stateArray_n26), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2775, new_AGEMA_signal_2774}) ) ;
    Precharger_reg new_AGEMA_gate_1721 ( .D (stateArray_n25), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2873, new_AGEMA_signal_2872}) ) ;
    Precharger_reg new_AGEMA_gate_1722 ( .D (KeyArray_n46), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2923, new_AGEMA_signal_2922}) ) ;
    Precharger_reg new_AGEMA_gate_1723 ( .D (KeyArray_n45), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_2973, new_AGEMA_signal_2972}) ) ;
    Precharger_reg new_AGEMA_gate_1724 ( .D (KeyArray_n44), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3071, new_AGEMA_signal_3070}) ) ;
    Precharger_reg new_AGEMA_gate_1725 ( .D (KeyArray_n43), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3169, new_AGEMA_signal_3168}) ) ;
    Precharger_reg new_AGEMA_gate_1726 ( .D (KeyArray_n42), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3267, new_AGEMA_signal_3266}) ) ;
    Precharger_reg new_AGEMA_gate_1727 ( .D (KeyArray_n41), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3365, new_AGEMA_signal_3364}) ) ;
    Precharger_reg new_AGEMA_gate_1728 ( .D (KeyArray_n40), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3463, new_AGEMA_signal_3462}) ) ;
    Precharger_reg new_AGEMA_gate_1729 ( .D (KeyArray_n39), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3561, new_AGEMA_signal_3560}) ) ;
    Precharger_reg new_AGEMA_gate_1730 ( .D (selMC), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3707, new_AGEMA_signal_3706}) ) ;
    Precharger_reg new_AGEMA_gate_1731 ( .D (intFinal), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3725, new_AGEMA_signal_3724}) ) ;
    Precharger_reg new_AGEMA_gate_1732 ( .D (MUX_StateInMC_n5), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3779, new_AGEMA_signal_3778}) ) ;
    Precharger_reg new_AGEMA_gate_1733 ( .D (MUX_StateInMC_n6), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3783, new_AGEMA_signal_3782}) ) ;
    Precharger_reg new_AGEMA_gate_1734 ( .D (KeyArray_n37), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3839, new_AGEMA_signal_3838}) ) ;
    Precharger_reg new_AGEMA_gate_1735 ( .D (KeyArray_n36), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3857, new_AGEMA_signal_3856}) ) ;
    Precharger_reg new_AGEMA_gate_1736 ( .D (KeyArray_n35), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3891, new_AGEMA_signal_3890}) ) ;
    Precharger_reg new_AGEMA_gate_1737 ( .D (KeyArray_n34), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3925, new_AGEMA_signal_3924}) ) ;
    Precharger_reg new_AGEMA_gate_1738 ( .D (KeyArray_n33), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3959, new_AGEMA_signal_3958}) ) ;
    Precharger_reg new_AGEMA_gate_1739 ( .D (KeyArray_n32), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_3993, new_AGEMA_signal_3992}) ) ;
    Precharger_reg new_AGEMA_gate_1740 ( .D (KeyArray_n31), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4027, new_AGEMA_signal_4026}) ) ;
    Precharger_reg new_AGEMA_gate_1741 ( .D (KeyArray_n30), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4045, new_AGEMA_signal_4044}) ) ;
    Precharger_reg new_AGEMA_gate_1742 ( .D (stateArray_n23), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4095, new_AGEMA_signal_4094}) ) ;
    Precharger_reg new_AGEMA_gate_1743 ( .D (stateArray_n22), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4129, new_AGEMA_signal_4128}) ) ;
    Precharger_reg new_AGEMA_gate_1744 ( .D (n12), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4269, new_AGEMA_signal_4268}) ) ;
    Precharger_reg new_AGEMA_gate_1745 ( .D (intselXOR), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4303, new_AGEMA_signal_4302}) ) ;
    Precharger_reg new_AGEMA_gate_1746 ( .D (stateArray_n20), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4339, new_AGEMA_signal_4338}) ) ;
    Precharger_reg new_AGEMA_gate_1747 ( .D (stateArray_n19), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4373, new_AGEMA_signal_4372}) ) ;
    Precharger_reg new_AGEMA_gate_1748 ( .D (stateArray_n18), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4407, new_AGEMA_signal_4406}) ) ;
    Precharger_reg new_AGEMA_gate_1749 ( .D (stateArray_n17), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4441, new_AGEMA_signal_4440}) ) ;
    Precharger_reg new_AGEMA_gate_1750 ( .D (stateArray_n16), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4475, new_AGEMA_signal_4474}) ) ;
    Precharger_reg new_AGEMA_gate_1751 ( .D (stateArray_n15), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4509, new_AGEMA_signal_4508}) ) ;
    Precharger_reg new_AGEMA_gate_1752 ( .D (stateArray_n14), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4543, new_AGEMA_signal_4542}) ) ;
    Precharger_reg new_AGEMA_gate_1753 ( .D (stateArray_n13), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4577, new_AGEMA_signal_4576}) ) ;
    Precharger_reg new_AGEMA_gate_1754 ( .D (KeyArray_n28), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4653, new_AGEMA_signal_4652}) ) ;
    Precharger_reg new_AGEMA_gate_1755 ( .D (KeyArray_n27), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4671, new_AGEMA_signal_4670}) ) ;
    Precharger_reg new_AGEMA_gate_1756 ( .D (KeyArray_n26), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4705, new_AGEMA_signal_4704}) ) ;
    Precharger_reg new_AGEMA_gate_1757 ( .D (KeyArray_n25), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4739, new_AGEMA_signal_4738}) ) ;
    Precharger_reg new_AGEMA_gate_1758 ( .D (KeyArray_n24), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4773, new_AGEMA_signal_4772}) ) ;
    Precharger_reg new_AGEMA_gate_1759 ( .D (KeyArray_n23), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4807, new_AGEMA_signal_4806}) ) ;
    Precharger_reg new_AGEMA_gate_1760 ( .D (KeyArray_n22), .mid_rst (mid_rst), .clk (clk), .Q ({new_AGEMA_signal_4825, new_AGEMA_signal_4824}) ) ;
    ClockController_LMDPL ClockControllerInst ( .clk (clk), .Po_rst (Po_rst), .pre1 (LMDPL_pre1), .pre2 (LMDPL_pre2), .mid_rst (mid_rst) ) ;
    Precharger PrechargeCell_0 ( .D (plaintext_s1[127]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2375, new_AGEMA_signal_2374}) ) ;
    Precharger PrechargeCell_1 ( .D (plaintext_s1[126]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2369, new_AGEMA_signal_2368}) ) ;
    Precharger PrechargeCell_2 ( .D (plaintext_s1[125]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2363, new_AGEMA_signal_2362}) ) ;
    Precharger PrechargeCell_3 ( .D (plaintext_s1[124]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2357, new_AGEMA_signal_2356}) ) ;
    Precharger PrechargeCell_4 ( .D (plaintext_s1[123]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2351, new_AGEMA_signal_2350}) ) ;
    Precharger PrechargeCell_5 ( .D (plaintext_s1[122]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2345, new_AGEMA_signal_2344}) ) ;
    Precharger PrechargeCell_6 ( .D (plaintext_s1[121]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2339, new_AGEMA_signal_2338}) ) ;
    Precharger PrechargeCell_7 ( .D (plaintext_s1[120]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2333, new_AGEMA_signal_2332}) ) ;
    Precharger PrechargeCell_8 ( .D (plaintext_s1[119]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2423, new_AGEMA_signal_2422}) ) ;
    Precharger PrechargeCell_9 ( .D (plaintext_s1[118]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2417, new_AGEMA_signal_2416}) ) ;
    Precharger PrechargeCell_10 ( .D (plaintext_s1[117]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2411, new_AGEMA_signal_2410}) ) ;
    Precharger PrechargeCell_11 ( .D (plaintext_s1[116]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2405, new_AGEMA_signal_2404}) ) ;
    Precharger PrechargeCell_12 ( .D (plaintext_s1[115]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2399, new_AGEMA_signal_2398}) ) ;
    Precharger PrechargeCell_13 ( .D (plaintext_s1[114]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2393, new_AGEMA_signal_2392}) ) ;
    Precharger PrechargeCell_14 ( .D (plaintext_s1[113]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2387, new_AGEMA_signal_2386}) ) ;
    Precharger PrechargeCell_15 ( .D (plaintext_s1[112]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2381, new_AGEMA_signal_2380}) ) ;
    Precharger PrechargeCell_16 ( .D (plaintext_s1[111]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2473, new_AGEMA_signal_2472}) ) ;
    Precharger PrechargeCell_17 ( .D (plaintext_s1[110]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2467, new_AGEMA_signal_2466}) ) ;
    Precharger PrechargeCell_18 ( .D (plaintext_s1[109]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2461, new_AGEMA_signal_2460}) ) ;
    Precharger PrechargeCell_19 ( .D (plaintext_s1[108]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2455, new_AGEMA_signal_2454}) ) ;
    Precharger PrechargeCell_20 ( .D (plaintext_s1[107]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2449, new_AGEMA_signal_2448}) ) ;
    Precharger PrechargeCell_21 ( .D (plaintext_s1[106]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2443, new_AGEMA_signal_2442}) ) ;
    Precharger PrechargeCell_22 ( .D (plaintext_s1[105]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2437, new_AGEMA_signal_2436}) ) ;
    Precharger PrechargeCell_23 ( .D (plaintext_s1[104]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2431, new_AGEMA_signal_2430}) ) ;
    Precharger PrechargeCell_24 ( .D (plaintext_s1[103]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4201, new_AGEMA_signal_4200}) ) ;
    Precharger PrechargeCell_25 ( .D (plaintext_s1[102]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4197, new_AGEMA_signal_4196}) ) ;
    Precharger PrechargeCell_26 ( .D (plaintext_s1[101]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4193, new_AGEMA_signal_4192}) ) ;
    Precharger PrechargeCell_27 ( .D (plaintext_s1[100]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4189, new_AGEMA_signal_4188}) ) ;
    Precharger PrechargeCell_28 ( .D (plaintext_s1[99]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4185, new_AGEMA_signal_4184}) ) ;
    Precharger PrechargeCell_29 ( .D (plaintext_s1[98]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4181, new_AGEMA_signal_4180}) ) ;
    Precharger PrechargeCell_30 ( .D (plaintext_s1[97]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4177, new_AGEMA_signal_4176}) ) ;
    Precharger PrechargeCell_31 ( .D (plaintext_s1[96]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4173, new_AGEMA_signal_4172}) ) ;
    Precharger PrechargeCell_32 ( .D (plaintext_s1[95]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2523, new_AGEMA_signal_2522}) ) ;
    Precharger PrechargeCell_33 ( .D (plaintext_s1[94]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2517, new_AGEMA_signal_2516}) ) ;
    Precharger PrechargeCell_34 ( .D (plaintext_s1[93]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2511, new_AGEMA_signal_2510}) ) ;
    Precharger PrechargeCell_35 ( .D (plaintext_s1[92]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2505, new_AGEMA_signal_2504}) ) ;
    Precharger PrechargeCell_36 ( .D (plaintext_s1[91]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2499, new_AGEMA_signal_2498}) ) ;
    Precharger PrechargeCell_37 ( .D (plaintext_s1[90]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2493, new_AGEMA_signal_2492}) ) ;
    Precharger PrechargeCell_38 ( .D (plaintext_s1[89]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2487, new_AGEMA_signal_2486}) ) ;
    Precharger PrechargeCell_39 ( .D (plaintext_s1[88]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2481, new_AGEMA_signal_2480}) ) ;
    Precharger PrechargeCell_40 ( .D (plaintext_s1[87]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2571, new_AGEMA_signal_2570}) ) ;
    Precharger PrechargeCell_41 ( .D (plaintext_s1[86]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2565, new_AGEMA_signal_2564}) ) ;
    Precharger PrechargeCell_42 ( .D (plaintext_s1[85]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2559, new_AGEMA_signal_2558}) ) ;
    Precharger PrechargeCell_43 ( .D (plaintext_s1[84]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2553, new_AGEMA_signal_2552}) ) ;
    Precharger PrechargeCell_44 ( .D (plaintext_s1[83]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2547, new_AGEMA_signal_2546}) ) ;
    Precharger PrechargeCell_45 ( .D (plaintext_s1[82]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2541, new_AGEMA_signal_2540}) ) ;
    Precharger PrechargeCell_46 ( .D (plaintext_s1[81]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2535, new_AGEMA_signal_2534}) ) ;
    Precharger PrechargeCell_47 ( .D (plaintext_s1[80]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2529, new_AGEMA_signal_2528}) ) ;
    Precharger PrechargeCell_48 ( .D (plaintext_s1[79]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2621, new_AGEMA_signal_2620}) ) ;
    Precharger PrechargeCell_49 ( .D (plaintext_s1[78]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2615, new_AGEMA_signal_2614}) ) ;
    Precharger PrechargeCell_50 ( .D (plaintext_s1[77]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2609, new_AGEMA_signal_2608}) ) ;
    Precharger PrechargeCell_51 ( .D (plaintext_s1[76]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2603, new_AGEMA_signal_2602}) ) ;
    Precharger PrechargeCell_52 ( .D (plaintext_s1[75]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2597, new_AGEMA_signal_2596}) ) ;
    Precharger PrechargeCell_53 ( .D (plaintext_s1[74]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2591, new_AGEMA_signal_2590}) ) ;
    Precharger PrechargeCell_54 ( .D (plaintext_s1[73]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2585, new_AGEMA_signal_2584}) ) ;
    Precharger PrechargeCell_55 ( .D (plaintext_s1[72]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2579, new_AGEMA_signal_2578}) ) ;
    Precharger PrechargeCell_56 ( .D (plaintext_s1[71]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4233, new_AGEMA_signal_4232}) ) ;
    Precharger PrechargeCell_57 ( .D (plaintext_s1[70]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4229, new_AGEMA_signal_4228}) ) ;
    Precharger PrechargeCell_58 ( .D (plaintext_s1[69]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4225, new_AGEMA_signal_4224}) ) ;
    Precharger PrechargeCell_59 ( .D (plaintext_s1[68]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4221, new_AGEMA_signal_4220}) ) ;
    Precharger PrechargeCell_60 ( .D (plaintext_s1[67]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4217, new_AGEMA_signal_4216}) ) ;
    Precharger PrechargeCell_61 ( .D (plaintext_s1[66]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4213, new_AGEMA_signal_4212}) ) ;
    Precharger PrechargeCell_62 ( .D (plaintext_s1[65]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4209, new_AGEMA_signal_4208}) ) ;
    Precharger PrechargeCell_63 ( .D (plaintext_s1[64]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4205, new_AGEMA_signal_4204}) ) ;
    Precharger PrechargeCell_64 ( .D (plaintext_s1[63]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2671, new_AGEMA_signal_2670}) ) ;
    Precharger PrechargeCell_65 ( .D (plaintext_s1[62]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2665, new_AGEMA_signal_2664}) ) ;
    Precharger PrechargeCell_66 ( .D (plaintext_s1[61]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2659, new_AGEMA_signal_2658}) ) ;
    Precharger PrechargeCell_67 ( .D (plaintext_s1[60]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2653, new_AGEMA_signal_2652}) ) ;
    Precharger PrechargeCell_68 ( .D (plaintext_s1[59]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2647, new_AGEMA_signal_2646}) ) ;
    Precharger PrechargeCell_69 ( .D (plaintext_s1[58]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2641, new_AGEMA_signal_2640}) ) ;
    Precharger PrechargeCell_70 ( .D (plaintext_s1[57]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2635, new_AGEMA_signal_2634}) ) ;
    Precharger PrechargeCell_71 ( .D (plaintext_s1[56]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2629, new_AGEMA_signal_2628}) ) ;
    Precharger PrechargeCell_72 ( .D (plaintext_s1[55]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2719, new_AGEMA_signal_2718}) ) ;
    Precharger PrechargeCell_73 ( .D (plaintext_s1[54]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2713, new_AGEMA_signal_2712}) ) ;
    Precharger PrechargeCell_74 ( .D (plaintext_s1[53]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2707, new_AGEMA_signal_2706}) ) ;
    Precharger PrechargeCell_75 ( .D (plaintext_s1[52]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2701, new_AGEMA_signal_2700}) ) ;
    Precharger PrechargeCell_76 ( .D (plaintext_s1[51]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2695, new_AGEMA_signal_2694}) ) ;
    Precharger PrechargeCell_77 ( .D (plaintext_s1[50]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2689, new_AGEMA_signal_2688}) ) ;
    Precharger PrechargeCell_78 ( .D (plaintext_s1[49]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2683, new_AGEMA_signal_2682}) ) ;
    Precharger PrechargeCell_79 ( .D (plaintext_s1[48]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2677, new_AGEMA_signal_2676}) ) ;
    Precharger PrechargeCell_80 ( .D (plaintext_s1[47]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2769, new_AGEMA_signal_2768}) ) ;
    Precharger PrechargeCell_81 ( .D (plaintext_s1[46]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2763, new_AGEMA_signal_2762}) ) ;
    Precharger PrechargeCell_82 ( .D (plaintext_s1[45]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2757, new_AGEMA_signal_2756}) ) ;
    Precharger PrechargeCell_83 ( .D (plaintext_s1[44]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2751, new_AGEMA_signal_2750}) ) ;
    Precharger PrechargeCell_84 ( .D (plaintext_s1[43]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2745, new_AGEMA_signal_2744}) ) ;
    Precharger PrechargeCell_85 ( .D (plaintext_s1[42]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2739, new_AGEMA_signal_2738}) ) ;
    Precharger PrechargeCell_86 ( .D (plaintext_s1[41]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2733, new_AGEMA_signal_2732}) ) ;
    Precharger PrechargeCell_87 ( .D (plaintext_s1[40]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2727, new_AGEMA_signal_2726}) ) ;
    Precharger PrechargeCell_88 ( .D (plaintext_s1[39]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4265, new_AGEMA_signal_4264}) ) ;
    Precharger PrechargeCell_89 ( .D (plaintext_s1[38]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4261, new_AGEMA_signal_4260}) ) ;
    Precharger PrechargeCell_90 ( .D (plaintext_s1[37]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4257, new_AGEMA_signal_4256}) ) ;
    Precharger PrechargeCell_91 ( .D (plaintext_s1[36]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4253, new_AGEMA_signal_4252}) ) ;
    Precharger PrechargeCell_92 ( .D (plaintext_s1[35]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4249, new_AGEMA_signal_4248}) ) ;
    Precharger PrechargeCell_93 ( .D (plaintext_s1[34]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4245, new_AGEMA_signal_4244}) ) ;
    Precharger PrechargeCell_94 ( .D (plaintext_s1[33]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4241, new_AGEMA_signal_4240}) ) ;
    Precharger PrechargeCell_95 ( .D (plaintext_s1[32]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4237, new_AGEMA_signal_4236}) ) ;
    Precharger PrechargeCell_96 ( .D (plaintext_s1[31]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2819, new_AGEMA_signal_2818}) ) ;
    Precharger PrechargeCell_97 ( .D (plaintext_s1[30]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2813, new_AGEMA_signal_2812}) ) ;
    Precharger PrechargeCell_98 ( .D (plaintext_s1[29]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2807, new_AGEMA_signal_2806}) ) ;
    Precharger PrechargeCell_99 ( .D (plaintext_s1[28]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2801, new_AGEMA_signal_2800}) ) ;
    Precharger PrechargeCell_100 ( .D (plaintext_s1[27]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2795, new_AGEMA_signal_2794}) ) ;
    Precharger PrechargeCell_101 ( .D (plaintext_s1[26]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2789, new_AGEMA_signal_2788}) ) ;
    Precharger PrechargeCell_102 ( .D (plaintext_s1[25]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2783, new_AGEMA_signal_2782}) ) ;
    Precharger PrechargeCell_103 ( .D (plaintext_s1[24]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2777, new_AGEMA_signal_2776}) ) ;
    Precharger PrechargeCell_104 ( .D (plaintext_s1[23]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2867, new_AGEMA_signal_2866}) ) ;
    Precharger PrechargeCell_105 ( .D (plaintext_s1[22]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2861, new_AGEMA_signal_2860}) ) ;
    Precharger PrechargeCell_106 ( .D (plaintext_s1[21]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2855, new_AGEMA_signal_2854}) ) ;
    Precharger PrechargeCell_107 ( .D (plaintext_s1[20]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2849, new_AGEMA_signal_2848}) ) ;
    Precharger PrechargeCell_108 ( .D (plaintext_s1[19]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2843, new_AGEMA_signal_2842}) ) ;
    Precharger PrechargeCell_109 ( .D (plaintext_s1[18]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2837, new_AGEMA_signal_2836}) ) ;
    Precharger PrechargeCell_110 ( .D (plaintext_s1[17]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2831, new_AGEMA_signal_2830}) ) ;
    Precharger PrechargeCell_111 ( .D (plaintext_s1[16]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2825, new_AGEMA_signal_2824}) ) ;
    Precharger PrechargeCell_112 ( .D (plaintext_s1[15]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2917, new_AGEMA_signal_2916}) ) ;
    Precharger PrechargeCell_113 ( .D (plaintext_s1[14]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2911, new_AGEMA_signal_2910}) ) ;
    Precharger PrechargeCell_114 ( .D (plaintext_s1[13]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2905, new_AGEMA_signal_2904}) ) ;
    Precharger PrechargeCell_115 ( .D (plaintext_s1[12]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2899, new_AGEMA_signal_2898}) ) ;
    Precharger PrechargeCell_116 ( .D (plaintext_s1[11]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2893, new_AGEMA_signal_2892}) ) ;
    Precharger PrechargeCell_117 ( .D (plaintext_s1[10]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2887, new_AGEMA_signal_2886}) ) ;
    Precharger PrechargeCell_118 ( .D (plaintext_s1[9]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2881, new_AGEMA_signal_2880}) ) ;
    Precharger PrechargeCell_119 ( .D (plaintext_s1[8]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2875, new_AGEMA_signal_2874}) ) ;
    Precharger PrechargeCell_120 ( .D (plaintext_s1[7]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_5137, new_AGEMA_signal_5136}) ) ;
    Precharger PrechargeCell_121 ( .D (plaintext_s1[6]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_5133, new_AGEMA_signal_5132}) ) ;
    Precharger PrechargeCell_122 ( .D (plaintext_s1[5]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_5129, new_AGEMA_signal_5128}) ) ;
    Precharger PrechargeCell_123 ( .D (plaintext_s1[4]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_5125, new_AGEMA_signal_5124}) ) ;
    Precharger PrechargeCell_124 ( .D (plaintext_s1[3]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_5121, new_AGEMA_signal_5120}) ) ;
    Precharger PrechargeCell_125 ( .D (plaintext_s1[2]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_5117, new_AGEMA_signal_5116}) ) ;
    Precharger PrechargeCell_126 ( .D (plaintext_s1[1]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_5113, new_AGEMA_signal_5112}) ) ;
    Precharger PrechargeCell_127 ( .D (plaintext_s1[0]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_5091, new_AGEMA_signal_5090}) ) ;
    Precharger PrechargeCell_128 ( .D (key_s1[127]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4623, new_AGEMA_signal_4622}) ) ;
    Precharger PrechargeCell_129 ( .D (key_s1[126]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4619, new_AGEMA_signal_4618}) ) ;
    Precharger PrechargeCell_130 ( .D (key_s1[125]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4615, new_AGEMA_signal_4614}) ) ;
    Precharger PrechargeCell_131 ( .D (key_s1[124]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4611, new_AGEMA_signal_4610}) ) ;
    Precharger PrechargeCell_132 ( .D (key_s1[123]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4607, new_AGEMA_signal_4606}) ) ;
    Precharger PrechargeCell_133 ( .D (key_s1[122]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4603, new_AGEMA_signal_4602}) ) ;
    Precharger PrechargeCell_134 ( .D (key_s1[121]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4599, new_AGEMA_signal_4598}) ) ;
    Precharger PrechargeCell_135 ( .D (key_s1[120]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_4595, new_AGEMA_signal_4594}) ) ;
    Precharger PrechargeCell_136 ( .D (key_s1[119]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2967, new_AGEMA_signal_2966}) ) ;
    Precharger PrechargeCell_137 ( .D (key_s1[118]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2961, new_AGEMA_signal_2960}) ) ;
    Precharger PrechargeCell_138 ( .D (key_s1[117]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2955, new_AGEMA_signal_2954}) ) ;
    Precharger PrechargeCell_139 ( .D (key_s1[116]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2949, new_AGEMA_signal_2948}) ) ;
    Precharger PrechargeCell_140 ( .D (key_s1[115]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2943, new_AGEMA_signal_2942}) ) ;
    Precharger PrechargeCell_141 ( .D (key_s1[114]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2937, new_AGEMA_signal_2936}) ) ;
    Precharger PrechargeCell_142 ( .D (key_s1[113]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2931, new_AGEMA_signal_2930}) ) ;
    Precharger PrechargeCell_143 ( .D (key_s1[112]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2925, new_AGEMA_signal_2924}) ) ;
    Precharger PrechargeCell_144 ( .D (key_s1[111]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3017, new_AGEMA_signal_3016}) ) ;
    Precharger PrechargeCell_145 ( .D (key_s1[110]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3011, new_AGEMA_signal_3010}) ) ;
    Precharger PrechargeCell_146 ( .D (key_s1[109]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3005, new_AGEMA_signal_3004}) ) ;
    Precharger PrechargeCell_147 ( .D (key_s1[108]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2999, new_AGEMA_signal_2998}) ) ;
    Precharger PrechargeCell_148 ( .D (key_s1[107]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2993, new_AGEMA_signal_2992}) ) ;
    Precharger PrechargeCell_149 ( .D (key_s1[106]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2987, new_AGEMA_signal_2986}) ) ;
    Precharger PrechargeCell_150 ( .D (key_s1[105]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2981, new_AGEMA_signal_2980}) ) ;
    Precharger PrechargeCell_151 ( .D (key_s1[104]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_2975, new_AGEMA_signal_2974}) ) ;
    Precharger PrechargeCell_152 ( .D (key_s1[103]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3065, new_AGEMA_signal_3064}) ) ;
    Precharger PrechargeCell_153 ( .D (key_s1[102]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3059, new_AGEMA_signal_3058}) ) ;
    Precharger PrechargeCell_154 ( .D (key_s1[101]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3053, new_AGEMA_signal_3052}) ) ;
    Precharger PrechargeCell_155 ( .D (key_s1[100]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3047, new_AGEMA_signal_3046}) ) ;
    Precharger PrechargeCell_156 ( .D (key_s1[99]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3041, new_AGEMA_signal_3040}) ) ;
    Precharger PrechargeCell_157 ( .D (key_s1[98]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3035, new_AGEMA_signal_3034}) ) ;
    Precharger PrechargeCell_158 ( .D (key_s1[97]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3029, new_AGEMA_signal_3028}) ) ;
    Precharger PrechargeCell_159 ( .D (key_s1[96]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3023, new_AGEMA_signal_3022}) ) ;
    Precharger PrechargeCell_160 ( .D (key_s1[95]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3115, new_AGEMA_signal_3114}) ) ;
    Precharger PrechargeCell_161 ( .D (key_s1[94]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3109, new_AGEMA_signal_3108}) ) ;
    Precharger PrechargeCell_162 ( .D (key_s1[93]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3103, new_AGEMA_signal_3102}) ) ;
    Precharger PrechargeCell_163 ( .D (key_s1[92]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3097, new_AGEMA_signal_3096}) ) ;
    Precharger PrechargeCell_164 ( .D (key_s1[91]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3091, new_AGEMA_signal_3090}) ) ;
    Precharger PrechargeCell_165 ( .D (key_s1[90]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3085, new_AGEMA_signal_3084}) ) ;
    Precharger PrechargeCell_166 ( .D (key_s1[89]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3079, new_AGEMA_signal_3078}) ) ;
    Precharger PrechargeCell_167 ( .D (key_s1[88]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3073, new_AGEMA_signal_3072}) ) ;
    Precharger PrechargeCell_168 ( .D (key_s1[87]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3163, new_AGEMA_signal_3162}) ) ;
    Precharger PrechargeCell_169 ( .D (key_s1[86]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3157, new_AGEMA_signal_3156}) ) ;
    Precharger PrechargeCell_170 ( .D (key_s1[85]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3151, new_AGEMA_signal_3150}) ) ;
    Precharger PrechargeCell_171 ( .D (key_s1[84]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3145, new_AGEMA_signal_3144}) ) ;
    Precharger PrechargeCell_172 ( .D (key_s1[83]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3139, new_AGEMA_signal_3138}) ) ;
    Precharger PrechargeCell_173 ( .D (key_s1[82]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3133, new_AGEMA_signal_3132}) ) ;
    Precharger PrechargeCell_174 ( .D (key_s1[81]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3127, new_AGEMA_signal_3126}) ) ;
    Precharger PrechargeCell_175 ( .D (key_s1[80]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3121, new_AGEMA_signal_3120}) ) ;
    Precharger PrechargeCell_176 ( .D (key_s1[79]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3213, new_AGEMA_signal_3212}) ) ;
    Precharger PrechargeCell_177 ( .D (key_s1[78]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3207, new_AGEMA_signal_3206}) ) ;
    Precharger PrechargeCell_178 ( .D (key_s1[77]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3201, new_AGEMA_signal_3200}) ) ;
    Precharger PrechargeCell_179 ( .D (key_s1[76]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3195, new_AGEMA_signal_3194}) ) ;
    Precharger PrechargeCell_180 ( .D (key_s1[75]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3189, new_AGEMA_signal_3188}) ) ;
    Precharger PrechargeCell_181 ( .D (key_s1[74]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3183, new_AGEMA_signal_3182}) ) ;
    Precharger PrechargeCell_182 ( .D (key_s1[73]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3177, new_AGEMA_signal_3176}) ) ;
    Precharger PrechargeCell_183 ( .D (key_s1[72]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3171, new_AGEMA_signal_3170}) ) ;
    Precharger PrechargeCell_184 ( .D (key_s1[71]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3261, new_AGEMA_signal_3260}) ) ;
    Precharger PrechargeCell_185 ( .D (key_s1[70]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3255, new_AGEMA_signal_3254}) ) ;
    Precharger PrechargeCell_186 ( .D (key_s1[69]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3249, new_AGEMA_signal_3248}) ) ;
    Precharger PrechargeCell_187 ( .D (key_s1[68]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3243, new_AGEMA_signal_3242}) ) ;
    Precharger PrechargeCell_188 ( .D (key_s1[67]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3237, new_AGEMA_signal_3236}) ) ;
    Precharger PrechargeCell_189 ( .D (key_s1[66]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3231, new_AGEMA_signal_3230}) ) ;
    Precharger PrechargeCell_190 ( .D (key_s1[65]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3225, new_AGEMA_signal_3224}) ) ;
    Precharger PrechargeCell_191 ( .D (key_s1[64]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3219, new_AGEMA_signal_3218}) ) ;
    Precharger PrechargeCell_192 ( .D (key_s1[63]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3311, new_AGEMA_signal_3310}) ) ;
    Precharger PrechargeCell_193 ( .D (key_s1[62]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3305, new_AGEMA_signal_3304}) ) ;
    Precharger PrechargeCell_194 ( .D (key_s1[61]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3299, new_AGEMA_signal_3298}) ) ;
    Precharger PrechargeCell_195 ( .D (key_s1[60]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3293, new_AGEMA_signal_3292}) ) ;
    Precharger PrechargeCell_196 ( .D (key_s1[59]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3287, new_AGEMA_signal_3286}) ) ;
    Precharger PrechargeCell_197 ( .D (key_s1[58]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3281, new_AGEMA_signal_3280}) ) ;
    Precharger PrechargeCell_198 ( .D (key_s1[57]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3275, new_AGEMA_signal_3274}) ) ;
    Precharger PrechargeCell_199 ( .D (key_s1[56]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3269, new_AGEMA_signal_3268}) ) ;
    Precharger PrechargeCell_200 ( .D (key_s1[55]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3359, new_AGEMA_signal_3358}) ) ;
    Precharger PrechargeCell_201 ( .D (key_s1[54]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3353, new_AGEMA_signal_3352}) ) ;
    Precharger PrechargeCell_202 ( .D (key_s1[53]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3347, new_AGEMA_signal_3346}) ) ;
    Precharger PrechargeCell_203 ( .D (key_s1[52]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3341, new_AGEMA_signal_3340}) ) ;
    Precharger PrechargeCell_204 ( .D (key_s1[51]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3335, new_AGEMA_signal_3334}) ) ;
    Precharger PrechargeCell_205 ( .D (key_s1[50]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3329, new_AGEMA_signal_3328}) ) ;
    Precharger PrechargeCell_206 ( .D (key_s1[49]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3323, new_AGEMA_signal_3322}) ) ;
    Precharger PrechargeCell_207 ( .D (key_s1[48]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3317, new_AGEMA_signal_3316}) ) ;
    Precharger PrechargeCell_208 ( .D (key_s1[47]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3409, new_AGEMA_signal_3408}) ) ;
    Precharger PrechargeCell_209 ( .D (key_s1[46]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3403, new_AGEMA_signal_3402}) ) ;
    Precharger PrechargeCell_210 ( .D (key_s1[45]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3397, new_AGEMA_signal_3396}) ) ;
    Precharger PrechargeCell_211 ( .D (key_s1[44]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3391, new_AGEMA_signal_3390}) ) ;
    Precharger PrechargeCell_212 ( .D (key_s1[43]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3385, new_AGEMA_signal_3384}) ) ;
    Precharger PrechargeCell_213 ( .D (key_s1[42]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3379, new_AGEMA_signal_3378}) ) ;
    Precharger PrechargeCell_214 ( .D (key_s1[41]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3373, new_AGEMA_signal_3372}) ) ;
    Precharger PrechargeCell_215 ( .D (key_s1[40]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3367, new_AGEMA_signal_3366}) ) ;
    Precharger PrechargeCell_216 ( .D (key_s1[39]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3457, new_AGEMA_signal_3456}) ) ;
    Precharger PrechargeCell_217 ( .D (key_s1[38]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3451, new_AGEMA_signal_3450}) ) ;
    Precharger PrechargeCell_218 ( .D (key_s1[37]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3445, new_AGEMA_signal_3444}) ) ;
    Precharger PrechargeCell_219 ( .D (key_s1[36]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3439, new_AGEMA_signal_3438}) ) ;
    Precharger PrechargeCell_220 ( .D (key_s1[35]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3433, new_AGEMA_signal_3432}) ) ;
    Precharger PrechargeCell_221 ( .D (key_s1[34]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3427, new_AGEMA_signal_3426}) ) ;
    Precharger PrechargeCell_222 ( .D (key_s1[33]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3421, new_AGEMA_signal_3420}) ) ;
    Precharger PrechargeCell_223 ( .D (key_s1[32]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3415, new_AGEMA_signal_3414}) ) ;
    Precharger PrechargeCell_224 ( .D (key_s1[31]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3507, new_AGEMA_signal_3506}) ) ;
    Precharger PrechargeCell_225 ( .D (key_s1[30]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3501, new_AGEMA_signal_3500}) ) ;
    Precharger PrechargeCell_226 ( .D (key_s1[29]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3495, new_AGEMA_signal_3494}) ) ;
    Precharger PrechargeCell_227 ( .D (key_s1[28]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3489, new_AGEMA_signal_3488}) ) ;
    Precharger PrechargeCell_228 ( .D (key_s1[27]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3483, new_AGEMA_signal_3482}) ) ;
    Precharger PrechargeCell_229 ( .D (key_s1[26]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3477, new_AGEMA_signal_3476}) ) ;
    Precharger PrechargeCell_230 ( .D (key_s1[25]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3471, new_AGEMA_signal_3470}) ) ;
    Precharger PrechargeCell_231 ( .D (key_s1[24]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3465, new_AGEMA_signal_3464}) ) ;
    Precharger PrechargeCell_232 ( .D (key_s1[23]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3555, new_AGEMA_signal_3554}) ) ;
    Precharger PrechargeCell_233 ( .D (key_s1[22]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3549, new_AGEMA_signal_3548}) ) ;
    Precharger PrechargeCell_234 ( .D (key_s1[21]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3543, new_AGEMA_signal_3542}) ) ;
    Precharger PrechargeCell_235 ( .D (key_s1[20]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3537, new_AGEMA_signal_3536}) ) ;
    Precharger PrechargeCell_236 ( .D (key_s1[19]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3531, new_AGEMA_signal_3530}) ) ;
    Precharger PrechargeCell_237 ( .D (key_s1[18]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3525, new_AGEMA_signal_3524}) ) ;
    Precharger PrechargeCell_238 ( .D (key_s1[17]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3519, new_AGEMA_signal_3518}) ) ;
    Precharger PrechargeCell_239 ( .D (key_s1[16]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3513, new_AGEMA_signal_3512}) ) ;
    Precharger PrechargeCell_240 ( .D (key_s1[15]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3605, new_AGEMA_signal_3604}) ) ;
    Precharger PrechargeCell_241 ( .D (key_s1[14]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3599, new_AGEMA_signal_3598}) ) ;
    Precharger PrechargeCell_242 ( .D (key_s1[13]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3593, new_AGEMA_signal_3592}) ) ;
    Precharger PrechargeCell_243 ( .D (key_s1[12]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3587, new_AGEMA_signal_3586}) ) ;
    Precharger PrechargeCell_244 ( .D (key_s1[11]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3581, new_AGEMA_signal_3580}) ) ;
    Precharger PrechargeCell_245 ( .D (key_s1[10]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3575, new_AGEMA_signal_3574}) ) ;
    Precharger PrechargeCell_246 ( .D (key_s1[9]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3569, new_AGEMA_signal_3568}) ) ;
    Precharger PrechargeCell_247 ( .D (key_s1[8]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3563, new_AGEMA_signal_3562}) ) ;
    Precharger PrechargeCell_248 ( .D (key_s1[7]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3639, new_AGEMA_signal_3638}) ) ;
    Precharger PrechargeCell_249 ( .D (key_s1[6]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3635, new_AGEMA_signal_3634}) ) ;
    Precharger PrechargeCell_250 ( .D (key_s1[5]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3631, new_AGEMA_signal_3630}) ) ;
    Precharger PrechargeCell_251 ( .D (key_s1[4]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3627, new_AGEMA_signal_3626}) ) ;
    Precharger PrechargeCell_252 ( .D (key_s1[3]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3623, new_AGEMA_signal_3622}) ) ;
    Precharger PrechargeCell_253 ( .D (key_s1[2]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3619, new_AGEMA_signal_3618}) ) ;
    Precharger PrechargeCell_254 ( .D (key_s1[1]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3615, new_AGEMA_signal_3614}) ) ;
    Precharger PrechargeCell_255 ( .D (key_s1[0]), .pre (LMDPL_pre2), .Q ({new_AGEMA_signal_3611, new_AGEMA_signal_3610}) ) ;

    /* register cells */
    reg_sr_LMDPL ctrl_seq6_SFF_0_Q_reg_FF_FF ( .D (ctrl_seq6_SFF_0_QD), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (ctrl_seq6In_1_), .QN () ) ;
    reg_sr_LMDPL ctrl_seq6_SFF_1_Q_reg_FF_FF ( .D (ctrl_seq6_SFF_1_QD), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (ctrl_seq6In_2_), .QN () ) ;
    reg_sr_LMDPL ctrl_seq6_SFF_2_Q_reg_FF_FF ( .D (ctrl_seq6_SFF_2_QD), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (ctrl_seq6In_3_), .QN () ) ;
    reg_sr_LMDPL ctrl_seq6_SFF_3_Q_reg_FF_FF ( .D (ctrl_seq6_SFF_3_QD), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (ctrl_seq6In_4_), .QN () ) ;
    reg_sr_LMDPL ctrl_seq6_SFF_4_Q_reg_FF_FF ( .D (ctrl_seq6_SFF_4_QD), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (ctrl_seq6Out_4_), .QN () ) ;
    reg_sr_LMDPL ctrl_seq4_SFF_0_Q_reg_FF_FF ( .D (ctrl_seq4_SFF_0_QD), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (ctrl_seq4In_1_), .QN () ) ;
    reg_sr_LMDPL ctrl_seq4_SFF_1_Q_reg_FF_FF ( .D (ctrl_seq4_SFF_1_QD), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (ctrl_seq4Out_1_), .QN () ) ;
    reg_sr_LMDPL ctrl_CSselMC_reg_FF_FF ( .D (ctrl_N14), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (ctrl_n6), .QN () ) ;
    reg_sr_LMDPL ctrl_CSenRC_reg_FF_FF ( .D (selSR), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (enRCon), .QN () ) ;
    reg_LMDPL stateArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4341, new_AGEMA_signal_4340, stateArray_S00reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1987, ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_LMDPL stateArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4343, new_AGEMA_signal_4342, stateArray_S00reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1993, ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_LMDPL stateArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4345, new_AGEMA_signal_4344, stateArray_S00reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1999, ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_LMDPL stateArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4347, new_AGEMA_signal_4346, stateArray_S00reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2005, ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_LMDPL stateArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4349, new_AGEMA_signal_4348, stateArray_S00reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2011, ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_LMDPL stateArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4351, new_AGEMA_signal_4350, stateArray_S00reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2017, ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_LMDPL stateArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4353, new_AGEMA_signal_4352, stateArray_S00reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2023, ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_LMDPL stateArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4355, new_AGEMA_signal_4354, stateArray_S00reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2029, ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_LMDPL stateArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4357, new_AGEMA_signal_4356, stateArray_S01reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2335, ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_LMDPL stateArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4359, new_AGEMA_signal_4358, stateArray_S01reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2341, ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_LMDPL stateArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4361, new_AGEMA_signal_4360, stateArray_S01reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2347, ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_LMDPL stateArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4363, new_AGEMA_signal_4362, stateArray_S01reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2353, ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_LMDPL stateArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4365, new_AGEMA_signal_4364, stateArray_S01reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2359, ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_LMDPL stateArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4367, new_AGEMA_signal_4366, stateArray_S01reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2365, ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_LMDPL stateArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4369, new_AGEMA_signal_4368, stateArray_S01reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2371, ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_LMDPL stateArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4371, new_AGEMA_signal_4370, stateArray_S01reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2377, ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_LMDPL stateArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4375, new_AGEMA_signal_4374, stateArray_S02reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2383, ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_LMDPL stateArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4377, new_AGEMA_signal_4376, stateArray_S02reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2389, ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_LMDPL stateArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4379, new_AGEMA_signal_4378, stateArray_S02reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2395, ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_LMDPL stateArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4381, new_AGEMA_signal_4380, stateArray_S02reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2401, ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_LMDPL stateArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4383, new_AGEMA_signal_4382, stateArray_S02reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2407, ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_LMDPL stateArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4385, new_AGEMA_signal_4384, stateArray_S02reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2413, ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_LMDPL stateArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4387, new_AGEMA_signal_4386, stateArray_S02reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2419, ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_LMDPL stateArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4389, new_AGEMA_signal_4388, stateArray_S02reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2425, ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_LMDPL stateArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4391, new_AGEMA_signal_4390, stateArray_S03reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2433, ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_LMDPL stateArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4393, new_AGEMA_signal_4392, stateArray_S03reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2439, ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_LMDPL stateArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4395, new_AGEMA_signal_4394, stateArray_S03reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2445, ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_LMDPL stateArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4397, new_AGEMA_signal_4396, stateArray_S03reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2451, ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_LMDPL stateArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4399, new_AGEMA_signal_4398, stateArray_S03reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2457, ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_LMDPL stateArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4401, new_AGEMA_signal_4400, stateArray_S03reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2463, ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_LMDPL stateArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4403, new_AGEMA_signal_4402, stateArray_S03reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2469, ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_LMDPL stateArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4405, new_AGEMA_signal_4404, stateArray_S03reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2475, ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_LMDPL stateArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4409, new_AGEMA_signal_4408, stateArray_S10reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2141, ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_LMDPL stateArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4411, new_AGEMA_signal_4410, stateArray_S10reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2137, ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_LMDPL stateArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4413, new_AGEMA_signal_4412, stateArray_S10reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2135, ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_LMDPL stateArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4415, new_AGEMA_signal_4414, stateArray_S10reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2145, ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_LMDPL stateArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4417, new_AGEMA_signal_4416, stateArray_S10reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2131, ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_LMDPL stateArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4419, new_AGEMA_signal_4418, stateArray_S10reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2127, ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_LMDPL stateArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4421, new_AGEMA_signal_4420, stateArray_S10reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2123, ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_LMDPL stateArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4423, new_AGEMA_signal_4422, stateArray_S10reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2121, ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_LMDPL stateArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4425, new_AGEMA_signal_4424, stateArray_S11reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2483, ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_LMDPL stateArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4427, new_AGEMA_signal_4426, stateArray_S11reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2489, ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_LMDPL stateArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4429, new_AGEMA_signal_4428, stateArray_S11reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2495, ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_LMDPL stateArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4431, new_AGEMA_signal_4430, stateArray_S11reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2501, ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_LMDPL stateArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4433, new_AGEMA_signal_4432, stateArray_S11reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2507, ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_LMDPL stateArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4435, new_AGEMA_signal_4434, stateArray_S11reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2513, ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_LMDPL stateArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4437, new_AGEMA_signal_4436, stateArray_S11reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2519, ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_LMDPL stateArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4439, new_AGEMA_signal_4438, stateArray_S11reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2525, ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_LMDPL stateArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4443, new_AGEMA_signal_4442, stateArray_S12reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2531, ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_LMDPL stateArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4445, new_AGEMA_signal_4444, stateArray_S12reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2537, ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_LMDPL stateArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4447, new_AGEMA_signal_4446, stateArray_S12reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2543, ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_LMDPL stateArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4449, new_AGEMA_signal_4448, stateArray_S12reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2549, ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_LMDPL stateArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4451, new_AGEMA_signal_4450, stateArray_S12reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2555, ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_LMDPL stateArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4453, new_AGEMA_signal_4452, stateArray_S12reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2561, ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_LMDPL stateArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4455, new_AGEMA_signal_4454, stateArray_S12reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2567, ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_LMDPL stateArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4457, new_AGEMA_signal_4456, stateArray_S12reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2573, ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_LMDPL stateArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4459, new_AGEMA_signal_4458, stateArray_S13reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2581, ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_LMDPL stateArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4461, new_AGEMA_signal_4460, stateArray_S13reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2587, ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_LMDPL stateArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4463, new_AGEMA_signal_4462, stateArray_S13reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2593, ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_LMDPL stateArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4465, new_AGEMA_signal_4464, stateArray_S13reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2599, ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_LMDPL stateArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4467, new_AGEMA_signal_4466, stateArray_S13reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2605, ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_LMDPL stateArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4469, new_AGEMA_signal_4468, stateArray_S13reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2611, ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_LMDPL stateArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4471, new_AGEMA_signal_4470, stateArray_S13reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2617, ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_LMDPL stateArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4473, new_AGEMA_signal_4472, stateArray_S13reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2623, ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_LMDPL stateArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4477, new_AGEMA_signal_4476, stateArray_S20reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2111, ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_LMDPL stateArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4479, new_AGEMA_signal_4478, stateArray_S20reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2105, ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_LMDPL stateArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4481, new_AGEMA_signal_4480, stateArray_S20reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2097, ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_LMDPL stateArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4483, new_AGEMA_signal_4482, stateArray_S20reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2091, ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_LMDPL stateArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4485, new_AGEMA_signal_4484, stateArray_S20reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2085, ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_LMDPL stateArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4487, new_AGEMA_signal_4486, stateArray_S20reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2079, ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_LMDPL stateArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4489, new_AGEMA_signal_4488, stateArray_S20reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2073, ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_LMDPL stateArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4491, new_AGEMA_signal_4490, stateArray_S20reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2067, ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_LMDPL stateArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4493, new_AGEMA_signal_4492, stateArray_S21reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2631, ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_LMDPL stateArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4495, new_AGEMA_signal_4494, stateArray_S21reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2637, ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_LMDPL stateArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4497, new_AGEMA_signal_4496, stateArray_S21reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2643, ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_LMDPL stateArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4499, new_AGEMA_signal_4498, stateArray_S21reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2649, ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_LMDPL stateArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4501, new_AGEMA_signal_4500, stateArray_S21reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2655, ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_LMDPL stateArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4503, new_AGEMA_signal_4502, stateArray_S21reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2661, ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_LMDPL stateArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4505, new_AGEMA_signal_4504, stateArray_S21reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2667, ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_LMDPL stateArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4507, new_AGEMA_signal_4506, stateArray_S21reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2673, ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_LMDPL stateArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4511, new_AGEMA_signal_4510, stateArray_S22reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2679, ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_LMDPL stateArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4513, new_AGEMA_signal_4512, stateArray_S22reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2685, ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_LMDPL stateArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4515, new_AGEMA_signal_4514, stateArray_S22reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2691, ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_LMDPL stateArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4517, new_AGEMA_signal_4516, stateArray_S22reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2697, ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_LMDPL stateArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4519, new_AGEMA_signal_4518, stateArray_S22reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2703, ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_LMDPL stateArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4521, new_AGEMA_signal_4520, stateArray_S22reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2709, ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_LMDPL stateArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4523, new_AGEMA_signal_4522, stateArray_S22reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2715, ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_LMDPL stateArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4525, new_AGEMA_signal_4524, stateArray_S22reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2721, ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_LMDPL stateArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4527, new_AGEMA_signal_4526, stateArray_S23reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2729, ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_LMDPL stateArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4529, new_AGEMA_signal_4528, stateArray_S23reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2735, ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_LMDPL stateArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4531, new_AGEMA_signal_4530, stateArray_S23reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2741, ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_LMDPL stateArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4533, new_AGEMA_signal_4532, stateArray_S23reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2747, ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_LMDPL stateArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4535, new_AGEMA_signal_4534, stateArray_S23reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2753, ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_LMDPL stateArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4537, new_AGEMA_signal_4536, stateArray_S23reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2759, ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_LMDPL stateArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4539, new_AGEMA_signal_4538, stateArray_S23reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2765, ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_LMDPL stateArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4541, new_AGEMA_signal_4540, stateArray_S23reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2771, ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_LMDPL stateArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4545, new_AGEMA_signal_4544, stateArray_S30reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2109, ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_LMDPL stateArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4547, new_AGEMA_signal_4546, stateArray_S30reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2103, ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_LMDPL stateArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4549, new_AGEMA_signal_4548, stateArray_S30reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2099, ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_LMDPL stateArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4551, new_AGEMA_signal_4550, stateArray_S30reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2093, ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_LMDPL stateArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4553, new_AGEMA_signal_4552, stateArray_S30reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2087, ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_LMDPL stateArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4555, new_AGEMA_signal_4554, stateArray_S30reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2081, ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_LMDPL stateArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4557, new_AGEMA_signal_4556, stateArray_S30reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2075, ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_LMDPL stateArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4559, new_AGEMA_signal_4558, stateArray_S30reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2069, ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_LMDPL stateArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4561, new_AGEMA_signal_4560, stateArray_S31reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2779, ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_LMDPL stateArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4563, new_AGEMA_signal_4562, stateArray_S31reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2785, ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_LMDPL stateArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4565, new_AGEMA_signal_4564, stateArray_S31reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2791, ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_LMDPL stateArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4567, new_AGEMA_signal_4566, stateArray_S31reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2797, ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_LMDPL stateArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4569, new_AGEMA_signal_4568, stateArray_S31reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2803, ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_LMDPL stateArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4571, new_AGEMA_signal_4570, stateArray_S31reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2809, ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_LMDPL stateArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4573, new_AGEMA_signal_4572, stateArray_S31reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2815, ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_LMDPL stateArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4575, new_AGEMA_signal_4574, stateArray_S31reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2821, ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_LMDPL stateArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4579, new_AGEMA_signal_4578, stateArray_S32reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2827, ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_LMDPL stateArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4581, new_AGEMA_signal_4580, stateArray_S32reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2833, ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_LMDPL stateArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4583, new_AGEMA_signal_4582, stateArray_S32reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2839, ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_LMDPL stateArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4585, new_AGEMA_signal_4584, stateArray_S32reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2845, ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_LMDPL stateArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4587, new_AGEMA_signal_4586, stateArray_S32reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2851, ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_LMDPL stateArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4589, new_AGEMA_signal_4588, stateArray_S32reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2857, ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_LMDPL stateArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4591, new_AGEMA_signal_4590, stateArray_S32reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2863, ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_LMDPL stateArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4593, new_AGEMA_signal_4592, stateArray_S32reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2869, ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_LMDPL stateArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5111, new_AGEMA_signal_5110, stateArray_S33reg_gff_1_SFF_0_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2877, ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_LMDPL stateArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5157, new_AGEMA_signal_5156, stateArray_S33reg_gff_1_SFF_1_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2883, ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_LMDPL stateArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5159, new_AGEMA_signal_5158, stateArray_S33reg_gff_1_SFF_2_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2889, ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_LMDPL stateArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5161, new_AGEMA_signal_5160, stateArray_S33reg_gff_1_SFF_3_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2895, ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_LMDPL stateArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5163, new_AGEMA_signal_5162, stateArray_S33reg_gff_1_SFF_4_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2901, ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_LMDPL stateArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5165, new_AGEMA_signal_5164, stateArray_S33reg_gff_1_SFF_5_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2907, ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_LMDPL stateArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5167, new_AGEMA_signal_5166, stateArray_S33reg_gff_1_SFF_6_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2913, ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_LMDPL stateArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5169, new_AGEMA_signal_5168, stateArray_S33reg_gff_1_SFF_7_QD}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2919, ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_LMDPL KeyArray_S00reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4867, new_AGEMA_signal_4866, KeyArray_S00reg_gff_1_SFF_0_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1989, new_AGEMA_signal_1988, keyStateIn[0]}) ) ;
    reg_LMDPL KeyArray_S00reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4869, new_AGEMA_signal_4868, KeyArray_S00reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_1995, new_AGEMA_signal_1994, keyStateIn[1]}) ) ;
    reg_LMDPL KeyArray_S00reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4871, new_AGEMA_signal_4870, KeyArray_S00reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2001, new_AGEMA_signal_2000, keyStateIn[2]}) ) ;
    reg_LMDPL KeyArray_S00reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4873, new_AGEMA_signal_4872, KeyArray_S00reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2007, new_AGEMA_signal_2006, keyStateIn[3]}) ) ;
    reg_LMDPL KeyArray_S00reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4875, new_AGEMA_signal_4874, KeyArray_S00reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2013, new_AGEMA_signal_2012, keyStateIn[4]}) ) ;
    reg_LMDPL KeyArray_S00reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4877, new_AGEMA_signal_4876, KeyArray_S00reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2019, new_AGEMA_signal_2018, keyStateIn[5]}) ) ;
    reg_LMDPL KeyArray_S00reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4879, new_AGEMA_signal_4878, KeyArray_S00reg_gff_1_SFF_6_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2025, new_AGEMA_signal_2024, keyStateIn[6]}) ) ;
    reg_LMDPL KeyArray_S00reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4881, new_AGEMA_signal_4880, KeyArray_S00reg_gff_1_SFF_7_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2031, new_AGEMA_signal_2030, keyStateIn[7]}) ) ;
    reg_LMDPL KeyArray_S01reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4655, new_AGEMA_signal_4654, KeyArray_S01reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2063, new_AGEMA_signal_2062, KeyArray_outS01ser_0_}) ) ;
    reg_LMDPL KeyArray_S01reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4657, new_AGEMA_signal_4656, KeyArray_S01reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2059, new_AGEMA_signal_2058, KeyArray_outS01ser_1_}) ) ;
    reg_LMDPL KeyArray_S01reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4659, new_AGEMA_signal_4658, KeyArray_S01reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2055, new_AGEMA_signal_2054, KeyArray_outS01ser_2_}) ) ;
    reg_LMDPL KeyArray_S01reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4661, new_AGEMA_signal_4660, KeyArray_S01reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2051, new_AGEMA_signal_2050, KeyArray_outS01ser_3_}) ) ;
    reg_LMDPL KeyArray_S01reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4663, new_AGEMA_signal_4662, KeyArray_S01reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2047, new_AGEMA_signal_2046, KeyArray_outS01ser_4_}) ) ;
    reg_LMDPL KeyArray_S01reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4665, new_AGEMA_signal_4664, KeyArray_S01reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2043, new_AGEMA_signal_2042, KeyArray_outS01ser_5_}) ) ;
    reg_LMDPL KeyArray_S01reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4667, new_AGEMA_signal_4666, KeyArray_S01reg_gff_1_SFF_6_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2039, new_AGEMA_signal_2038, KeyArray_outS01ser_6_}) ) ;
    reg_LMDPL KeyArray_S01reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4669, new_AGEMA_signal_4668, KeyArray_S01reg_gff_1_SFF_7_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2035, new_AGEMA_signal_2034, KeyArray_outS01ser_7_}) ) ;
    reg_LMDPL KeyArray_S02reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4673, new_AGEMA_signal_4672, KeyArray_S02reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2927, new_AGEMA_signal_2926, KeyArray_outS02ser[0]}) ) ;
    reg_LMDPL KeyArray_S02reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4675, new_AGEMA_signal_4674, KeyArray_S02reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2933, new_AGEMA_signal_2932, KeyArray_outS02ser[1]}) ) ;
    reg_LMDPL KeyArray_S02reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4677, new_AGEMA_signal_4676, KeyArray_S02reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2939, new_AGEMA_signal_2938, KeyArray_outS02ser[2]}) ) ;
    reg_LMDPL KeyArray_S02reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4679, new_AGEMA_signal_4678, KeyArray_S02reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2945, new_AGEMA_signal_2944, KeyArray_outS02ser[3]}) ) ;
    reg_LMDPL KeyArray_S02reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4681, new_AGEMA_signal_4680, KeyArray_S02reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2951, new_AGEMA_signal_2950, KeyArray_outS02ser[4]}) ) ;
    reg_LMDPL KeyArray_S02reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4683, new_AGEMA_signal_4682, KeyArray_S02reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2957, new_AGEMA_signal_2956, KeyArray_outS02ser[5]}) ) ;
    reg_LMDPL KeyArray_S02reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4685, new_AGEMA_signal_4684, KeyArray_S02reg_gff_1_SFF_6_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2963, new_AGEMA_signal_2962, KeyArray_outS02ser[6]}) ) ;
    reg_LMDPL KeyArray_S02reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4687, new_AGEMA_signal_4686, KeyArray_S02reg_gff_1_SFF_7_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2969, new_AGEMA_signal_2968, KeyArray_outS02ser[7]}) ) ;
    reg_LMDPL KeyArray_S03reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4689, new_AGEMA_signal_4688, KeyArray_S03reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2977, new_AGEMA_signal_2976, KeyArray_outS03ser[0]}) ) ;
    reg_LMDPL KeyArray_S03reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4691, new_AGEMA_signal_4690, KeyArray_S03reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2983, new_AGEMA_signal_2982, KeyArray_outS03ser[1]}) ) ;
    reg_LMDPL KeyArray_S03reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4693, new_AGEMA_signal_4692, KeyArray_S03reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2989, new_AGEMA_signal_2988, KeyArray_outS03ser[2]}) ) ;
    reg_LMDPL KeyArray_S03reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4695, new_AGEMA_signal_4694, KeyArray_S03reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_2995, new_AGEMA_signal_2994, KeyArray_outS03ser[3]}) ) ;
    reg_LMDPL KeyArray_S03reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4697, new_AGEMA_signal_4696, KeyArray_S03reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3001, new_AGEMA_signal_3000, KeyArray_outS03ser[4]}) ) ;
    reg_LMDPL KeyArray_S03reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4699, new_AGEMA_signal_4698, KeyArray_S03reg_gff_1_SFF_5_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3007, new_AGEMA_signal_3006, KeyArray_outS03ser[5]}) ) ;
    reg_LMDPL KeyArray_S03reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4701, new_AGEMA_signal_4700, KeyArray_S03reg_gff_1_SFF_6_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3013, new_AGEMA_signal_3012, KeyArray_outS03ser[6]}) ) ;
    reg_LMDPL KeyArray_S03reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4703, new_AGEMA_signal_4702, KeyArray_S03reg_gff_1_SFF_7_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3019, new_AGEMA_signal_3018, KeyArray_outS03ser[7]}) ) ;
    reg_LMDPL KeyArray_S10reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4707, new_AGEMA_signal_4706, KeyArray_S10reg_gff_1_SFF_0_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3025, new_AGEMA_signal_3024, KeyArray_outS10ser[0]}) ) ;
    reg_LMDPL KeyArray_S10reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4709, new_AGEMA_signal_4708, KeyArray_S10reg_gff_1_SFF_1_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3031, new_AGEMA_signal_3030, KeyArray_outS10ser[1]}) ) ;
    reg_LMDPL KeyArray_S10reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4711, new_AGEMA_signal_4710, KeyArray_S10reg_gff_1_SFF_2_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3037, new_AGEMA_signal_3036, KeyArray_outS10ser[2]}) ) ;
    reg_LMDPL KeyArray_S10reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4713, new_AGEMA_signal_4712, KeyArray_S10reg_gff_1_SFF_3_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3043, new_AGEMA_signal_3042, KeyArray_outS10ser[3]}) ) ;
    reg_LMDPL KeyArray_S10reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4715, new_AGEMA_signal_4714, KeyArray_S10reg_gff_1_SFF_4_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3049, new_AGEMA_signal_3048, KeyArray_outS10ser[4]}) ) ;
    reg_LMDPL KeyArray_S10reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4717, new_AGEMA_signal_4716, KeyArray_S10reg_gff_1_SFF_5_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3055, new_AGEMA_signal_3054, KeyArray_outS10ser[5]}) ) ;
    reg_LMDPL KeyArray_S10reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4719, new_AGEMA_signal_4718, KeyArray_S10reg_gff_1_SFF_6_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3061, new_AGEMA_signal_3060, KeyArray_outS10ser[6]}) ) ;
    reg_LMDPL KeyArray_S10reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4721, new_AGEMA_signal_4720, KeyArray_S10reg_gff_1_SFF_7_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3067, new_AGEMA_signal_3066, KeyArray_outS10ser[7]}) ) ;
    reg_LMDPL KeyArray_S11reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4723, new_AGEMA_signal_4722, KeyArray_S11reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3075, new_AGEMA_signal_3074, KeyArray_outS11ser[0]}) ) ;
    reg_LMDPL KeyArray_S11reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4725, new_AGEMA_signal_4724, KeyArray_S11reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3081, new_AGEMA_signal_3080, KeyArray_outS11ser[1]}) ) ;
    reg_LMDPL KeyArray_S11reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4727, new_AGEMA_signal_4726, KeyArray_S11reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3087, new_AGEMA_signal_3086, KeyArray_outS11ser[2]}) ) ;
    reg_LMDPL KeyArray_S11reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4729, new_AGEMA_signal_4728, KeyArray_S11reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3093, new_AGEMA_signal_3092, KeyArray_outS11ser[3]}) ) ;
    reg_LMDPL KeyArray_S11reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4731, new_AGEMA_signal_4730, KeyArray_S11reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3099, new_AGEMA_signal_3098, KeyArray_outS11ser[4]}) ) ;
    reg_LMDPL KeyArray_S11reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4733, new_AGEMA_signal_4732, KeyArray_S11reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3105, new_AGEMA_signal_3104, KeyArray_outS11ser[5]}) ) ;
    reg_LMDPL KeyArray_S11reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4735, new_AGEMA_signal_4734, KeyArray_S11reg_gff_1_SFF_6_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3111, new_AGEMA_signal_3110, KeyArray_outS11ser[6]}) ) ;
    reg_LMDPL KeyArray_S11reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4737, new_AGEMA_signal_4736, KeyArray_S11reg_gff_1_SFF_7_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3117, new_AGEMA_signal_3116, KeyArray_outS11ser[7]}) ) ;
    reg_LMDPL KeyArray_S12reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4271, new_AGEMA_signal_4270, KeyArray_S12reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3123, new_AGEMA_signal_3122, KeyArray_outS12ser[0]}) ) ;
    reg_LMDPL KeyArray_S12reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4273, new_AGEMA_signal_4272, KeyArray_S12reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3129, new_AGEMA_signal_3128, KeyArray_outS12ser[1]}) ) ;
    reg_LMDPL KeyArray_S12reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4275, new_AGEMA_signal_4274, KeyArray_S12reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3135, new_AGEMA_signal_3134, KeyArray_outS12ser[2]}) ) ;
    reg_LMDPL KeyArray_S12reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4277, new_AGEMA_signal_4276, KeyArray_S12reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3141, new_AGEMA_signal_3140, KeyArray_outS12ser[3]}) ) ;
    reg_LMDPL KeyArray_S12reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4279, new_AGEMA_signal_4278, KeyArray_S12reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3147, new_AGEMA_signal_3146, KeyArray_outS12ser[4]}) ) ;
    reg_LMDPL KeyArray_S12reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4281, new_AGEMA_signal_4280, KeyArray_S12reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3153, new_AGEMA_signal_3152, KeyArray_outS12ser[5]}) ) ;
    reg_LMDPL KeyArray_S12reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4283, new_AGEMA_signal_4282, KeyArray_S12reg_gff_1_SFF_6_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3159, new_AGEMA_signal_3158, KeyArray_outS12ser[6]}) ) ;
    reg_LMDPL KeyArray_S12reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4285, new_AGEMA_signal_4284, KeyArray_S12reg_gff_1_SFF_7_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3165, new_AGEMA_signal_3164, KeyArray_outS12ser[7]}) ) ;
    reg_LMDPL KeyArray_S13reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4287, new_AGEMA_signal_4286, KeyArray_S13reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3173, new_AGEMA_signal_3172, keySBIn[0]}) ) ;
    reg_LMDPL KeyArray_S13reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4289, new_AGEMA_signal_4288, KeyArray_S13reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3179, new_AGEMA_signal_3178, keySBIn[1]}) ) ;
    reg_LMDPL KeyArray_S13reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4291, new_AGEMA_signal_4290, KeyArray_S13reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3185, new_AGEMA_signal_3184, keySBIn[2]}) ) ;
    reg_LMDPL KeyArray_S13reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4293, new_AGEMA_signal_4292, KeyArray_S13reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3191, new_AGEMA_signal_3190, keySBIn[3]}) ) ;
    reg_LMDPL KeyArray_S13reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4295, new_AGEMA_signal_4294, KeyArray_S13reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3197, new_AGEMA_signal_3196, keySBIn[4]}) ) ;
    reg_LMDPL KeyArray_S13reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4297, new_AGEMA_signal_4296, KeyArray_S13reg_gff_1_SFF_5_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3203, new_AGEMA_signal_3202, keySBIn[5]}) ) ;
    reg_LMDPL KeyArray_S13reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4299, new_AGEMA_signal_4298, KeyArray_S13reg_gff_1_SFF_6_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3209, new_AGEMA_signal_3208, keySBIn[6]}) ) ;
    reg_LMDPL KeyArray_S13reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4301, new_AGEMA_signal_4300, KeyArray_S13reg_gff_1_SFF_7_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3215, new_AGEMA_signal_3214, keySBIn[7]}) ) ;
    reg_LMDPL KeyArray_S20reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4741, new_AGEMA_signal_4740, KeyArray_S20reg_gff_1_SFF_0_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3221, new_AGEMA_signal_3220, KeyArray_outS20ser[0]}) ) ;
    reg_LMDPL KeyArray_S20reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4743, new_AGEMA_signal_4742, KeyArray_S20reg_gff_1_SFF_1_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3227, new_AGEMA_signal_3226, KeyArray_outS20ser[1]}) ) ;
    reg_LMDPL KeyArray_S20reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4745, new_AGEMA_signal_4744, KeyArray_S20reg_gff_1_SFF_2_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3233, new_AGEMA_signal_3232, KeyArray_outS20ser[2]}) ) ;
    reg_LMDPL KeyArray_S20reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4747, new_AGEMA_signal_4746, KeyArray_S20reg_gff_1_SFF_3_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3239, new_AGEMA_signal_3238, KeyArray_outS20ser[3]}) ) ;
    reg_LMDPL KeyArray_S20reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4749, new_AGEMA_signal_4748, KeyArray_S20reg_gff_1_SFF_4_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3245, new_AGEMA_signal_3244, KeyArray_outS20ser[4]}) ) ;
    reg_LMDPL KeyArray_S20reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4751, new_AGEMA_signal_4750, KeyArray_S20reg_gff_1_SFF_5_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3251, new_AGEMA_signal_3250, KeyArray_outS20ser[5]}) ) ;
    reg_LMDPL KeyArray_S20reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4753, new_AGEMA_signal_4752, KeyArray_S20reg_gff_1_SFF_6_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3257, new_AGEMA_signal_3256, KeyArray_outS20ser[6]}) ) ;
    reg_LMDPL KeyArray_S20reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4755, new_AGEMA_signal_4754, KeyArray_S20reg_gff_1_SFF_7_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3263, new_AGEMA_signal_3262, KeyArray_outS20ser[7]}) ) ;
    reg_LMDPL KeyArray_S21reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4757, new_AGEMA_signal_4756, KeyArray_S21reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3271, new_AGEMA_signal_3270, KeyArray_outS21ser[0]}) ) ;
    reg_LMDPL KeyArray_S21reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4759, new_AGEMA_signal_4758, KeyArray_S21reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3277, new_AGEMA_signal_3276, KeyArray_outS21ser[1]}) ) ;
    reg_LMDPL KeyArray_S21reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4761, new_AGEMA_signal_4760, KeyArray_S21reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3283, new_AGEMA_signal_3282, KeyArray_outS21ser[2]}) ) ;
    reg_LMDPL KeyArray_S21reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4763, new_AGEMA_signal_4762, KeyArray_S21reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3289, new_AGEMA_signal_3288, KeyArray_outS21ser[3]}) ) ;
    reg_LMDPL KeyArray_S21reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4765, new_AGEMA_signal_4764, KeyArray_S21reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3295, new_AGEMA_signal_3294, KeyArray_outS21ser[4]}) ) ;
    reg_LMDPL KeyArray_S21reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4767, new_AGEMA_signal_4766, KeyArray_S21reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3301, new_AGEMA_signal_3300, KeyArray_outS21ser[5]}) ) ;
    reg_LMDPL KeyArray_S21reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4769, new_AGEMA_signal_4768, KeyArray_S21reg_gff_1_SFF_6_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3307, new_AGEMA_signal_3306, KeyArray_outS21ser[6]}) ) ;
    reg_LMDPL KeyArray_S21reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4771, new_AGEMA_signal_4770, KeyArray_S21reg_gff_1_SFF_7_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3313, new_AGEMA_signal_3312, KeyArray_outS21ser[7]}) ) ;
    reg_LMDPL KeyArray_S22reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4775, new_AGEMA_signal_4774, KeyArray_S22reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3319, new_AGEMA_signal_3318, KeyArray_outS22ser[0]}) ) ;
    reg_LMDPL KeyArray_S22reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4777, new_AGEMA_signal_4776, KeyArray_S22reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3325, new_AGEMA_signal_3324, KeyArray_outS22ser[1]}) ) ;
    reg_LMDPL KeyArray_S22reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4779, new_AGEMA_signal_4778, KeyArray_S22reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3331, new_AGEMA_signal_3330, KeyArray_outS22ser[2]}) ) ;
    reg_LMDPL KeyArray_S22reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4781, new_AGEMA_signal_4780, KeyArray_S22reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3337, new_AGEMA_signal_3336, KeyArray_outS22ser[3]}) ) ;
    reg_LMDPL KeyArray_S22reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4783, new_AGEMA_signal_4782, KeyArray_S22reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3343, new_AGEMA_signal_3342, KeyArray_outS22ser[4]}) ) ;
    reg_LMDPL KeyArray_S22reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4785, new_AGEMA_signal_4784, KeyArray_S22reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3349, new_AGEMA_signal_3348, KeyArray_outS22ser[5]}) ) ;
    reg_LMDPL KeyArray_S22reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4787, new_AGEMA_signal_4786, KeyArray_S22reg_gff_1_SFF_6_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3355, new_AGEMA_signal_3354, KeyArray_outS22ser[6]}) ) ;
    reg_LMDPL KeyArray_S22reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4789, new_AGEMA_signal_4788, KeyArray_S22reg_gff_1_SFF_7_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3361, new_AGEMA_signal_3360, KeyArray_outS22ser[7]}) ) ;
    reg_LMDPL KeyArray_S23reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4791, new_AGEMA_signal_4790, KeyArray_S23reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3369, new_AGEMA_signal_3368, KeyArray_outS23ser[0]}) ) ;
    reg_LMDPL KeyArray_S23reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4793, new_AGEMA_signal_4792, KeyArray_S23reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3375, new_AGEMA_signal_3374, KeyArray_outS23ser[1]}) ) ;
    reg_LMDPL KeyArray_S23reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4795, new_AGEMA_signal_4794, KeyArray_S23reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3381, new_AGEMA_signal_3380, KeyArray_outS23ser[2]}) ) ;
    reg_LMDPL KeyArray_S23reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4797, new_AGEMA_signal_4796, KeyArray_S23reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3387, new_AGEMA_signal_3386, KeyArray_outS23ser[3]}) ) ;
    reg_LMDPL KeyArray_S23reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4799, new_AGEMA_signal_4798, KeyArray_S23reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3393, new_AGEMA_signal_3392, KeyArray_outS23ser[4]}) ) ;
    reg_LMDPL KeyArray_S23reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4801, new_AGEMA_signal_4800, KeyArray_S23reg_gff_1_SFF_5_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3399, new_AGEMA_signal_3398, KeyArray_outS23ser[5]}) ) ;
    reg_LMDPL KeyArray_S23reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4803, new_AGEMA_signal_4802, KeyArray_S23reg_gff_1_SFF_6_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3405, new_AGEMA_signal_3404, KeyArray_outS23ser[6]}) ) ;
    reg_LMDPL KeyArray_S23reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4805, new_AGEMA_signal_4804, KeyArray_S23reg_gff_1_SFF_7_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3411, new_AGEMA_signal_3410, KeyArray_outS23ser[7]}) ) ;
    reg_LMDPL KeyArray_S30reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5141, new_AGEMA_signal_5140, KeyArray_S30reg_gff_1_SFF_0_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3417, new_AGEMA_signal_3416, KeyArray_outS30ser[0]}) ) ;
    reg_LMDPL KeyArray_S30reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5171, new_AGEMA_signal_5170, KeyArray_S30reg_gff_1_SFF_1_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3423, new_AGEMA_signal_3422, KeyArray_outS30ser[1]}) ) ;
    reg_LMDPL KeyArray_S30reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5173, new_AGEMA_signal_5172, KeyArray_S30reg_gff_1_SFF_2_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3429, new_AGEMA_signal_3428, KeyArray_outS30ser[2]}) ) ;
    reg_LMDPL KeyArray_S30reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5175, new_AGEMA_signal_5174, KeyArray_S30reg_gff_1_SFF_3_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3435, new_AGEMA_signal_3434, KeyArray_outS30ser[3]}) ) ;
    reg_LMDPL KeyArray_S30reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5177, new_AGEMA_signal_5176, KeyArray_S30reg_gff_1_SFF_4_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3441, new_AGEMA_signal_3440, KeyArray_outS30ser[4]}) ) ;
    reg_LMDPL KeyArray_S30reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5179, new_AGEMA_signal_5178, KeyArray_S30reg_gff_1_SFF_5_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3447, new_AGEMA_signal_3446, KeyArray_outS30ser[5]}) ) ;
    reg_LMDPL KeyArray_S30reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5181, new_AGEMA_signal_5180, KeyArray_S30reg_gff_1_SFF_6_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3453, new_AGEMA_signal_3452, KeyArray_outS30ser[6]}) ) ;
    reg_LMDPL KeyArray_S30reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_5183, new_AGEMA_signal_5182, KeyArray_S30reg_gff_1_SFF_7_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3459, new_AGEMA_signal_3458, KeyArray_outS30ser[7]}) ) ;
    reg_LMDPL KeyArray_S31reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4809, new_AGEMA_signal_4808, KeyArray_S31reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3467, new_AGEMA_signal_3466, KeyArray_outS31ser[0]}) ) ;
    reg_LMDPL KeyArray_S31reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4811, new_AGEMA_signal_4810, KeyArray_S31reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3473, new_AGEMA_signal_3472, KeyArray_outS31ser[1]}) ) ;
    reg_LMDPL KeyArray_S31reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4813, new_AGEMA_signal_4812, KeyArray_S31reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3479, new_AGEMA_signal_3478, KeyArray_outS31ser[2]}) ) ;
    reg_LMDPL KeyArray_S31reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4815, new_AGEMA_signal_4814, KeyArray_S31reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3485, new_AGEMA_signal_3484, KeyArray_outS31ser[3]}) ) ;
    reg_LMDPL KeyArray_S31reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4817, new_AGEMA_signal_4816, KeyArray_S31reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3491, new_AGEMA_signal_3490, KeyArray_outS31ser[4]}) ) ;
    reg_LMDPL KeyArray_S31reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4819, new_AGEMA_signal_4818, KeyArray_S31reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3497, new_AGEMA_signal_3496, KeyArray_outS31ser[5]}) ) ;
    reg_LMDPL KeyArray_S31reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4821, new_AGEMA_signal_4820, KeyArray_S31reg_gff_1_SFF_6_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3503, new_AGEMA_signal_3502, KeyArray_outS31ser[6]}) ) ;
    reg_LMDPL KeyArray_S31reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4823, new_AGEMA_signal_4822, KeyArray_S31reg_gff_1_SFF_7_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3509, new_AGEMA_signal_3508, KeyArray_outS31ser[7]}) ) ;
    reg_LMDPL KeyArray_S32reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4827, new_AGEMA_signal_4826, KeyArray_S32reg_gff_1_SFF_0_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3515, new_AGEMA_signal_3514, KeyArray_outS32ser[0]}) ) ;
    reg_LMDPL KeyArray_S32reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4829, new_AGEMA_signal_4828, KeyArray_S32reg_gff_1_SFF_1_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3521, new_AGEMA_signal_3520, KeyArray_outS32ser[1]}) ) ;
    reg_LMDPL KeyArray_S32reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4831, new_AGEMA_signal_4830, KeyArray_S32reg_gff_1_SFF_2_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3527, new_AGEMA_signal_3526, KeyArray_outS32ser[2]}) ) ;
    reg_LMDPL KeyArray_S32reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4833, new_AGEMA_signal_4832, KeyArray_S32reg_gff_1_SFF_3_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3533, new_AGEMA_signal_3532, KeyArray_outS32ser[3]}) ) ;
    reg_LMDPL KeyArray_S32reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4835, new_AGEMA_signal_4834, KeyArray_S32reg_gff_1_SFF_4_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3539, new_AGEMA_signal_3538, KeyArray_outS32ser[4]}) ) ;
    reg_LMDPL KeyArray_S32reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4837, new_AGEMA_signal_4836, KeyArray_S32reg_gff_1_SFF_5_n6}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3545, new_AGEMA_signal_3544, KeyArray_outS32ser[5]}) ) ;
    reg_LMDPL KeyArray_S32reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4839, new_AGEMA_signal_4838, KeyArray_S32reg_gff_1_SFF_6_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3551, new_AGEMA_signal_3550, KeyArray_outS32ser[6]}) ) ;
    reg_LMDPL KeyArray_S32reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4841, new_AGEMA_signal_4840, KeyArray_S32reg_gff_1_SFF_7_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3557, new_AGEMA_signal_3556, KeyArray_outS32ser[7]}) ) ;
    reg_LMDPL KeyArray_S33reg_gff_1_SFF_0_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4843, new_AGEMA_signal_4842, KeyArray_S33reg_gff_1_SFF_0_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3565, new_AGEMA_signal_3564, KeyArray_outS33ser[0]}) ) ;
    reg_LMDPL KeyArray_S33reg_gff_1_SFF_1_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4845, new_AGEMA_signal_4844, KeyArray_S33reg_gff_1_SFF_1_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3571, new_AGEMA_signal_3570, KeyArray_outS33ser[1]}) ) ;
    reg_LMDPL KeyArray_S33reg_gff_1_SFF_2_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4847, new_AGEMA_signal_4846, KeyArray_S33reg_gff_1_SFF_2_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3577, new_AGEMA_signal_3576, KeyArray_outS33ser[2]}) ) ;
    reg_LMDPL KeyArray_S33reg_gff_1_SFF_3_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4849, new_AGEMA_signal_4848, KeyArray_S33reg_gff_1_SFF_3_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3583, new_AGEMA_signal_3582, KeyArray_outS33ser[3]}) ) ;
    reg_LMDPL KeyArray_S33reg_gff_1_SFF_4_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4851, new_AGEMA_signal_4850, KeyArray_S33reg_gff_1_SFF_4_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3589, new_AGEMA_signal_3588, KeyArray_outS33ser[4]}) ) ;
    reg_LMDPL KeyArray_S33reg_gff_1_SFF_5_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4853, new_AGEMA_signal_4852, KeyArray_S33reg_gff_1_SFF_5_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3595, new_AGEMA_signal_3594, KeyArray_outS33ser[5]}) ) ;
    reg_LMDPL KeyArray_S33reg_gff_1_SFF_6_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4855, new_AGEMA_signal_4854, KeyArray_S33reg_gff_1_SFF_6_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3601, new_AGEMA_signal_3600, KeyArray_outS33ser[6]}) ) ;
    reg_LMDPL KeyArray_S33reg_gff_1_SFF_7_Q_reg_FF_FF ( .D ({new_AGEMA_signal_4857, new_AGEMA_signal_4856, KeyArray_S33reg_gff_1_SFF_7_n5}), .Po_rst (Po_rst), .en (LMDPL_pre1), .clk (clk), .Q ({new_AGEMA_signal_3607, new_AGEMA_signal_3606, KeyArray_outS33ser[7]}) ) ;
    reg_sr_LMDPL calcRCon_s_current_state_reg_0__FF_FF ( .D (calcRCon_n51), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (calcRCon_s_current_state_0_), .QN () ) ;
    reg_sr_LMDPL calcRCon_s_current_state_reg_1__FF_FF ( .D (calcRCon_n50), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (calcRCon_s_current_state_1_), .QN () ) ;
    reg_sr_LMDPL calcRCon_s_current_state_reg_2__FF_FF ( .D (calcRCon_n49), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (calcRCon_s_current_state_2_), .QN () ) ;
    reg_sr_LMDPL calcRCon_s_current_state_reg_3__FF_FF ( .D (calcRCon_n48), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (calcRCon_s_current_state_3_), .QN () ) ;
    reg_sr_LMDPL calcRCon_s_current_state_reg_4__FF_FF ( .D (calcRCon_n47), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (calcRCon_s_current_state_4_), .QN () ) ;
    reg_sr_LMDPL calcRCon_s_current_state_reg_5__FF_FF ( .D (calcRCon_n46), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (calcRCon_s_current_state_5_), .QN () ) ;
    reg_sr_LMDPL calcRCon_s_current_state_reg_6__FF_FF ( .D (calcRCon_n45), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (calcRCon_s_current_state_6_), .QN () ) ;
    reg_sr_LMDPL calcRCon_s_current_state_reg_7__FF_FF ( .D (calcRCon_n44), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (calcRCon_n3), .QN () ) ;
    reg_sr_LMDPL nReset_reg_FF_FF ( .D (n9), .clk (clk), .Po_rst (Po_rst), .en (LMDPL_pre1), .Q (nReset), .QN () ) ;
endmodule
