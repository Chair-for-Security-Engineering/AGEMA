module Reg1(x, y);
 input [325:0] x;
 output [324:0] y;

  assign y[0] = x[325];
  assign y[5] = x[0];
  assign y[6] = x[11];
  assign y[7] = x[22];
  assign y[8] = x[33];
  assign y[9] = x[44];
  assign y[10] = x[55];
  assign y[11] = x[60];
  assign y[12] = x[61];
  assign y[13] = x[62];
  assign y[14] = x[63];
  assign y[15] = x[1];
  assign y[16] = x[2];
  assign y[17] = x[3];
  assign y[18] = x[4];
  assign y[19] = x[5];
  assign y[20] = x[6];
  assign y[21] = x[7];
  assign y[22] = x[8];
  assign y[23] = x[9];
  assign y[24] = x[10];
  assign y[25] = x[12];
  assign y[26] = x[13];
  assign y[27] = x[14];
  assign y[28] = x[15];
  assign y[29] = x[16];
  assign y[30] = x[17];
  assign y[31] = x[18];
  assign y[32] = x[19];
  assign y[33] = x[20];
  assign y[34] = x[21];
  assign y[35] = x[23];
  assign y[36] = x[24];
  assign y[37] = x[25];
  assign y[38] = x[26];
  assign y[39] = x[27];
  assign y[40] = x[28];
  assign y[41] = x[29];
  assign y[42] = x[30];
  assign y[43] = x[31];
  assign y[44] = x[32];
  assign y[45] = x[34];
  assign y[46] = x[35];
  assign y[47] = x[36];
  assign y[48] = x[37];
  assign y[49] = x[38];
  assign y[50] = x[39];
  assign y[51] = x[40];
  assign y[52] = x[41];
  assign y[53] = x[42];
  assign y[54] = x[43];
  assign y[55] = x[45];
  assign y[56] = x[46];
  assign y[57] = x[47];
  assign y[58] = x[48];
  assign y[59] = x[49];
  assign y[60] = x[50];
  assign y[61] = x[51];
  assign y[62] = x[52];
  assign y[63] = x[53];
  assign y[64] = x[54];
  assign y[65] = x[56];
  assign y[66] = x[57];
  assign y[67] = x[58];
  assign y[68] = x[59];
  assign y[133] = x[64];
  assign y[134] = x[75];
  assign y[135] = x[86];
  assign y[136] = x[97];
  assign y[137] = x[108];
  assign y[138] = x[119];
  assign y[139] = x[124];
  assign y[140] = x[125];
  assign y[141] = x[126];
  assign y[142] = x[127];
  assign y[143] = x[65];
  assign y[144] = x[66];
  assign y[145] = x[67];
  assign y[146] = x[68];
  assign y[147] = x[69];
  assign y[148] = x[70];
  assign y[149] = x[71];
  assign y[150] = x[72];
  assign y[151] = x[73];
  assign y[152] = x[74];
  assign y[153] = x[76];
  assign y[154] = x[77];
  assign y[155] = x[78];
  assign y[156] = x[79];
  assign y[157] = x[80];
  assign y[158] = x[81];
  assign y[159] = x[82];
  assign y[160] = x[83];
  assign y[161] = x[84];
  assign y[162] = x[85];
  assign y[163] = x[87];
  assign y[164] = x[88];
  assign y[165] = x[89];
  assign y[166] = x[90];
  assign y[167] = x[91];
  assign y[168] = x[92];
  assign y[169] = x[93];
  assign y[170] = x[94];
  assign y[171] = x[95];
  assign y[172] = x[96];
  assign y[173] = x[98];
  assign y[174] = x[99];
  assign y[175] = x[100];
  assign y[176] = x[101];
  assign y[177] = x[102];
  assign y[178] = x[103];
  assign y[179] = x[104];
  assign y[180] = x[105];
  assign y[181] = x[106];
  assign y[182] = x[107];
  assign y[183] = x[109];
  assign y[184] = x[110];
  assign y[185] = x[111];
  assign y[186] = x[112];
  assign y[187] = x[113];
  assign y[188] = x[114];
  assign y[189] = x[115];
  assign y[190] = x[116];
  assign y[191] = x[117];
  assign y[192] = x[118];
  assign y[193] = x[120];
  assign y[194] = x[121];
  assign y[195] = x[122];
  assign y[196] = x[123];
  assign y[197] = x[256];
  assign y[198] = x[267];
  assign y[199] = x[278];
  assign y[200] = x[289];
  assign y[201] = x[300];
  assign y[202] = x[311];
  assign y[203] = x[316];
  assign y[204] = x[317];
  assign y[205] = x[318];
  assign y[206] = x[319];
  assign y[207] = x[257];
  assign y[208] = x[258];
  assign y[209] = x[259];
  assign y[210] = x[260];
  assign y[211] = x[261];
  assign y[212] = x[262];
  assign y[213] = x[263];
  assign y[214] = x[264];
  assign y[215] = x[265];
  assign y[216] = x[266];
  assign y[217] = x[268];
  assign y[218] = x[269];
  assign y[219] = x[270];
  assign y[220] = x[271];
  assign y[221] = x[272];
  assign y[222] = x[273];
  assign y[223] = x[274];
  assign y[224] = x[275];
  assign y[225] = x[276];
  assign y[226] = x[277];
  assign y[227] = x[279];
  assign y[228] = x[280];
  assign y[229] = x[281];
  assign y[230] = x[282];
  assign y[231] = x[283];
  assign y[232] = x[284];
  assign y[233] = x[285];
  assign y[234] = x[286];
  assign y[235] = x[287];
  assign y[236] = x[288];
  assign y[237] = x[290];
  assign y[238] = x[291];
  assign y[239] = x[292];
  assign y[240] = x[293];
  assign y[241] = x[294];
  assign y[242] = x[295];
  assign y[243] = x[296];
  assign y[244] = x[297];
  assign y[245] = x[298];
  assign y[246] = x[299];
  assign y[247] = x[301];
  assign y[248] = x[302];
  assign y[249] = x[303];
  assign y[250] = x[304];
  assign y[251] = x[305];
  assign y[252] = x[306];
  assign y[253] = x[307];
  assign y[254] = x[308];
  assign y[255] = x[309];
  assign y[256] = x[310];
  assign y[257] = x[312];
  assign y[258] = x[313];
  assign y[259] = x[314];
  assign y[260] = x[315];
  assign y[261] = x[128];
  assign y[262] = x[139];
  assign y[263] = x[150];
  assign y[264] = x[161];
  assign y[265] = x[172];
  assign y[266] = x[183];
  assign y[267] = x[188];
  assign y[268] = x[189];
  assign y[269] = x[190];
  assign y[270] = x[191];
  assign y[271] = x[129];
  assign y[272] = x[130];
  assign y[273] = x[131];
  assign y[274] = x[132];
  assign y[275] = x[133];
  assign y[276] = x[134];
  assign y[277] = x[135];
  assign y[278] = x[136];
  assign y[279] = x[137];
  assign y[280] = x[138];
  assign y[281] = x[140];
  assign y[282] = x[141];
  assign y[283] = x[142];
  assign y[284] = x[143];
  assign y[285] = x[144];
  assign y[286] = x[145];
  assign y[287] = x[146];
  assign y[288] = x[147];
  assign y[289] = x[148];
  assign y[290] = x[149];
  assign y[291] = x[151];
  assign y[292] = x[152];
  assign y[293] = x[153];
  assign y[294] = x[154];
  assign y[295] = x[155];
  assign y[296] = x[156];
  assign y[297] = x[157];
  assign y[298] = x[158];
  assign y[299] = x[159];
  assign y[300] = x[160];
  assign y[301] = x[162];
  assign y[302] = x[163];
  assign y[303] = x[164];
  assign y[304] = x[165];
  assign y[305] = x[166];
  assign y[306] = x[167];
  assign y[307] = x[168];
  assign y[308] = x[169];
  assign y[309] = x[170];
  assign y[310] = x[171];
  assign y[311] = x[173];
  assign y[312] = x[174];
  assign y[313] = x[175];
  assign y[314] = x[176];
  assign y[315] = x[177];
  assign y[316] = x[178];
  assign y[317] = x[179];
  assign y[318] = x[180];
  assign y[319] = x[181];
  assign y[320] = x[182];
  assign y[321] = x[184];
  assign y[322] = x[185];
  assign y[323] = x[186];
  assign y[324] = x[187];
  register_stage #(.WIDTH(68)) inst_0(.clk(x[320]), .D({x[321],x[322],x[323],x[324],x[192],x[203],x[214],x[225],x[236],x[247],x[252],x[253],x[254],x[255],x[193],x[194],x[195],x[196],x[197],x[198],x[199],x[200],x[201],x[202],x[204],x[205],x[206],x[207],x[208],x[209],x[210],x[211],x[212],x[213],x[215],x[216],x[217],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[237],x[238],x[239],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[248],x[249],x[250],x[251]}), .Q({y[1],y[2],y[3],y[4],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132]}));
endmodule

module Reg2(x, y);
 input [425:0] x;
 output [424:0] y;

  assign y[0] = x[421];
  assign y[1] = x[422];
  assign y[2] = x[423];
  assign y[3] = x[424];
  assign y[4] = x[425];
  assign y[25] = x[0];
  assign y[26] = x[1];
  assign y[27] = x[2];
  assign y[28] = x[3];
  assign y[29] = x[4];
  assign y[30] = x[55];
  assign y[31] = x[56];
  assign y[32] = x[57];
  assign y[33] = x[58];
  assign y[34] = x[59];
  assign y[35] = x[75];
  assign y[36] = x[76];
  assign y[37] = x[77];
  assign y[38] = x[78];
  assign y[39] = x[79];
  assign y[40] = x[5];
  assign y[41] = x[6];
  assign y[42] = x[7];
  assign y[43] = x[8];
  assign y[44] = x[9];
  assign y[45] = x[10];
  assign y[46] = x[11];
  assign y[47] = x[12];
  assign y[48] = x[13];
  assign y[49] = x[14];
  assign y[50] = x[15];
  assign y[51] = x[16];
  assign y[52] = x[17];
  assign y[53] = x[18];
  assign y[54] = x[19];
  assign y[55] = x[20];
  assign y[56] = x[21];
  assign y[57] = x[22];
  assign y[58] = x[23];
  assign y[59] = x[24];
  assign y[60] = x[25];
  assign y[61] = x[26];
  assign y[62] = x[27];
  assign y[63] = x[28];
  assign y[64] = x[29];
  assign y[65] = x[30];
  assign y[66] = x[31];
  assign y[67] = x[32];
  assign y[68] = x[33];
  assign y[69] = x[34];
  assign y[70] = x[35];
  assign y[71] = x[36];
  assign y[72] = x[37];
  assign y[73] = x[38];
  assign y[74] = x[39];
  assign y[75] = x[40];
  assign y[76] = x[41];
  assign y[77] = x[42];
  assign y[78] = x[43];
  assign y[79] = x[44];
  assign y[80] = x[45];
  assign y[81] = x[46];
  assign y[82] = x[47];
  assign y[83] = x[48];
  assign y[84] = x[49];
  assign y[85] = x[50];
  assign y[86] = x[51];
  assign y[87] = x[52];
  assign y[88] = x[53];
  assign y[89] = x[54];
  assign y[90] = x[60];
  assign y[91] = x[61];
  assign y[92] = x[62];
  assign y[93] = x[63];
  assign y[94] = x[64];
  assign y[95] = x[65];
  assign y[96] = x[66];
  assign y[97] = x[67];
  assign y[98] = x[68];
  assign y[99] = x[69];
  assign y[100] = x[70];
  assign y[101] = x[71];
  assign y[102] = x[72];
  assign y[103] = x[73];
  assign y[104] = x[74];
  assign y[185] = x[80];
  assign y[186] = x[81];
  assign y[187] = x[82];
  assign y[188] = x[83];
  assign y[189] = x[84];
  assign y[190] = x[135];
  assign y[191] = x[136];
  assign y[192] = x[137];
  assign y[193] = x[138];
  assign y[194] = x[139];
  assign y[195] = x[155];
  assign y[196] = x[156];
  assign y[197] = x[157];
  assign y[198] = x[158];
  assign y[199] = x[159];
  assign y[200] = x[85];
  assign y[201] = x[86];
  assign y[202] = x[87];
  assign y[203] = x[88];
  assign y[204] = x[89];
  assign y[205] = x[90];
  assign y[206] = x[91];
  assign y[207] = x[92];
  assign y[208] = x[93];
  assign y[209] = x[94];
  assign y[210] = x[95];
  assign y[211] = x[96];
  assign y[212] = x[97];
  assign y[213] = x[98];
  assign y[214] = x[99];
  assign y[215] = x[100];
  assign y[216] = x[101];
  assign y[217] = x[102];
  assign y[218] = x[103];
  assign y[219] = x[104];
  assign y[220] = x[105];
  assign y[221] = x[106];
  assign y[222] = x[107];
  assign y[223] = x[108];
  assign y[224] = x[109];
  assign y[225] = x[110];
  assign y[226] = x[111];
  assign y[227] = x[112];
  assign y[228] = x[113];
  assign y[229] = x[114];
  assign y[230] = x[115];
  assign y[231] = x[116];
  assign y[232] = x[117];
  assign y[233] = x[118];
  assign y[234] = x[119];
  assign y[235] = x[120];
  assign y[236] = x[121];
  assign y[237] = x[122];
  assign y[238] = x[123];
  assign y[239] = x[124];
  assign y[240] = x[125];
  assign y[241] = x[126];
  assign y[242] = x[127];
  assign y[243] = x[128];
  assign y[244] = x[129];
  assign y[245] = x[130];
  assign y[246] = x[131];
  assign y[247] = x[132];
  assign y[248] = x[133];
  assign y[249] = x[134];
  assign y[250] = x[140];
  assign y[251] = x[141];
  assign y[252] = x[142];
  assign y[253] = x[143];
  assign y[254] = x[144];
  assign y[255] = x[145];
  assign y[256] = x[146];
  assign y[257] = x[147];
  assign y[258] = x[148];
  assign y[259] = x[149];
  assign y[260] = x[150];
  assign y[261] = x[151];
  assign y[262] = x[152];
  assign y[263] = x[153];
  assign y[264] = x[154];
  assign y[265] = x[320];
  assign y[266] = x[321];
  assign y[267] = x[322];
  assign y[268] = x[323];
  assign y[269] = x[324];
  assign y[270] = x[375];
  assign y[271] = x[376];
  assign y[272] = x[377];
  assign y[273] = x[378];
  assign y[274] = x[379];
  assign y[275] = x[395];
  assign y[276] = x[396];
  assign y[277] = x[397];
  assign y[278] = x[398];
  assign y[279] = x[399];
  assign y[280] = x[325];
  assign y[281] = x[326];
  assign y[282] = x[327];
  assign y[283] = x[328];
  assign y[284] = x[329];
  assign y[285] = x[330];
  assign y[286] = x[331];
  assign y[287] = x[332];
  assign y[288] = x[333];
  assign y[289] = x[334];
  assign y[290] = x[335];
  assign y[291] = x[336];
  assign y[292] = x[337];
  assign y[293] = x[338];
  assign y[294] = x[339];
  assign y[295] = x[340];
  assign y[296] = x[341];
  assign y[297] = x[342];
  assign y[298] = x[343];
  assign y[299] = x[344];
  assign y[300] = x[345];
  assign y[301] = x[346];
  assign y[302] = x[347];
  assign y[303] = x[348];
  assign y[304] = x[349];
  assign y[305] = x[350];
  assign y[306] = x[351];
  assign y[307] = x[352];
  assign y[308] = x[353];
  assign y[309] = x[354];
  assign y[310] = x[355];
  assign y[311] = x[356];
  assign y[312] = x[357];
  assign y[313] = x[358];
  assign y[314] = x[359];
  assign y[315] = x[360];
  assign y[316] = x[361];
  assign y[317] = x[362];
  assign y[318] = x[363];
  assign y[319] = x[364];
  assign y[320] = x[365];
  assign y[321] = x[366];
  assign y[322] = x[367];
  assign y[323] = x[368];
  assign y[324] = x[369];
  assign y[325] = x[370];
  assign y[326] = x[371];
  assign y[327] = x[372];
  assign y[328] = x[373];
  assign y[329] = x[374];
  assign y[330] = x[380];
  assign y[331] = x[381];
  assign y[332] = x[382];
  assign y[333] = x[383];
  assign y[334] = x[384];
  assign y[335] = x[385];
  assign y[336] = x[386];
  assign y[337] = x[387];
  assign y[338] = x[388];
  assign y[339] = x[389];
  assign y[340] = x[390];
  assign y[341] = x[391];
  assign y[342] = x[392];
  assign y[343] = x[393];
  assign y[344] = x[394];
  assign y[345] = x[160];
  assign y[346] = x[161];
  assign y[347] = x[162];
  assign y[348] = x[163];
  assign y[349] = x[164];
  assign y[350] = x[215];
  assign y[351] = x[216];
  assign y[352] = x[217];
  assign y[353] = x[218];
  assign y[354] = x[219];
  assign y[355] = x[235];
  assign y[356] = x[236];
  assign y[357] = x[237];
  assign y[358] = x[238];
  assign y[359] = x[239];
  assign y[360] = x[165];
  assign y[361] = x[166];
  assign y[362] = x[167];
  assign y[363] = x[168];
  assign y[364] = x[169];
  assign y[365] = x[170];
  assign y[366] = x[171];
  assign y[367] = x[172];
  assign y[368] = x[173];
  assign y[369] = x[174];
  assign y[370] = x[175];
  assign y[371] = x[176];
  assign y[372] = x[177];
  assign y[373] = x[178];
  assign y[374] = x[179];
  assign y[375] = x[180];
  assign y[376] = x[181];
  assign y[377] = x[182];
  assign y[378] = x[183];
  assign y[379] = x[184];
  assign y[380] = x[185];
  assign y[381] = x[186];
  assign y[382] = x[187];
  assign y[383] = x[188];
  assign y[384] = x[189];
  assign y[385] = x[190];
  assign y[386] = x[191];
  assign y[387] = x[192];
  assign y[388] = x[193];
  assign y[389] = x[194];
  assign y[390] = x[195];
  assign y[391] = x[196];
  assign y[392] = x[197];
  assign y[393] = x[198];
  assign y[394] = x[199];
  assign y[395] = x[200];
  assign y[396] = x[201];
  assign y[397] = x[202];
  assign y[398] = x[203];
  assign y[399] = x[204];
  assign y[400] = x[205];
  assign y[401] = x[206];
  assign y[402] = x[207];
  assign y[403] = x[208];
  assign y[404] = x[209];
  assign y[405] = x[210];
  assign y[406] = x[211];
  assign y[407] = x[212];
  assign y[408] = x[213];
  assign y[409] = x[214];
  assign y[410] = x[220];
  assign y[411] = x[221];
  assign y[412] = x[222];
  assign y[413] = x[223];
  assign y[414] = x[224];
  assign y[415] = x[225];
  assign y[416] = x[226];
  assign y[417] = x[227];
  assign y[418] = x[228];
  assign y[419] = x[229];
  assign y[420] = x[230];
  assign y[421] = x[231];
  assign y[422] = x[232];
  assign y[423] = x[233];
  assign y[424] = x[234];
  register_stage #(.WIDTH(100)) inst_0(.clk(x[400]), .D({x[401],x[402],x[403],x[404],x[405],x[406],x[407],x[408],x[409],x[410],x[411],x[412],x[413],x[414],x[415],x[416],x[417],x[418],x[419],x[420],x[240],x[241],x[242],x[243],x[244],x[295],x[296],x[297],x[298],x[299],x[315],x[316],x[317],x[318],x[319],x[245],x[246],x[247],x[248],x[249],x[250],x[251],x[252],x[253],x[254],x[255],x[256],x[257],x[258],x[259],x[260],x[261],x[262],x[263],x[264],x[265],x[266],x[267],x[268],x[269],x[270],x[271],x[272],x[273],x[274],x[275],x[276],x[277],x[278],x[279],x[280],x[281],x[282],x[283],x[284],x[285],x[286],x[287],x[288],x[289],x[290],x[291],x[292],x[293],x[294],x[300],x[301],x[302],x[303],x[304],x[305],x[306],x[307],x[308],x[309],x[310],x[311],x[312],x[313],x[314]}), .Q({y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx195(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx196(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx197(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx198(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx199(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx200(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx201(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx202(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx203(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx204(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx205(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx206(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx207(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx208(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx209(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx210(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx211(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx212(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx213(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx214(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx215(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx216(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx217(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx218(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx219(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx220(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx221(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx222(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx223(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx224(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx225(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx226(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx227(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx228(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx229(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx230(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx231(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx232(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx233(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx234(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx235(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx236(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx237(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx238(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx239(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx240(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx241(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx242(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx243(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx244(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx245(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx246(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx247(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx248(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx249(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx250(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx251(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx252(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx253(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx254(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx255(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx256(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx257(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx258(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx259(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx260(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx261(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx262(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx263(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx264(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx265(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx266(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx267(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx268(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx269(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx270(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx271(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx272(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx273(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx274(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx275(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx276(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx277(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx278(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx279(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx280(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx281(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx282(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx283(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx284(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx285(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx286(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx287(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx288(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx289(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx290(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx291(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx292(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx293(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx294(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx295(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx296(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx297(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx298(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx299(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx300(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx301(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx302(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx303(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx304(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx305(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx306(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx307(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx308(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx309(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx310(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx311(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx312(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx313(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx314(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx315(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx316(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx317(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx318(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx319(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx320(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx321(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx322(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx323(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx324(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx325(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx326(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx327(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx328(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx329(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx330(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx331(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx332(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx333(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx334(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx335(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx336(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx337(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx338(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx339(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx340(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx341(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx342(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx343(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx344(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx345(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx346(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx347(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx348(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx349(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx350(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx351(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx352(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx353(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx354(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx355(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx356(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx357(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx358(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx359(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx360(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx361(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx362(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx363(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx364(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx365(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx366(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx367(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx368(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx369(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx370(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx371(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx372(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx373(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx374(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx375(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx376(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx377(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx378(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx379(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx380(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx381(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx382(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx383(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx384(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx385(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx386(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx387(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx388(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx389(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx390(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx391(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx392(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx393(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx394(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx395(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx396(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx397(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx398(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx399(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx400(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx401(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx402(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx403(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx404(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx405(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx406(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx407(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx408(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx409(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx410(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx411(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx412(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx413(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx414(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx415(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx416(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx417(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx418(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx419(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx420(x, y);
 input [4:0] x;
 output y;

 wire t;
  assign t = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign y = t ^ x[4];
endmodule

module Fx421(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx422(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx423(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx424(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [734:0] x;
 output [409:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx4 Fx4_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx5 Fx5_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx9 Fx9_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx10 Fx10_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx14 Fx14_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx15 Fx15_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx19 Fx19_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx20 Fx20_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx24 Fx24_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx25 Fx25_inst(.x({x[19], x[18], x[17], x[16], x[15]}), .y(y[10]));
  Fx26 Fx26_inst(.x({x[20], x[18]}), .y(y[11]));
  Fx27 Fx27_inst(.x({x[21], x[17]}), .y(y[12]));
  Fx28 Fx28_inst(.x({x[22], x[16]}), .y(y[13]));
  Fx29 Fx29_inst(.x({x[23], x[15]}), .y(y[14]));
  Fx30 Fx30_inst(.x({x[28], x[27], x[26], x[25], x[24]}), .y(y[15]));
  Fx31 Fx31_inst(.x({x[29], x[27]}), .y(y[16]));
  Fx32 Fx32_inst(.x({x[30], x[26]}), .y(y[17]));
  Fx33 Fx33_inst(.x({x[31], x[25]}), .y(y[18]));
  Fx34 Fx34_inst(.x({x[32], x[24]}), .y(y[19]));
  Fx35 Fx35_inst(.x({x[37], x[36], x[35], x[34], x[33]}), .y(y[20]));
  Fx36 Fx36_inst(.x({x[38], x[36]}), .y(y[21]));
  Fx37 Fx37_inst(.x({x[39], x[35]}), .y(y[22]));
  Fx38 Fx38_inst(.x({x[40], x[34]}), .y(y[23]));
  Fx39 Fx39_inst(.x({x[41], x[33]}), .y(y[24]));
  Fx40 Fx40_inst(.x({x[46], x[45], x[44], x[43], x[42]}), .y(y[25]));
  Fx41 Fx41_inst(.x({x[47], x[45]}), .y(y[26]));
  Fx42 Fx42_inst(.x({x[48], x[44]}), .y(y[27]));
  Fx43 Fx43_inst(.x({x[49], x[43]}), .y(y[28]));
  Fx44 Fx44_inst(.x({x[50], x[42]}), .y(y[29]));
  Fx45 Fx45_inst(.x({x[55], x[54], x[53], x[52], x[51]}), .y(y[30]));
  Fx46 Fx46_inst(.x({x[56], x[54]}), .y(y[31]));
  Fx47 Fx47_inst(.x({x[57], x[53]}), .y(y[32]));
  Fx48 Fx48_inst(.x({x[58], x[52]}), .y(y[33]));
  Fx49 Fx49_inst(.x({x[59], x[51]}), .y(y[34]));
  Fx50 Fx50_inst(.x({x[64], x[63], x[62], x[61], x[60]}), .y(y[35]));
  Fx51 Fx51_inst(.x({x[65], x[63]}), .y(y[36]));
  Fx52 Fx52_inst(.x({x[66], x[62]}), .y(y[37]));
  Fx53 Fx53_inst(.x({x[67], x[61]}), .y(y[38]));
  Fx54 Fx54_inst(.x({x[68], x[60]}), .y(y[39]));
  Fx55 Fx55_inst(.x({x[73], x[72], x[71], x[70], x[69]}), .y(y[40]));
  Fx56 Fx56_inst(.x({x[74], x[72]}), .y(y[41]));
  Fx57 Fx57_inst(.x({x[75], x[71]}), .y(y[42]));
  Fx58 Fx58_inst(.x({x[76], x[70]}), .y(y[43]));
  Fx59 Fx59_inst(.x({x[77], x[69]}), .y(y[44]));
  Fx60 Fx60_inst(.x({x[82], x[81], x[80], x[79], x[78]}), .y(y[45]));
  Fx61 Fx61_inst(.x({x[83], x[81]}), .y(y[46]));
  Fx62 Fx62_inst(.x({x[84], x[80]}), .y(y[47]));
  Fx63 Fx63_inst(.x({x[85], x[79]}), .y(y[48]));
  Fx64 Fx64_inst(.x({x[86], x[78]}), .y(y[49]));
  Fx65 Fx65_inst(.x({x[91], x[90], x[89], x[88], x[87]}), .y(y[50]));
  Fx66 Fx66_inst(.x({x[92], x[90]}), .y(y[51]));
  Fx67 Fx67_inst(.x({x[93], x[89]}), .y(y[52]));
  Fx68 Fx68_inst(.x({x[94], x[88]}), .y(y[53]));
  Fx69 Fx69_inst(.x({x[95], x[87]}), .y(y[54]));
  Fx70 Fx70_inst(.x({x[100], x[99], x[98], x[97], x[96]}), .y(y[55]));
  Fx71 Fx71_inst(.x({x[101], x[99]}), .y(y[56]));
  Fx72 Fx72_inst(.x({x[102], x[98]}), .y(y[57]));
  Fx73 Fx73_inst(.x({x[103], x[97]}), .y(y[58]));
  Fx74 Fx74_inst(.x({x[104], x[96]}), .y(y[59]));
  Fx75 Fx75_inst(.x({x[109], x[108], x[107], x[106], x[105]}), .y(y[60]));
  Fx76 Fx76_inst(.x({x[110], x[108]}), .y(y[61]));
  Fx77 Fx77_inst(.x({x[111], x[107]}), .y(y[62]));
  Fx78 Fx78_inst(.x({x[112], x[106]}), .y(y[63]));
  Fx79 Fx79_inst(.x({x[113], x[105]}), .y(y[64]));
  Fx80 Fx80_inst(.x({x[118], x[117], x[116], x[115], x[114]}), .y(y[65]));
  Fx81 Fx81_inst(.x({x[119], x[117]}), .y(y[66]));
  Fx82 Fx82_inst(.x({x[120], x[116]}), .y(y[67]));
  Fx83 Fx83_inst(.x({x[121], x[115]}), .y(y[68]));
  Fx84 Fx84_inst(.x({x[122], x[114]}), .y(y[69]));
  Fx85 Fx85_inst(.x({x[127], x[126], x[125], x[124], x[123]}), .y(y[70]));
  Fx86 Fx86_inst(.x({x[128], x[126]}), .y(y[71]));
  Fx87 Fx87_inst(.x({x[129], x[125]}), .y(y[72]));
  Fx88 Fx88_inst(.x({x[130], x[124]}), .y(y[73]));
  Fx89 Fx89_inst(.x({x[131], x[123]}), .y(y[74]));
  Fx90 Fx90_inst(.x({x[136], x[135], x[134], x[133], x[132]}), .y(y[75]));
  Fx91 Fx91_inst(.x({x[137], x[135]}), .y(y[76]));
  Fx92 Fx92_inst(.x({x[138], x[134]}), .y(y[77]));
  Fx93 Fx93_inst(.x({x[139], x[133]}), .y(y[78]));
  Fx94 Fx94_inst(.x({x[140], x[132]}), .y(y[79]));
  Fx95 Fx95_inst(.x({x[145], x[144], x[143], x[142], x[141]}), .y(y[80]));
  Fx96 Fx96_inst(.x({x[146], x[144]}), .y(y[81]));
  Fx97 Fx97_inst(.x({x[147], x[143]}), .y(y[82]));
  Fx98 Fx98_inst(.x({x[148], x[142]}), .y(y[83]));
  Fx99 Fx99_inst(.x({x[149], x[141]}), .y(y[84]));
  Fx100 Fx100_inst(.x({x[154], x[153], x[152], x[151], x[150]}), .y(y[85]));
  Fx101 Fx101_inst(.x({x[155], x[153]}), .y(y[86]));
  Fx102 Fx102_inst(.x({x[156], x[152]}), .y(y[87]));
  Fx103 Fx103_inst(.x({x[157], x[151]}), .y(y[88]));
  Fx104 Fx104_inst(.x({x[158], x[150]}), .y(y[89]));
  Fx105 Fx105_inst(.x({x[163], x[162], x[161], x[160], x[159]}), .y(y[90]));
  Fx106 Fx106_inst(.x({x[164], x[162]}), .y(y[91]));
  Fx107 Fx107_inst(.x({x[165], x[161]}), .y(y[92]));
  Fx108 Fx108_inst(.x({x[166], x[160]}), .y(y[93]));
  Fx109 Fx109_inst(.x({x[167], x[159]}), .y(y[94]));
  Fx110 Fx110_inst(.x({x[172], x[171], x[170], x[169], x[168]}), .y(y[95]));
  Fx111 Fx111_inst(.x({x[173], x[171]}), .y(y[96]));
  Fx112 Fx112_inst(.x({x[174], x[170]}), .y(y[97]));
  Fx113 Fx113_inst(.x({x[175], x[169]}), .y(y[98]));
  Fx114 Fx114_inst(.x({x[176], x[168]}), .y(y[99]));
  Fx115 Fx115_inst(.x({x[181], x[180], x[179], x[178], x[177]}), .y(y[100]));
  Fx116 Fx116_inst(.x({x[182], x[180]}), .y(y[101]));
  Fx117 Fx117_inst(.x({x[183], x[179]}), .y(y[102]));
  Fx118 Fx118_inst(.x({x[184], x[178]}), .y(y[103]));
  Fx119 Fx119_inst(.x({x[185], x[177]}), .y(y[104]));
  Fx120 Fx120_inst(.x({x[190], x[189], x[188], x[187], x[186]}), .y(y[105]));
  Fx121 Fx121_inst(.x({x[191], x[189]}), .y(y[106]));
  Fx122 Fx122_inst(.x({x[192], x[188]}), .y(y[107]));
  Fx123 Fx123_inst(.x({x[193], x[187]}), .y(y[108]));
  Fx124 Fx124_inst(.x({x[194], x[186]}), .y(y[109]));
  Fx125 Fx125_inst(.x({x[199], x[198], x[197], x[196], x[195]}), .y(y[110]));
  Fx126 Fx126_inst(.x({x[200], x[198]}), .y(y[111]));
  Fx127 Fx127_inst(.x({x[201], x[197]}), .y(y[112]));
  Fx128 Fx128_inst(.x({x[202], x[196]}), .y(y[113]));
  Fx129 Fx129_inst(.x({x[203], x[195]}), .y(y[114]));
  Fx130 Fx130_inst(.x({x[208], x[207], x[206], x[205], x[204]}), .y(y[115]));
  Fx131 Fx131_inst(.x({x[209], x[207]}), .y(y[116]));
  Fx132 Fx132_inst(.x({x[210], x[206]}), .y(y[117]));
  Fx133 Fx133_inst(.x({x[211], x[205]}), .y(y[118]));
  Fx134 Fx134_inst(.x({x[212], x[204]}), .y(y[119]));
  Fx135 Fx135_inst(.x({x[217], x[216], x[215], x[214], x[213]}), .y(y[120]));
  Fx136 Fx136_inst(.x({x[218], x[216]}), .y(y[121]));
  Fx137 Fx137_inst(.x({x[219], x[215]}), .y(y[122]));
  Fx138 Fx138_inst(.x({x[220], x[214]}), .y(y[123]));
  Fx139 Fx139_inst(.x({x[221], x[213]}), .y(y[124]));
  Fx140 Fx140_inst(.x({x[226], x[225], x[224], x[223], x[222]}), .y(y[125]));
  Fx141 Fx141_inst(.x({x[227], x[225]}), .y(y[126]));
  Fx142 Fx142_inst(.x({x[228], x[224]}), .y(y[127]));
  Fx143 Fx143_inst(.x({x[229], x[223]}), .y(y[128]));
  Fx144 Fx144_inst(.x({x[230], x[222]}), .y(y[129]));
  Fx145 Fx145_inst(.x({x[235], x[234], x[233], x[232], x[231]}), .y(y[130]));
  Fx146 Fx146_inst(.x({x[236], x[234]}), .y(y[131]));
  Fx147 Fx147_inst(.x({x[237], x[233]}), .y(y[132]));
  Fx148 Fx148_inst(.x({x[238], x[232]}), .y(y[133]));
  Fx149 Fx149_inst(.x({x[239], x[231]}), .y(y[134]));
  Fx150 Fx150_inst(.x({x[244], x[243], x[242], x[241], x[240]}), .y(y[135]));
  Fx151 Fx151_inst(.x({x[245], x[243]}), .y(y[136]));
  Fx152 Fx152_inst(.x({x[246], x[242]}), .y(y[137]));
  Fx153 Fx153_inst(.x({x[247], x[241]}), .y(y[138]));
  Fx154 Fx154_inst(.x({x[248], x[240]}), .y(y[139]));
  Fx155 Fx155_inst(.x({x[253], x[252], x[251], x[250], x[249]}), .y(y[140]));
  Fx156 Fx156_inst(.x({x[254], x[252]}), .y(y[141]));
  Fx157 Fx157_inst(.x({x[255], x[251]}), .y(y[142]));
  Fx158 Fx158_inst(.x({x[256], x[250]}), .y(y[143]));
  Fx159 Fx159_inst(.x({x[257], x[249]}), .y(y[144]));
  Fx160 Fx160_inst(.x({x[262], x[261], x[260], x[259], x[258]}), .y(y[145]));
  Fx161 Fx161_inst(.x({x[263], x[261]}), .y(y[146]));
  Fx162 Fx162_inst(.x({x[264], x[260]}), .y(y[147]));
  Fx163 Fx163_inst(.x({x[265], x[259]}), .y(y[148]));
  Fx164 Fx164_inst(.x({x[266], x[258]}), .y(y[149]));
  Fx165 Fx165_inst(.x({x[271], x[270], x[269], x[268], x[267]}), .y(y[150]));
  Fx166 Fx166_inst(.x({x[272], x[270]}), .y(y[151]));
  Fx167 Fx167_inst(.x({x[273], x[269]}), .y(y[152]));
  Fx168 Fx168_inst(.x({x[274], x[268]}), .y(y[153]));
  Fx169 Fx169_inst(.x({x[275], x[267]}), .y(y[154]));
  Fx170 Fx170_inst(.x({x[280], x[279], x[278], x[277], x[276]}), .y(y[155]));
  Fx171 Fx171_inst(.x({x[281], x[279]}), .y(y[156]));
  Fx172 Fx172_inst(.x({x[282], x[278]}), .y(y[157]));
  Fx173 Fx173_inst(.x({x[283], x[277]}), .y(y[158]));
  Fx174 Fx174_inst(.x({x[284], x[276]}), .y(y[159]));
  Fx175 Fx175_inst(.x({x[289], x[288], x[287], x[286], x[285]}), .y(y[160]));
  Fx176 Fx176_inst(.x({x[290], x[288]}), .y(y[161]));
  Fx177 Fx177_inst(.x({x[291], x[287]}), .y(y[162]));
  Fx178 Fx178_inst(.x({x[292], x[286]}), .y(y[163]));
  Fx179 Fx179_inst(.x({x[293], x[285]}), .y(y[164]));
  Fx180 Fx180_inst(.x({x[298], x[297], x[296], x[295], x[294]}), .y(y[165]));
  Fx181 Fx181_inst(.x({x[299], x[297]}), .y(y[166]));
  Fx182 Fx182_inst(.x({x[300], x[296]}), .y(y[167]));
  Fx183 Fx183_inst(.x({x[301], x[295]}), .y(y[168]));
  Fx184 Fx184_inst(.x({x[302], x[294]}), .y(y[169]));
  Fx185 Fx185_inst(.x({x[307], x[306], x[305], x[304], x[303]}), .y(y[170]));
  Fx186 Fx186_inst(.x({x[308], x[306]}), .y(y[171]));
  Fx187 Fx187_inst(.x({x[309], x[305]}), .y(y[172]));
  Fx188 Fx188_inst(.x({x[310], x[304]}), .y(y[173]));
  Fx189 Fx189_inst(.x({x[311], x[303]}), .y(y[174]));
  Fx190 Fx190_inst(.x({x[316], x[315], x[314], x[313], x[312]}), .y(y[175]));
  Fx191 Fx191_inst(.x({x[317], x[315]}), .y(y[176]));
  Fx192 Fx192_inst(.x({x[318], x[314]}), .y(y[177]));
  Fx193 Fx193_inst(.x({x[319], x[313]}), .y(y[178]));
  Fx194 Fx194_inst(.x({x[320], x[312]}), .y(y[179]));
  Fx195 Fx195_inst(.x({x[325], x[324], x[323], x[322], x[321]}), .y(y[180]));
  Fx196 Fx196_inst(.x({x[326], x[324]}), .y(y[181]));
  Fx197 Fx197_inst(.x({x[327], x[323]}), .y(y[182]));
  Fx198 Fx198_inst(.x({x[328], x[322]}), .y(y[183]));
  Fx199 Fx199_inst(.x({x[329], x[321]}), .y(y[184]));
  Fx200 Fx200_inst(.x({x[334], x[333], x[332], x[331], x[330]}), .y(y[185]));
  Fx201 Fx201_inst(.x({x[335], x[333]}), .y(y[186]));
  Fx202 Fx202_inst(.x({x[336], x[332]}), .y(y[187]));
  Fx203 Fx203_inst(.x({x[337], x[331]}), .y(y[188]));
  Fx204 Fx204_inst(.x({x[338], x[330]}), .y(y[189]));
  Fx205 Fx205_inst(.x({x[343], x[342], x[341], x[340], x[339]}), .y(y[190]));
  Fx206 Fx206_inst(.x({x[344], x[342]}), .y(y[191]));
  Fx207 Fx207_inst(.x({x[345], x[341]}), .y(y[192]));
  Fx208 Fx208_inst(.x({x[346], x[340]}), .y(y[193]));
  Fx209 Fx209_inst(.x({x[347], x[339]}), .y(y[194]));
  Fx210 Fx210_inst(.x({x[352], x[351], x[350], x[349], x[348]}), .y(y[195]));
  Fx211 Fx211_inst(.x({x[353], x[351]}), .y(y[196]));
  Fx212 Fx212_inst(.x({x[354], x[350]}), .y(y[197]));
  Fx213 Fx213_inst(.x({x[355], x[349]}), .y(y[198]));
  Fx214 Fx214_inst(.x({x[356], x[348]}), .y(y[199]));
  Fx215 Fx215_inst(.x({x[361], x[360], x[359], x[358], x[357]}), .y(y[200]));
  Fx216 Fx216_inst(.x({x[362], x[360]}), .y(y[201]));
  Fx217 Fx217_inst(.x({x[363], x[359]}), .y(y[202]));
  Fx218 Fx218_inst(.x({x[364], x[358]}), .y(y[203]));
  Fx219 Fx219_inst(.x({x[365], x[357]}), .y(y[204]));
  Fx220 Fx220_inst(.x({x[370], x[369], x[368], x[367], x[366]}), .y(y[205]));
  Fx221 Fx221_inst(.x({x[371], x[369]}), .y(y[206]));
  Fx222 Fx222_inst(.x({x[372], x[368]}), .y(y[207]));
  Fx223 Fx223_inst(.x({x[373], x[367]}), .y(y[208]));
  Fx224 Fx224_inst(.x({x[374], x[366]}), .y(y[209]));
  Fx225 Fx225_inst(.x({x[379], x[378], x[377], x[376], x[375]}), .y(y[210]));
  Fx226 Fx226_inst(.x({x[380], x[378]}), .y(y[211]));
  Fx227 Fx227_inst(.x({x[381], x[377]}), .y(y[212]));
  Fx228 Fx228_inst(.x({x[382], x[376]}), .y(y[213]));
  Fx229 Fx229_inst(.x({x[383], x[375]}), .y(y[214]));
  Fx230 Fx230_inst(.x({x[388], x[387], x[386], x[385], x[384]}), .y(y[215]));
  Fx231 Fx231_inst(.x({x[389], x[387]}), .y(y[216]));
  Fx232 Fx232_inst(.x({x[390], x[386]}), .y(y[217]));
  Fx233 Fx233_inst(.x({x[391], x[385]}), .y(y[218]));
  Fx234 Fx234_inst(.x({x[392], x[384]}), .y(y[219]));
  Fx235 Fx235_inst(.x({x[397], x[396], x[395], x[394], x[393]}), .y(y[220]));
  Fx236 Fx236_inst(.x({x[398], x[396]}), .y(y[221]));
  Fx237 Fx237_inst(.x({x[399], x[395]}), .y(y[222]));
  Fx238 Fx238_inst(.x({x[400], x[394]}), .y(y[223]));
  Fx239 Fx239_inst(.x({x[401], x[393]}), .y(y[224]));
  Fx240 Fx240_inst(.x({x[406], x[405], x[404], x[403], x[402]}), .y(y[225]));
  Fx241 Fx241_inst(.x({x[407], x[405]}), .y(y[226]));
  Fx242 Fx242_inst(.x({x[408], x[404]}), .y(y[227]));
  Fx243 Fx243_inst(.x({x[409], x[403]}), .y(y[228]));
  Fx244 Fx244_inst(.x({x[410], x[402]}), .y(y[229]));
  Fx245 Fx245_inst(.x({x[415], x[414], x[413], x[412], x[411]}), .y(y[230]));
  Fx246 Fx246_inst(.x({x[416], x[414]}), .y(y[231]));
  Fx247 Fx247_inst(.x({x[417], x[413]}), .y(y[232]));
  Fx248 Fx248_inst(.x({x[418], x[412]}), .y(y[233]));
  Fx249 Fx249_inst(.x({x[419], x[411]}), .y(y[234]));
  Fx250 Fx250_inst(.x({x[424], x[423], x[422], x[421], x[420]}), .y(y[235]));
  Fx251 Fx251_inst(.x({x[425], x[423]}), .y(y[236]));
  Fx252 Fx252_inst(.x({x[426], x[422]}), .y(y[237]));
  Fx253 Fx253_inst(.x({x[427], x[421]}), .y(y[238]));
  Fx254 Fx254_inst(.x({x[428], x[420]}), .y(y[239]));
  Fx255 Fx255_inst(.x({x[433], x[432], x[431], x[430], x[429]}), .y(y[240]));
  Fx256 Fx256_inst(.x({x[434], x[432]}), .y(y[241]));
  Fx257 Fx257_inst(.x({x[435], x[431]}), .y(y[242]));
  Fx258 Fx258_inst(.x({x[436], x[430]}), .y(y[243]));
  Fx259 Fx259_inst(.x({x[437], x[429]}), .y(y[244]));
  Fx260 Fx260_inst(.x({x[442], x[441], x[440], x[439], x[438]}), .y(y[245]));
  Fx261 Fx261_inst(.x({x[443], x[441]}), .y(y[246]));
  Fx262 Fx262_inst(.x({x[444], x[440]}), .y(y[247]));
  Fx263 Fx263_inst(.x({x[445], x[439]}), .y(y[248]));
  Fx264 Fx264_inst(.x({x[446], x[438]}), .y(y[249]));
  Fx265 Fx265_inst(.x({x[451], x[450], x[449], x[448], x[447]}), .y(y[250]));
  Fx266 Fx266_inst(.x({x[452], x[450]}), .y(y[251]));
  Fx267 Fx267_inst(.x({x[453], x[449]}), .y(y[252]));
  Fx268 Fx268_inst(.x({x[454], x[448]}), .y(y[253]));
  Fx269 Fx269_inst(.x({x[455], x[447]}), .y(y[254]));
  Fx270 Fx270_inst(.x({x[460], x[459], x[458], x[457], x[456]}), .y(y[255]));
  Fx271 Fx271_inst(.x({x[461], x[459]}), .y(y[256]));
  Fx272 Fx272_inst(.x({x[462], x[458]}), .y(y[257]));
  Fx273 Fx273_inst(.x({x[463], x[457]}), .y(y[258]));
  Fx274 Fx274_inst(.x({x[464], x[456]}), .y(y[259]));
  Fx275 Fx275_inst(.x({x[469], x[468], x[467], x[466], x[465]}), .y(y[260]));
  Fx276 Fx276_inst(.x({x[470], x[468]}), .y(y[261]));
  Fx277 Fx277_inst(.x({x[471], x[467]}), .y(y[262]));
  Fx278 Fx278_inst(.x({x[472], x[466]}), .y(y[263]));
  Fx279 Fx279_inst(.x({x[473], x[465]}), .y(y[264]));
  Fx280 Fx280_inst(.x({x[478], x[477], x[476], x[475], x[474]}), .y(y[265]));
  Fx281 Fx281_inst(.x({x[479], x[477]}), .y(y[266]));
  Fx282 Fx282_inst(.x({x[480], x[476]}), .y(y[267]));
  Fx283 Fx283_inst(.x({x[481], x[475]}), .y(y[268]));
  Fx284 Fx284_inst(.x({x[482], x[474]}), .y(y[269]));
  Fx285 Fx285_inst(.x({x[487], x[486], x[485], x[484], x[483]}), .y(y[270]));
  Fx286 Fx286_inst(.x({x[488], x[486]}), .y(y[271]));
  Fx287 Fx287_inst(.x({x[489], x[485]}), .y(y[272]));
  Fx288 Fx288_inst(.x({x[490], x[484]}), .y(y[273]));
  Fx289 Fx289_inst(.x({x[491], x[483]}), .y(y[274]));
  Fx290 Fx290_inst(.x({x[496], x[495], x[494], x[493], x[492]}), .y(y[275]));
  Fx291 Fx291_inst(.x({x[497], x[495]}), .y(y[276]));
  Fx292 Fx292_inst(.x({x[498], x[494]}), .y(y[277]));
  Fx293 Fx293_inst(.x({x[499], x[493]}), .y(y[278]));
  Fx294 Fx294_inst(.x({x[500], x[492]}), .y(y[279]));
  Fx295 Fx295_inst(.x({x[505], x[504], x[503], x[502], x[501]}), .y(y[280]));
  Fx296 Fx296_inst(.x({x[506], x[504]}), .y(y[281]));
  Fx297 Fx297_inst(.x({x[507], x[503]}), .y(y[282]));
  Fx298 Fx298_inst(.x({x[508], x[502]}), .y(y[283]));
  Fx299 Fx299_inst(.x({x[509], x[501]}), .y(y[284]));
  Fx300 Fx300_inst(.x({x[514], x[513], x[512], x[511], x[510]}), .y(y[285]));
  Fx301 Fx301_inst(.x({x[515], x[513]}), .y(y[286]));
  Fx302 Fx302_inst(.x({x[516], x[512]}), .y(y[287]));
  Fx303 Fx303_inst(.x({x[517], x[511]}), .y(y[288]));
  Fx304 Fx304_inst(.x({x[518], x[510]}), .y(y[289]));
  Fx305 Fx305_inst(.x({x[523], x[522], x[521], x[520], x[519]}), .y(y[290]));
  Fx306 Fx306_inst(.x({x[524], x[522]}), .y(y[291]));
  Fx307 Fx307_inst(.x({x[525], x[521]}), .y(y[292]));
  Fx308 Fx308_inst(.x({x[526], x[520]}), .y(y[293]));
  Fx309 Fx309_inst(.x({x[527], x[519]}), .y(y[294]));
  Fx310 Fx310_inst(.x({x[532], x[531], x[530], x[529], x[528]}), .y(y[295]));
  Fx311 Fx311_inst(.x({x[533], x[531]}), .y(y[296]));
  Fx312 Fx312_inst(.x({x[534], x[530]}), .y(y[297]));
  Fx313 Fx313_inst(.x({x[535], x[529]}), .y(y[298]));
  Fx314 Fx314_inst(.x({x[536], x[528]}), .y(y[299]));
  Fx315 Fx315_inst(.x({x[541], x[540], x[539], x[538], x[537]}), .y(y[300]));
  Fx316 Fx316_inst(.x({x[542], x[540]}), .y(y[301]));
  Fx317 Fx317_inst(.x({x[543], x[539]}), .y(y[302]));
  Fx318 Fx318_inst(.x({x[544], x[538]}), .y(y[303]));
  Fx319 Fx319_inst(.x({x[545], x[537]}), .y(y[304]));
  Fx320 Fx320_inst(.x({x[550], x[549], x[548], x[547], x[546]}), .y(y[305]));
  Fx321 Fx321_inst(.x({x[551], x[549]}), .y(y[306]));
  Fx322 Fx322_inst(.x({x[552], x[548]}), .y(y[307]));
  Fx323 Fx323_inst(.x({x[553], x[547]}), .y(y[308]));
  Fx324 Fx324_inst(.x({x[554], x[546]}), .y(y[309]));
  Fx325 Fx325_inst(.x({x[559], x[558], x[557], x[556], x[555]}), .y(y[310]));
  Fx326 Fx326_inst(.x({x[560], x[558]}), .y(y[311]));
  Fx327 Fx327_inst(.x({x[561], x[557]}), .y(y[312]));
  Fx328 Fx328_inst(.x({x[562], x[556]}), .y(y[313]));
  Fx329 Fx329_inst(.x({x[563], x[555]}), .y(y[314]));
  Fx330 Fx330_inst(.x({x[568], x[567], x[566], x[565], x[564]}), .y(y[315]));
  Fx331 Fx331_inst(.x({x[569], x[567]}), .y(y[316]));
  Fx332 Fx332_inst(.x({x[570], x[566]}), .y(y[317]));
  Fx333 Fx333_inst(.x({x[571], x[565]}), .y(y[318]));
  Fx334 Fx334_inst(.x({x[572], x[564]}), .y(y[319]));
  Fx335 Fx335_inst(.x({x[577], x[576], x[575], x[574], x[573]}), .y(y[320]));
  Fx336 Fx336_inst(.x({x[578], x[576]}), .y(y[321]));
  Fx337 Fx337_inst(.x({x[579], x[575]}), .y(y[322]));
  Fx338 Fx338_inst(.x({x[580], x[574]}), .y(y[323]));
  Fx339 Fx339_inst(.x({x[581], x[573]}), .y(y[324]));
  Fx340 Fx340_inst(.x({x[586], x[585], x[584], x[583], x[582]}), .y(y[325]));
  Fx341 Fx341_inst(.x({x[587], x[585]}), .y(y[326]));
  Fx342 Fx342_inst(.x({x[588], x[584]}), .y(y[327]));
  Fx343 Fx343_inst(.x({x[589], x[583]}), .y(y[328]));
  Fx344 Fx344_inst(.x({x[590], x[582]}), .y(y[329]));
  Fx345 Fx345_inst(.x({x[595], x[594], x[593], x[592], x[591]}), .y(y[330]));
  Fx346 Fx346_inst(.x({x[596], x[594]}), .y(y[331]));
  Fx347 Fx347_inst(.x({x[597], x[593]}), .y(y[332]));
  Fx348 Fx348_inst(.x({x[598], x[592]}), .y(y[333]));
  Fx349 Fx349_inst(.x({x[599], x[591]}), .y(y[334]));
  Fx350 Fx350_inst(.x({x[604], x[603], x[602], x[601], x[600]}), .y(y[335]));
  Fx351 Fx351_inst(.x({x[605], x[603]}), .y(y[336]));
  Fx352 Fx352_inst(.x({x[606], x[602]}), .y(y[337]));
  Fx353 Fx353_inst(.x({x[607], x[601]}), .y(y[338]));
  Fx354 Fx354_inst(.x({x[608], x[600]}), .y(y[339]));
  Fx355 Fx355_inst(.x({x[613], x[612], x[611], x[610], x[609]}), .y(y[340]));
  Fx356 Fx356_inst(.x({x[614], x[612]}), .y(y[341]));
  Fx357 Fx357_inst(.x({x[615], x[611]}), .y(y[342]));
  Fx358 Fx358_inst(.x({x[616], x[610]}), .y(y[343]));
  Fx359 Fx359_inst(.x({x[617], x[609]}), .y(y[344]));
  Fx360 Fx360_inst(.x({x[622], x[621], x[620], x[619], x[618]}), .y(y[345]));
  Fx361 Fx361_inst(.x({x[623], x[621]}), .y(y[346]));
  Fx362 Fx362_inst(.x({x[624], x[620]}), .y(y[347]));
  Fx363 Fx363_inst(.x({x[625], x[619]}), .y(y[348]));
  Fx364 Fx364_inst(.x({x[626], x[618]}), .y(y[349]));
  Fx365 Fx365_inst(.x({x[631], x[630], x[629], x[628], x[627]}), .y(y[350]));
  Fx366 Fx366_inst(.x({x[632], x[630]}), .y(y[351]));
  Fx367 Fx367_inst(.x({x[633], x[629]}), .y(y[352]));
  Fx368 Fx368_inst(.x({x[634], x[628]}), .y(y[353]));
  Fx369 Fx369_inst(.x({x[635], x[627]}), .y(y[354]));
  Fx370 Fx370_inst(.x({x[640], x[639], x[638], x[637], x[636]}), .y(y[355]));
  Fx371 Fx371_inst(.x({x[641], x[639]}), .y(y[356]));
  Fx372 Fx372_inst(.x({x[642], x[638]}), .y(y[357]));
  Fx373 Fx373_inst(.x({x[643], x[637]}), .y(y[358]));
  Fx374 Fx374_inst(.x({x[644], x[636]}), .y(y[359]));
  Fx375 Fx375_inst(.x({x[649], x[648], x[647], x[646], x[645]}), .y(y[360]));
  Fx376 Fx376_inst(.x({x[650], x[648]}), .y(y[361]));
  Fx377 Fx377_inst(.x({x[651], x[647]}), .y(y[362]));
  Fx378 Fx378_inst(.x({x[652], x[646]}), .y(y[363]));
  Fx379 Fx379_inst(.x({x[653], x[645]}), .y(y[364]));
  Fx380 Fx380_inst(.x({x[658], x[657], x[656], x[655], x[654]}), .y(y[365]));
  Fx381 Fx381_inst(.x({x[659], x[657]}), .y(y[366]));
  Fx382 Fx382_inst(.x({x[660], x[656]}), .y(y[367]));
  Fx383 Fx383_inst(.x({x[661], x[655]}), .y(y[368]));
  Fx384 Fx384_inst(.x({x[662], x[654]}), .y(y[369]));
  Fx385 Fx385_inst(.x({x[667], x[666], x[665], x[664], x[663]}), .y(y[370]));
  Fx386 Fx386_inst(.x({x[668], x[666]}), .y(y[371]));
  Fx387 Fx387_inst(.x({x[669], x[665]}), .y(y[372]));
  Fx388 Fx388_inst(.x({x[670], x[664]}), .y(y[373]));
  Fx389 Fx389_inst(.x({x[671], x[663]}), .y(y[374]));
  Fx390 Fx390_inst(.x({x[676], x[675], x[674], x[673], x[672]}), .y(y[375]));
  Fx391 Fx391_inst(.x({x[677], x[675]}), .y(y[376]));
  Fx392 Fx392_inst(.x({x[678], x[674]}), .y(y[377]));
  Fx393 Fx393_inst(.x({x[679], x[673]}), .y(y[378]));
  Fx394 Fx394_inst(.x({x[680], x[672]}), .y(y[379]));
  Fx395 Fx395_inst(.x({x[685], x[684], x[683], x[682], x[681]}), .y(y[380]));
  Fx396 Fx396_inst(.x({x[686], x[684]}), .y(y[381]));
  Fx397 Fx397_inst(.x({x[687], x[683]}), .y(y[382]));
  Fx398 Fx398_inst(.x({x[688], x[682]}), .y(y[383]));
  Fx399 Fx399_inst(.x({x[689], x[681]}), .y(y[384]));
  Fx400 Fx400_inst(.x({x[694], x[693], x[692], x[691], x[690]}), .y(y[385]));
  Fx401 Fx401_inst(.x({x[695], x[693]}), .y(y[386]));
  Fx402 Fx402_inst(.x({x[696], x[692]}), .y(y[387]));
  Fx403 Fx403_inst(.x({x[697], x[691]}), .y(y[388]));
  Fx404 Fx404_inst(.x({x[698], x[690]}), .y(y[389]));
  Fx405 Fx405_inst(.x({x[703], x[702], x[701], x[700], x[699]}), .y(y[390]));
  Fx406 Fx406_inst(.x({x[704], x[702]}), .y(y[391]));
  Fx407 Fx407_inst(.x({x[705], x[701]}), .y(y[392]));
  Fx408 Fx408_inst(.x({x[706], x[700]}), .y(y[393]));
  Fx409 Fx409_inst(.x({x[707], x[699]}), .y(y[394]));
  Fx410 Fx410_inst(.x({x[712], x[711], x[710], x[709], x[708]}), .y(y[395]));
  Fx411 Fx411_inst(.x({x[713], x[711]}), .y(y[396]));
  Fx412 Fx412_inst(.x({x[714], x[710]}), .y(y[397]));
  Fx413 Fx413_inst(.x({x[715], x[709]}), .y(y[398]));
  Fx414 Fx414_inst(.x({x[716], x[708]}), .y(y[399]));
  Fx415 Fx415_inst(.x({x[721], x[720], x[719], x[718], x[717]}), .y(y[400]));
  Fx416 Fx416_inst(.x({x[722], x[720]}), .y(y[401]));
  Fx417 Fx417_inst(.x({x[723], x[719]}), .y(y[402]));
  Fx418 Fx418_inst(.x({x[724], x[718]}), .y(y[403]));
  Fx419 Fx419_inst(.x({x[725], x[717]}), .y(y[404]));
  Fx420 Fx420_inst(.x({x[730], x[729], x[728], x[727], x[726]}), .y(y[405]));
  Fx421 Fx421_inst(.x({x[731], x[729]}), .y(y[406]));
  Fx422 Fx422_inst(.x({x[732], x[728]}), .y(y[407]));
  Fx423 Fx423_inst(.x({x[733], x[727]}), .y(y[408]));
  Fx424 Fx424_inst(.x({x[734], x[726]}), .y(y[409]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind66(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind67(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind68(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind69(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind70(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind71(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind72(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind73(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind74(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind75(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind76(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind77(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind78(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind79(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind80(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind81(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind82(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind83(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind84(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind85(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind86(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind87(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind88(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind89(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind90(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind91(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind92(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind93(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind94(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind95(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind96(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind97(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind98(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind99(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind100(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind101(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind102(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind103(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind104(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind105(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind106(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind107(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind108(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind109(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind110(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind111(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind112(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind113(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind114(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind115(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind116(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind117(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind118(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind119(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind120(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind121(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind122(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind123(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind124(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind125(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind126(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind127(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind128(x, y);
 input [4:0] x;
 output y;

 wire [2:0] t;
  assign t[0] = x[3] ^ x[4];
  assign t[1] = t[2] ^ x[2];
  assign t[2] = (x[0] & x[1]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind129(x, y);
 input [11:0] x;
 output y;

 wire [9:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[2] = t[6] ^ x[2];
  assign t[3] = t[7] ^ x[5];
  assign t[4] = t[8] ^ x[8];
  assign t[5] = t[9] ^ x[11];
  assign t[6] = (x[0] & x[1]);
  assign t[7] = (x[3] & x[4]);
  assign t[8] = (x[6] & x[7]);
  assign t[9] = (x[9] & x[10]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind130(x, y);
 input [28:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[15] ? x[10] : x[9];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[16]);
  assign t[16] = ~(t[23]);
  assign t[17] = t[25] ^ x[2];
  assign t[18] = t[26] ^ x[8];
  assign t[19] = t[27] ^ x[13];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[28] ^ x[16];
  assign t[21] = t[29] ^ x[19];
  assign t[22] = t[30] ^ x[22];
  assign t[23] = t[31] ^ x[25];
  assign t[24] = t[32] ^ x[28];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[6] & x[7]);
  assign t[27] = (x[11] & x[12]);
  assign t[28] = (x[14] & x[15]);
  assign t[29] = (x[17] & x[18]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[20] & x[21]);
  assign t[31] = (x[23] & x[24]);
  assign t[32] = (x[26] & x[27]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[7];
  assign t[7] = ~(t[18] ^ t[12]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[13] | t[14]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind131(x, y);
 input [28:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[15] ? x[10] : x[9];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[16]);
  assign t[16] = ~(t[23]);
  assign t[17] = t[25] ^ x[2];
  assign t[18] = t[26] ^ x[8];
  assign t[19] = t[27] ^ x[13];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[28] ^ x[16];
  assign t[21] = t[29] ^ x[19];
  assign t[22] = t[30] ^ x[22];
  assign t[23] = t[31] ^ x[25];
  assign t[24] = t[32] ^ x[28];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[6] & x[7]);
  assign t[27] = (x[11] & x[12]);
  assign t[28] = (x[14] & x[15]);
  assign t[29] = (x[17] & x[18]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[20] & x[21]);
  assign t[31] = (x[23] & x[24]);
  assign t[32] = (x[26] & x[27]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[7];
  assign t[7] = ~(t[18] ^ t[12]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[13] | t[14]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind132(x, y);
 input [28:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[15] ? x[10] : x[9];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[16]);
  assign t[16] = ~(t[23]);
  assign t[17] = t[25] ^ x[2];
  assign t[18] = t[26] ^ x[8];
  assign t[19] = t[27] ^ x[13];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[28] ^ x[16];
  assign t[21] = t[29] ^ x[19];
  assign t[22] = t[30] ^ x[22];
  assign t[23] = t[31] ^ x[25];
  assign t[24] = t[32] ^ x[28];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[6] & x[7]);
  assign t[27] = (x[11] & x[12]);
  assign t[28] = (x[14] & x[15]);
  assign t[29] = (x[17] & x[18]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[20] & x[21]);
  assign t[31] = (x[23] & x[24]);
  assign t[32] = (x[26] & x[27]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[7];
  assign t[7] = ~(t[18] ^ t[12]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[13] | t[14]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind133(x, y);
 input [28:0] x;
 output y;

 wire [64:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[15] ^ t[16]);
  assign t[12] = ~(t[51] ^ t[52]);
  assign t[13] = ~(t[53] & t[54]);
  assign t[14] = ~(t[55] & t[56]);
  assign t[15] = t[17] ? x[10] : x[9];
  assign t[16] = ~(t[18] & t[19]);
  assign t[17] = ~(t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[55]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[25] | t[27]);
  assign t[23] = ~(t[28]);
  assign t[24] = ~(t[29] | t[30]);
  assign t[25] = ~(t[55]);
  assign t[26] = t[53] ? t[32] : t[31];
  assign t[27] = t[53] ? t[34] : t[33];
  assign t[28] = ~(t[35] | t[36]);
  assign t[29] = ~(t[25]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[53] ? t[37] : t[33];
  assign t[31] = ~(t[38] & t[39]);
  assign t[32] = ~(t[40] & t[39]);
  assign t[33] = ~(x[4] & t[41]);
  assign t[34] = ~(t[42] & t[39]);
  assign t[35] = ~(t[29] | t[43]);
  assign t[36] = ~(t[29] | t[44]);
  assign t[37] = ~(t[56] & t[42]);
  assign t[38] = x[4] & t[54];
  assign t[39] = ~(t[56]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(x[4] | t[54]);
  assign t[41] = ~(t[54] | t[56]);
  assign t[42] = ~(x[4] | t[45]);
  assign t[43] = t[53] ? t[46] : t[34];
  assign t[44] = t[53] ? t[31] : t[47];
  assign t[45] = ~(t[54]);
  assign t[46] = ~(x[4] & t[48]);
  assign t[47] = ~(t[40] & t[56]);
  assign t[48] = ~(t[54] | t[39]);
  assign t[49] = t[57] ^ x[2];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[58] ^ x[8];
  assign t[51] = t[59] ^ x[13];
  assign t[52] = t[60] ^ x[16];
  assign t[53] = t[61] ^ x[19];
  assign t[54] = t[62] ^ x[22];
  assign t[55] = t[63] ^ x[25];
  assign t[56] = t[64] ^ x[28];
  assign t[57] = (x[0] & x[1]);
  assign t[58] = (x[6] & x[7]);
  assign t[59] = (x[11] & x[12]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = (x[14] & x[15]);
  assign t[61] = (x[17] & x[18]);
  assign t[62] = (x[20] & x[21]);
  assign t[63] = (x[23] & x[24]);
  assign t[64] = (x[26] & x[27]);
  assign t[6] = ~(t[7] ^ t[11]);
  assign t[7] = ~(t[50] ^ t[12]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[13] | t[14]);
  assign y = t[0] ? t[1] : t[49];
endmodule

module R1ind134(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind135(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind136(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind137(x, y);
 input [37:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[59] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[60] ^ t[61]);
  assign t[14] = ~(t[62] & t[63]);
  assign t[15] = ~(t[64] & t[65]);
  assign t[16] = ~(t[66] ^ t[67]);
  assign t[17] = t[19] ? x[10] : x[9];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[64]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[27] | t[29]);
  assign t[25] = ~(t[30] & t[31]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[64]);
  assign t[28] = t[62] ? t[35] : t[34];
  assign t[29] = t[62] ? t[37] : t[36];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[38] | t[39]);
  assign t[31] = ~(t[27] & t[40]);
  assign t[32] = ~(t[41] & t[42]);
  assign t[33] = t[27] | t[43];
  assign t[34] = ~(t[44] & t[45]);
  assign t[35] = ~(t[46] & t[45]);
  assign t[36] = ~(x[4] & t[47]);
  assign t[37] = ~(t[48] & t[45]);
  assign t[38] = ~(t[27] | t[49]);
  assign t[39] = ~(t[50] | t[51]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[36] & t[52]);
  assign t[41] = t[65] & t[53];
  assign t[42] = t[44] | t[46];
  assign t[43] = t[62] ? t[36] : t[37];
  assign t[44] = ~(x[4] | t[63]);
  assign t[45] = ~(t[65]);
  assign t[46] = x[4] & t[63];
  assign t[47] = ~(t[63] | t[65]);
  assign t[48] = ~(x[4] | t[54]);
  assign t[49] = t[62] ? t[34] : t[35];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[27]);
  assign t[51] = t[62] ? t[37] : t[55];
  assign t[52] = ~(t[65] & t[48]);
  assign t[53] = ~(t[27] | t[62]);
  assign t[54] = ~(t[63]);
  assign t[55] = ~(x[4] & t[56]);
  assign t[56] = ~(t[63] | t[45]);
  assign t[57] = t[68] ^ x[2];
  assign t[58] = t[69] ^ x[8];
  assign t[59] = t[70] ^ x[13];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[16];
  assign t[61] = t[72] ^ x[19];
  assign t[62] = t[73] ^ x[22];
  assign t[63] = t[74] ^ x[25];
  assign t[64] = t[75] ^ x[28];
  assign t[65] = t[76] ^ x[31];
  assign t[66] = t[77] ^ x[34];
  assign t[67] = t[78] ^ x[37];
  assign t[68] = (x[0] & x[1]);
  assign t[69] = (x[6] & x[7]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[11] & x[12]);
  assign t[71] = (x[14] & x[15]);
  assign t[72] = (x[17] & x[18]);
  assign t[73] = (x[20] & x[21]);
  assign t[74] = (x[23] & x[24]);
  assign t[75] = (x[26] & x[27]);
  assign t[76] = (x[29] & x[30]);
  assign t[77] = (x[32] & x[33]);
  assign t[78] = (x[35] & x[36]);
  assign t[7] = ~(t[58] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[57];
endmodule

module R1ind138(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind139(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind140(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind141(x, y);
 input [37:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[51] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[52] ^ t[53]);
  assign t[14] = ~(t[54] & t[55]);
  assign t[15] = ~(t[56] & t[57]);
  assign t[16] = ~(t[58] ^ t[59]);
  assign t[17] = t[19] ? x[10] : x[9];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[56]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[27] | t[29]);
  assign t[25] = t[57] & t[30];
  assign t[26] = ~(t[31]);
  assign t[27] = ~(t[32]);
  assign t[28] = t[54] ? t[34] : t[33];
  assign t[29] = t[54] ? t[36] : t[35];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[32] | t[54]);
  assign t[31] = ~(t[37] | t[38]);
  assign t[32] = ~(t[56]);
  assign t[33] = ~(t[57] & t[39]);
  assign t[34] = ~(x[4] & t[40]);
  assign t[35] = ~(t[41] & t[57]);
  assign t[36] = ~(t[42] & t[43]);
  assign t[37] = ~(t[32] | t[44]);
  assign t[38] = ~(t[32] | t[45]);
  assign t[39] = ~(x[4] | t[46]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[55] | t[57]);
  assign t[41] = ~(x[4] | t[55]);
  assign t[42] = x[4] & t[55];
  assign t[43] = ~(t[57]);
  assign t[44] = t[54] ? t[36] : t[47];
  assign t[45] = t[54] ? t[48] : t[34];
  assign t[46] = ~(t[55]);
  assign t[47] = ~(t[41] & t[43]);
  assign t[48] = ~(t[39] & t[43]);
  assign t[49] = t[60] ^ x[2];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[61] ^ x[8];
  assign t[51] = t[62] ^ x[13];
  assign t[52] = t[63] ^ x[16];
  assign t[53] = t[64] ^ x[19];
  assign t[54] = t[65] ^ x[22];
  assign t[55] = t[66] ^ x[25];
  assign t[56] = t[67] ^ x[28];
  assign t[57] = t[68] ^ x[31];
  assign t[58] = t[69] ^ x[34];
  assign t[59] = t[70] ^ x[37];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = (x[0] & x[1]);
  assign t[61] = (x[6] & x[7]);
  assign t[62] = (x[11] & x[12]);
  assign t[63] = (x[14] & x[15]);
  assign t[64] = (x[17] & x[18]);
  assign t[65] = (x[20] & x[21]);
  assign t[66] = (x[23] & x[24]);
  assign t[67] = (x[26] & x[27]);
  assign t[68] = (x[29] & x[30]);
  assign t[69] = (x[32] & x[33]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[35] & x[36]);
  assign t[7] = ~(t[50] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[49];
endmodule

module R1ind142(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind143(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind144(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind145(x, y);
 input [37:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[62] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[63] ^ t[64]);
  assign t[14] = ~(t[65] & t[66]);
  assign t[15] = ~(t[67] & t[68]);
  assign t[16] = ~(t[69] ^ t[70]);
  assign t[17] = t[19] ? x[10] : x[9];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[67]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28] & t[29]);
  assign t[25] = ~(t[26] | t[30]);
  assign t[26] = ~(t[31]);
  assign t[27] = t[65] ? t[33] : t[32];
  assign t[28] = ~(t[34] | t[35]);
  assign t[29] = ~(t[36] | t[37]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[65] ? t[39] : t[38];
  assign t[31] = ~(t[67]);
  assign t[32] = ~(t[40] & t[41]);
  assign t[33] = ~(x[4] & t[42]);
  assign t[34] = ~(t[26] | t[43]);
  assign t[35] = ~(t[44] & t[45]);
  assign t[36] = ~(t[31] | t[46]);
  assign t[37] = ~(t[31] | t[47]);
  assign t[38] = ~(t[48] & t[68]);
  assign t[39] = ~(t[49] & t[41]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(x[4] | t[50]);
  assign t[41] = ~(t[68]);
  assign t[42] = ~(t[66] | t[41]);
  assign t[43] = t[65] ? t[38] : t[39];
  assign t[44] = ~(t[51] | t[52]);
  assign t[45] = ~(t[31] & t[53]);
  assign t[46] = t[65] ? t[54] : t[39];
  assign t[47] = t[65] ? t[32] : t[55];
  assign t[48] = x[4] & t[66];
  assign t[49] = ~(x[4] | t[66]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[66]);
  assign t[51] = ~(t[31] | t[56]);
  assign t[52] = ~(t[26] | t[57]);
  assign t[53] = ~(t[55] & t[58]);
  assign t[54] = ~(t[48] & t[41]);
  assign t[55] = ~(x[4] & t[59]);
  assign t[56] = t[65] ? t[39] : t[54];
  assign t[57] = t[65] ? t[32] : t[33];
  assign t[58] = ~(t[68] & t[40]);
  assign t[59] = ~(t[66] | t[68]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[2];
  assign t[61] = t[72] ^ x[8];
  assign t[62] = t[73] ^ x[13];
  assign t[63] = t[74] ^ x[16];
  assign t[64] = t[75] ^ x[19];
  assign t[65] = t[76] ^ x[22];
  assign t[66] = t[77] ^ x[25];
  assign t[67] = t[78] ^ x[28];
  assign t[68] = t[79] ^ x[31];
  assign t[69] = t[80] ^ x[34];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[81] ^ x[37];
  assign t[71] = (x[0] & x[1]);
  assign t[72] = (x[6] & x[7]);
  assign t[73] = (x[11] & x[12]);
  assign t[74] = (x[14] & x[15]);
  assign t[75] = (x[17] & x[18]);
  assign t[76] = (x[20] & x[21]);
  assign t[77] = (x[23] & x[24]);
  assign t[78] = (x[26] & x[27]);
  assign t[79] = (x[29] & x[30]);
  assign t[7] = ~(t[61] ^ t[13]);
  assign t[80] = (x[32] & x[33]);
  assign t[81] = (x[35] & x[36]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[60];
endmodule

module R1ind146(x, y);
 input [31:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[20] ^ t[13]);
  assign t[13] = ~(t[21] ^ t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[25]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[8];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[29] ^ x[13];
  assign t[21] = t[30] ^ x[16];
  assign t[22] = t[31] ^ x[19];
  assign t[23] = t[32] ^ x[22];
  assign t[24] = t[33] ^ x[25];
  assign t[25] = t[34] ^ x[28];
  assign t[26] = t[35] ^ x[31];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[6] & x[7]);
  assign t[29] = (x[11] & x[12]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[14] & x[15]);
  assign t[31] = (x[17] & x[18]);
  assign t[32] = (x[20] & x[21]);
  assign t[33] = (x[23] & x[24]);
  assign t[34] = (x[26] & x[27]);
  assign t[35] = (x[29] & x[30]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[19] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[18];
endmodule

module R1ind147(x, y);
 input [31:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[20] ^ t[13]);
  assign t[13] = ~(t[21] ^ t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[25]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[8];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[29] ^ x[13];
  assign t[21] = t[30] ^ x[16];
  assign t[22] = t[31] ^ x[19];
  assign t[23] = t[32] ^ x[22];
  assign t[24] = t[33] ^ x[25];
  assign t[25] = t[34] ^ x[28];
  assign t[26] = t[35] ^ x[31];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[6] & x[7]);
  assign t[29] = (x[11] & x[12]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[14] & x[15]);
  assign t[31] = (x[17] & x[18]);
  assign t[32] = (x[20] & x[21]);
  assign t[33] = (x[23] & x[24]);
  assign t[34] = (x[26] & x[27]);
  assign t[35] = (x[29] & x[30]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[19] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[18];
endmodule

module R1ind148(x, y);
 input [31:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[20] ^ t[13]);
  assign t[13] = ~(t[21] ^ t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[25]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[8];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[29] ^ x[13];
  assign t[21] = t[30] ^ x[16];
  assign t[22] = t[31] ^ x[19];
  assign t[23] = t[32] ^ x[22];
  assign t[24] = t[33] ^ x[25];
  assign t[25] = t[34] ^ x[28];
  assign t[26] = t[35] ^ x[31];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[6] & x[7]);
  assign t[29] = (x[11] & x[12]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[14] & x[15]);
  assign t[31] = (x[17] & x[18]);
  assign t[32] = (x[20] & x[21]);
  assign t[33] = (x[23] & x[24]);
  assign t[34] = (x[26] & x[27]);
  assign t[35] = (x[29] & x[30]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[19] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[18];
endmodule

module R1ind149(x, y);
 input [31:0] x;
 output y;

 wire [61:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[46] ^ t[13]);
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[13] = ~(t[47] ^ t[48]);
  assign t[14] = ~(t[49] & t[50]);
  assign t[15] = ~(t[51] & t[52]);
  assign t[16] = t[18] ? x[10] : x[9];
  assign t[17] = t[19] | t[20];
  assign t[18] = ~(t[21]);
  assign t[19] = ~(t[22] & t[23]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[51]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[28] & t[29]);
  assign t[24] = ~(t[30]);
  assign t[25] = t[49] ? t[32] : t[31];
  assign t[26] = ~(t[30] | t[33]);
  assign t[27] = ~(t[30] | t[34]);
  assign t[28] = ~(t[50] | t[35]);
  assign t[29] = t[24] & t[49];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[51]);
  assign t[31] = ~(x[4] & t[36]);
  assign t[32] = ~(t[52] & t[37]);
  assign t[33] = t[49] ? t[39] : t[38];
  assign t[34] = t[49] ? t[40] : t[31];
  assign t[35] = ~(t[52]);
  assign t[36] = ~(t[50] | t[52]);
  assign t[37] = ~(x[4] | t[41]);
  assign t[38] = ~(t[42] & t[35]);
  assign t[39] = ~(t[43] & t[35]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[37] & t[35]);
  assign t[41] = ~(t[50]);
  assign t[42] = ~(x[4] | t[50]);
  assign t[43] = x[4] & t[50];
  assign t[44] = t[53] ^ x[2];
  assign t[45] = t[54] ^ x[8];
  assign t[46] = t[55] ^ x[13];
  assign t[47] = t[56] ^ x[16];
  assign t[48] = t[57] ^ x[19];
  assign t[49] = t[58] ^ x[22];
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[59] ^ x[25];
  assign t[51] = t[60] ^ x[28];
  assign t[52] = t[61] ^ x[31];
  assign t[53] = (x[0] & x[1]);
  assign t[54] = (x[6] & x[7]);
  assign t[55] = (x[11] & x[12]);
  assign t[56] = (x[14] & x[15]);
  assign t[57] = (x[17] & x[18]);
  assign t[58] = (x[20] & x[21]);
  assign t[59] = (x[23] & x[24]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = (x[26] & x[27]);
  assign t[61] = (x[29] & x[30]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[7] = ~(t[45] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[44];
endmodule

module R1ind150(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind151(x, y);
 input [37:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[14] ? x[22] : x[21];
  assign t[12] = ~(t[23] ^ t[15]);
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[26] ^ t[27]);
  assign t[16] = ~(t[20]);
  assign t[17] = t[28] ^ x[2];
  assign t[18] = t[29] ^ x[8];
  assign t[19] = t[30] ^ x[11];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[14];
  assign t[21] = t[32] ^ x[17];
  assign t[22] = t[33] ^ x[20];
  assign t[23] = t[34] ^ x[25];
  assign t[24] = t[35] ^ x[28];
  assign t[25] = t[36] ^ x[31];
  assign t[26] = t[37] ^ x[34];
  assign t[27] = t[38] ^ x[37];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[23] & x[24]);
  assign t[35] = (x[26] & x[27]);
  assign t[36] = (x[29] & x[30]);
  assign t[37] = (x[32] & x[33]);
  assign t[38] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[22] ^ t[13]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind152(x, y);
 input [37:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[14] ? x[22] : x[21];
  assign t[12] = ~(t[23] ^ t[15]);
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[26] ^ t[27]);
  assign t[16] = ~(t[20]);
  assign t[17] = t[28] ^ x[2];
  assign t[18] = t[29] ^ x[8];
  assign t[19] = t[30] ^ x[11];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[14];
  assign t[21] = t[32] ^ x[17];
  assign t[22] = t[33] ^ x[20];
  assign t[23] = t[34] ^ x[25];
  assign t[24] = t[35] ^ x[28];
  assign t[25] = t[36] ^ x[31];
  assign t[26] = t[37] ^ x[34];
  assign t[27] = t[38] ^ x[37];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[23] & x[24]);
  assign t[35] = (x[26] & x[27]);
  assign t[36] = (x[29] & x[30]);
  assign t[37] = (x[32] & x[33]);
  assign t[38] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[22] ^ t[13]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind153(x, y);
 input [37:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[52] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[53] ^ t[54]);
  assign t[14] = ~(t[55] & t[56]);
  assign t[15] = ~(t[57] & t[58]);
  assign t[16] = ~(t[59] ^ t[60]);
  assign t[17] = t[19] ? x[10] : x[9];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[57]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[28]);
  assign t[25] = ~(t[26] | t[29]);
  assign t[26] = ~(t[30]);
  assign t[27] = t[55] ? t[32] : t[31];
  assign t[28] = ~(t[33] | t[34]);
  assign t[29] = t[55] ? t[36] : t[35];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[57]);
  assign t[31] = ~(t[37] & t[38]);
  assign t[32] = ~(t[39] & t[58]);
  assign t[33] = ~(t[26] | t[40]);
  assign t[34] = ~(t[26] | t[41]);
  assign t[35] = ~(x[4] & t[42]);
  assign t[36] = ~(t[58] & t[43]);
  assign t[37] = ~(x[4] | t[56]);
  assign t[38] = ~(t[58]);
  assign t[39] = x[4] & t[56];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[55] ? t[45] : t[44];
  assign t[41] = t[55] ? t[47] : t[46];
  assign t[42] = ~(t[56] | t[58]);
  assign t[43] = ~(x[4] | t[48]);
  assign t[44] = ~(t[43] & t[38]);
  assign t[45] = ~(x[4] & t[49]);
  assign t[46] = ~(t[37] & t[58]);
  assign t[47] = ~(t[39] & t[38]);
  assign t[48] = ~(t[56]);
  assign t[49] = ~(t[56] | t[38]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[61] ^ x[2];
  assign t[51] = t[62] ^ x[8];
  assign t[52] = t[63] ^ x[13];
  assign t[53] = t[64] ^ x[16];
  assign t[54] = t[65] ^ x[19];
  assign t[55] = t[66] ^ x[22];
  assign t[56] = t[67] ^ x[25];
  assign t[57] = t[68] ^ x[28];
  assign t[58] = t[69] ^ x[31];
  assign t[59] = t[70] ^ x[34];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[37];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[6] & x[7]);
  assign t[63] = (x[11] & x[12]);
  assign t[64] = (x[14] & x[15]);
  assign t[65] = (x[17] & x[18]);
  assign t[66] = (x[20] & x[21]);
  assign t[67] = (x[23] & x[24]);
  assign t[68] = (x[26] & x[27]);
  assign t[69] = (x[29] & x[30]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[32] & x[33]);
  assign t[71] = (x[35] & x[36]);
  assign t[7] = ~(t[51] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[50];
endmodule

module R1ind154(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind155(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind156(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[10] : x[9];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind157(x, y);
 input [37:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[52] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[53] ^ t[54]);
  assign t[14] = ~(t[55] & t[56]);
  assign t[15] = ~(t[57] & t[58]);
  assign t[16] = ~(t[59] ^ t[60]);
  assign t[17] = t[19] ? x[10] : x[9];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[57]);
  assign t[23] = ~(t[27] & t[28]);
  assign t[24] = t[29] | t[30];
  assign t[25] = t[58] & t[31];
  assign t[26] = t[32] | t[33];
  assign t[27] = ~(t[31] & t[34]);
  assign t[28] = ~(t[35] & t[36]);
  assign t[29] = ~(t[37] | t[38]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[37] | t[39]);
  assign t[31] = ~(t[40] | t[55]);
  assign t[32] = ~(x[4] | t[56]);
  assign t[33] = x[4] & t[56];
  assign t[34] = ~(t[41] & t[42]);
  assign t[35] = ~(t[56] | t[43]);
  assign t[36] = t[37] & t[55];
  assign t[37] = ~(t[40]);
  assign t[38] = t[55] ? t[41] : t[44];
  assign t[39] = t[55] ? t[46] : t[45];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[57]);
  assign t[41] = ~(t[58] & t[47]);
  assign t[42] = ~(x[4] & t[35]);
  assign t[43] = ~(t[58]);
  assign t[44] = ~(x[4] & t[48]);
  assign t[45] = ~(t[33] & t[43]);
  assign t[46] = ~(t[32] & t[58]);
  assign t[47] = ~(x[4] | t[49]);
  assign t[48] = ~(t[56] | t[58]);
  assign t[49] = ~(t[56]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[61] ^ x[2];
  assign t[51] = t[62] ^ x[8];
  assign t[52] = t[63] ^ x[13];
  assign t[53] = t[64] ^ x[16];
  assign t[54] = t[65] ^ x[19];
  assign t[55] = t[66] ^ x[22];
  assign t[56] = t[67] ^ x[25];
  assign t[57] = t[68] ^ x[28];
  assign t[58] = t[69] ^ x[31];
  assign t[59] = t[70] ^ x[34];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[37];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[6] & x[7]);
  assign t[63] = (x[11] & x[12]);
  assign t[64] = (x[14] & x[15]);
  assign t[65] = (x[17] & x[18]);
  assign t[66] = (x[20] & x[21]);
  assign t[67] = (x[23] & x[24]);
  assign t[68] = (x[26] & x[27]);
  assign t[69] = (x[29] & x[30]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[32] & x[33]);
  assign t[71] = (x[35] & x[36]);
  assign t[7] = ~(t[51] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[50];
endmodule

module R1ind158(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind159(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind160(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind161(x, y);
 input [37:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[52] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[53] ^ t[54]);
  assign t[14] = ~(t[55] & t[56]);
  assign t[15] = ~(t[57] & t[58]);
  assign t[16] = ~(t[59] ^ t[60]);
  assign t[17] = t[19] ? x[9] : x[10];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] & t[26]);
  assign t[22] = ~(t[57]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[29] & t[30]);
  assign t[25] = ~(t[56] | t[31]);
  assign t[26] = t[27] & t[55];
  assign t[27] = ~(t[32]);
  assign t[28] = t[55] ? t[34] : t[33];
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[32] & t[37]);
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[57]);
  assign t[33] = ~(t[38] & t[31]);
  assign t[34] = ~(t[39] & t[58]);
  assign t[35] = ~(t[32] | t[40]);
  assign t[36] = ~(t[27] | t[41]);
  assign t[37] = ~(t[42] & t[43]);
  assign t[38] = ~(x[4] | t[56]);
  assign t[39] = x[4] & t[56];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[55] ? t[33] : t[44];
  assign t[41] = t[55] ? t[46] : t[45];
  assign t[42] = ~(x[4] & t[47]);
  assign t[43] = ~(t[58] & t[48]);
  assign t[44] = ~(t[39] & t[31]);
  assign t[45] = ~(x[4] & t[25]);
  assign t[46] = ~(t[48] & t[31]);
  assign t[47] = ~(t[56] | t[58]);
  assign t[48] = ~(x[4] | t[49]);
  assign t[49] = ~(t[56]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = t[61] ^ x[2];
  assign t[51] = t[62] ^ x[8];
  assign t[52] = t[63] ^ x[13];
  assign t[53] = t[64] ^ x[16];
  assign t[54] = t[65] ^ x[19];
  assign t[55] = t[66] ^ x[22];
  assign t[56] = t[67] ^ x[25];
  assign t[57] = t[68] ^ x[28];
  assign t[58] = t[69] ^ x[31];
  assign t[59] = t[70] ^ x[34];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[37];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[6] & x[7]);
  assign t[63] = (x[11] & x[12]);
  assign t[64] = (x[14] & x[15]);
  assign t[65] = (x[17] & x[18]);
  assign t[66] = (x[20] & x[21]);
  assign t[67] = (x[23] & x[24]);
  assign t[68] = (x[26] & x[27]);
  assign t[69] = (x[29] & x[30]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[32] & x[33]);
  assign t[71] = (x[35] & x[36]);
  assign t[7] = ~(t[51] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[50];
endmodule

module R1ind162(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind163(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind164(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind165(x, y);
 input [37:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[66] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[67] ^ t[68]);
  assign t[14] = ~(t[69] & t[70]);
  assign t[15] = ~(t[71] & t[72]);
  assign t[16] = ~(t[73] ^ t[74]);
  assign t[17] = t[19] ? x[9] : x[10];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[71]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[27] | t[29]);
  assign t[25] = t[30] | t[31];
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[34]);
  assign t[28] = t[69] ? t[36] : t[35];
  assign t[29] = t[69] ? t[38] : t[37];
  assign t[2] = ~(t[5]);
  assign t[30] = ~(t[39] & t[40]);
  assign t[31] = ~(t[27] | t[41]);
  assign t[32] = ~(t[42] | t[43]);
  assign t[33] = t[34] | t[44];
  assign t[34] = ~(t[71]);
  assign t[35] = ~(t[45] & t[46]);
  assign t[36] = ~(t[47] & t[72]);
  assign t[37] = ~(t[72] & t[48]);
  assign t[38] = ~(x[4] & t[49]);
  assign t[39] = ~(t[50] | t[51]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[52] & t[53]);
  assign t[41] = t[69] ? t[37] : t[38];
  assign t[42] = ~(t[54]);
  assign t[43] = ~(t[27] | t[55]);
  assign t[44] = t[69] ? t[38] : t[56];
  assign t[45] = ~(x[4] | t[70]);
  assign t[46] = ~(t[72]);
  assign t[47] = x[4] & t[70];
  assign t[48] = ~(x[4] | t[57]);
  assign t[49] = ~(t[70] | t[72]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[34] | t[58]);
  assign t[51] = ~(t[34] | t[59]);
  assign t[52] = ~(t[70] | t[46]);
  assign t[53] = t[27] & t[69];
  assign t[54] = ~(t[60] & t[61]);
  assign t[55] = t[69] ? t[62] : t[56];
  assign t[56] = ~(t[48] & t[46]);
  assign t[57] = ~(t[70]);
  assign t[58] = t[69] ? t[63] : t[35];
  assign t[59] = t[69] ? t[56] : t[38];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = ~(t[34] | t[69]);
  assign t[61] = ~(t[37] & t[62]);
  assign t[62] = ~(x[4] & t[52]);
  assign t[63] = ~(t[47] & t[46]);
  assign t[64] = t[75] ^ x[2];
  assign t[65] = t[76] ^ x[8];
  assign t[66] = t[77] ^ x[13];
  assign t[67] = t[78] ^ x[16];
  assign t[68] = t[79] ^ x[19];
  assign t[69] = t[80] ^ x[22];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = t[81] ^ x[25];
  assign t[71] = t[82] ^ x[28];
  assign t[72] = t[83] ^ x[31];
  assign t[73] = t[84] ^ x[34];
  assign t[74] = t[85] ^ x[37];
  assign t[75] = (x[0] & x[1]);
  assign t[76] = (x[6] & x[7]);
  assign t[77] = (x[11] & x[12]);
  assign t[78] = (x[14] & x[15]);
  assign t[79] = (x[17] & x[18]);
  assign t[7] = ~(t[65] ^ t[13]);
  assign t[80] = (x[20] & x[21]);
  assign t[81] = (x[23] & x[24]);
  assign t[82] = (x[26] & x[27]);
  assign t[83] = (x[29] & x[30]);
  assign t[84] = (x[32] & x[33]);
  assign t[85] = (x[35] & x[36]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[64];
endmodule

module R1ind166(x, y);
 input [31:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[20] ^ t[13]);
  assign t[13] = ~(t[21] ^ t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[25]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[8];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[29] ^ x[13];
  assign t[21] = t[30] ^ x[16];
  assign t[22] = t[31] ^ x[19];
  assign t[23] = t[32] ^ x[22];
  assign t[24] = t[33] ^ x[25];
  assign t[25] = t[34] ^ x[28];
  assign t[26] = t[35] ^ x[31];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[6] & x[7]);
  assign t[29] = (x[11] & x[12]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[14] & x[15]);
  assign t[31] = (x[17] & x[18]);
  assign t[32] = (x[20] & x[21]);
  assign t[33] = (x[23] & x[24]);
  assign t[34] = (x[26] & x[27]);
  assign t[35] = (x[29] & x[30]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[19] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[18];
endmodule

module R1ind167(x, y);
 input [31:0] x;
 output y;

 wire [33:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[18] ? x[9] : x[10];
  assign t[12] = ~(t[19] ^ t[13]);
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[14] = ~(t[22] & t[23]);
  assign t[15] = ~(t[18] & t[24]);
  assign t[16] = t[25] ^ x[2];
  assign t[17] = t[26] ^ x[8];
  assign t[18] = t[27] ^ x[13];
  assign t[19] = t[28] ^ x[16];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[29] ^ x[19];
  assign t[21] = t[30] ^ x[22];
  assign t[22] = t[31] ^ x[25];
  assign t[23] = t[32] ^ x[28];
  assign t[24] = t[33] ^ x[31];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[6] & x[7]);
  assign t[27] = (x[11] & x[12]);
  assign t[28] = (x[14] & x[15]);
  assign t[29] = (x[17] & x[18]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[20] & x[21]);
  assign t[31] = (x[23] & x[24]);
  assign t[32] = (x[26] & x[27]);
  assign t[33] = (x[29] & x[30]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[17] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[16];
endmodule

module R1ind168(x, y);
 input [31:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[20] ^ t[13]);
  assign t[13] = ~(t[21] ^ t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[25]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[8];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[29] ^ x[13];
  assign t[21] = t[30] ^ x[16];
  assign t[22] = t[31] ^ x[19];
  assign t[23] = t[32] ^ x[22];
  assign t[24] = t[33] ^ x[25];
  assign t[25] = t[34] ^ x[28];
  assign t[26] = t[35] ^ x[31];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[6] & x[7]);
  assign t[29] = (x[11] & x[12]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[14] & x[15]);
  assign t[31] = (x[17] & x[18]);
  assign t[32] = (x[20] & x[21]);
  assign t[33] = (x[23] & x[24]);
  assign t[34] = (x[26] & x[27]);
  assign t[35] = (x[29] & x[30]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[19] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[18];
endmodule

module R1ind169(x, y);
 input [31:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[53] ^ t[13]);
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[13] = ~(t[54] ^ t[55]);
  assign t[14] = ~(t[56] & t[57]);
  assign t[15] = ~(t[58] & t[59]);
  assign t[16] = t[18] ? x[9] : x[10];
  assign t[17] = ~(t[19] & t[20]);
  assign t[18] = ~(t[21]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[58]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[26] | t[28]);
  assign t[24] = ~(t[29] | t[30]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[26] = ~(t[29]);
  assign t[27] = t[56] ? t[34] : t[33];
  assign t[28] = t[56] ? t[36] : t[35];
  assign t[29] = ~(t[58]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[56] ? t[34] : t[35];
  assign t[31] = ~(t[37] | t[38]);
  assign t[32] = ~(t[39] & t[40]);
  assign t[33] = ~(t[41] & t[59]);
  assign t[34] = ~(t[42] & t[43]);
  assign t[35] = ~(t[41] & t[43]);
  assign t[36] = ~(t[42] & t[59]);
  assign t[37] = ~(t[29] | t[44]);
  assign t[38] = ~(t[29] | t[45]);
  assign t[39] = ~(t[57] | t[43]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[26] & t[56];
  assign t[41] = x[4] & t[57];
  assign t[42] = ~(x[4] | t[57]);
  assign t[43] = ~(t[59]);
  assign t[44] = t[56] ? t[35] : t[34];
  assign t[45] = t[56] ? t[47] : t[46];
  assign t[46] = ~(x[4] & t[48]);
  assign t[47] = ~(t[49] & t[43]);
  assign t[48] = ~(t[57] | t[59]);
  assign t[49] = ~(x[4] | t[50]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[57]);
  assign t[51] = t[60] ^ x[2];
  assign t[52] = t[61] ^ x[8];
  assign t[53] = t[62] ^ x[13];
  assign t[54] = t[63] ^ x[16];
  assign t[55] = t[64] ^ x[19];
  assign t[56] = t[65] ^ x[22];
  assign t[57] = t[66] ^ x[25];
  assign t[58] = t[67] ^ x[28];
  assign t[59] = t[68] ^ x[31];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = (x[0] & x[1]);
  assign t[61] = (x[6] & x[7]);
  assign t[62] = (x[11] & x[12]);
  assign t[63] = (x[14] & x[15]);
  assign t[64] = (x[17] & x[18]);
  assign t[65] = (x[20] & x[21]);
  assign t[66] = (x[23] & x[24]);
  assign t[67] = (x[26] & x[27]);
  assign t[68] = (x[29] & x[30]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[7] = ~(t[52] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[51];
endmodule

module R1ind170(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind171(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind172(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind173(x, y);
 input [37:0] x;
 output y;

 wire [74:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[55] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[56] ^ t[57]);
  assign t[14] = ~(t[58] & t[59]);
  assign t[15] = ~(t[60] & t[61]);
  assign t[16] = ~(t[62] ^ t[63]);
  assign t[17] = t[19] ? x[9] : x[10];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[60]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[29] | t[30]);
  assign t[25] = ~(t[29] | t[31]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[60]);
  assign t[28] = t[58] ? t[35] : t[34];
  assign t[29] = ~(t[27]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[58] ? t[37] : t[36];
  assign t[31] = t[58] ? t[38] : t[34];
  assign t[32] = ~(t[39] | t[40]);
  assign t[33] = t[27] | t[41];
  assign t[34] = ~(t[42] & t[43]);
  assign t[35] = ~(t[44] & t[43]);
  assign t[36] = ~(x[4] & t[45]);
  assign t[37] = ~(t[46] & t[43]);
  assign t[38] = ~(t[44] & t[61]);
  assign t[39] = ~(t[29] | t[47]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[29] | t[48]);
  assign t[41] = t[58] ? t[49] : t[37];
  assign t[42] = x[4] & t[59];
  assign t[43] = ~(t[61]);
  assign t[44] = ~(x[4] | t[59]);
  assign t[45] = ~(t[59] | t[43]);
  assign t[46] = ~(x[4] | t[50]);
  assign t[47] = t[58] ? t[51] : t[35];
  assign t[48] = t[58] ? t[34] : t[38];
  assign t[49] = ~(x[4] & t[52]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[59]);
  assign t[51] = ~(t[42] & t[61]);
  assign t[52] = ~(t[59] | t[61]);
  assign t[53] = t[64] ^ x[2];
  assign t[54] = t[65] ^ x[8];
  assign t[55] = t[66] ^ x[13];
  assign t[56] = t[67] ^ x[16];
  assign t[57] = t[68] ^ x[19];
  assign t[58] = t[69] ^ x[22];
  assign t[59] = t[70] ^ x[25];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[28];
  assign t[61] = t[72] ^ x[31];
  assign t[62] = t[73] ^ x[34];
  assign t[63] = t[74] ^ x[37];
  assign t[64] = (x[0] & x[1]);
  assign t[65] = (x[6] & x[7]);
  assign t[66] = (x[11] & x[12]);
  assign t[67] = (x[14] & x[15]);
  assign t[68] = (x[17] & x[18]);
  assign t[69] = (x[20] & x[21]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[23] & x[24]);
  assign t[71] = (x[26] & x[27]);
  assign t[72] = (x[29] & x[30]);
  assign t[73] = (x[32] & x[33]);
  assign t[74] = (x[35] & x[36]);
  assign t[7] = ~(t[54] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[53];
endmodule

module R1ind174(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind175(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind176(x, y);
 input [37:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[16] ? x[9] : x[10];
  assign t[12] = ~(t[21] ^ t[17]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = ~(t[18]);
  assign t[17] = ~(t[28] ^ t[29]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[30] ^ x[2];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[8];
  assign t[21] = t[32] ^ x[13];
  assign t[22] = t[33] ^ x[16];
  assign t[23] = t[34] ^ x[19];
  assign t[24] = t[35] ^ x[22];
  assign t[25] = t[36] ^ x[25];
  assign t[26] = t[37] ^ x[28];
  assign t[27] = t[38] ^ x[31];
  assign t[28] = t[39] ^ x[34];
  assign t[29] = t[40] ^ x[37];
  assign t[2] = ~(t[5]);
  assign t[30] = (x[0] & x[1]);
  assign t[31] = (x[6] & x[7]);
  assign t[32] = (x[11] & x[12]);
  assign t[33] = (x[14] & x[15]);
  assign t[34] = (x[17] & x[18]);
  assign t[35] = (x[20] & x[21]);
  assign t[36] = (x[23] & x[24]);
  assign t[37] = (x[26] & x[27]);
  assign t[38] = (x[29] & x[30]);
  assign t[39] = (x[32] & x[33]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = (x[35] & x[36]);
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[20] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[19];
endmodule

module R1ind177(x, y);
 input [37:0] x;
 output y;

 wire [80:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[61] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[62] ^ t[63]);
  assign t[14] = ~(t[64] & t[65]);
  assign t[15] = ~(t[66] & t[67]);
  assign t[16] = ~(t[68] ^ t[69]);
  assign t[17] = t[19] ? x[9] : x[10];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[66]);
  assign t[23] = ~(t[27] & t[28]);
  assign t[24] = ~(t[29] & t[30]);
  assign t[25] = ~(t[31] | t[32]);
  assign t[26] = ~(t[31] | t[33]);
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = ~(t[36] & t[37]);
  assign t[29] = ~(t[38] & t[39]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[36] | t[40];
  assign t[31] = ~(t[36]);
  assign t[32] = t[64] ? t[42] : t[41];
  assign t[33] = t[64] ? t[44] : t[43];
  assign t[34] = ~(t[36] | t[45]);
  assign t[35] = ~(t[31] | t[46]);
  assign t[36] = ~(t[66]);
  assign t[37] = ~(t[47] & t[48]);
  assign t[38] = t[67] & t[49];
  assign t[39] = t[50] | t[51];
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = t[64] ? t[47] : t[52];
  assign t[41] = ~(t[50] & t[53]);
  assign t[42] = ~(t[51] & t[67]);
  assign t[43] = ~(t[50] & t[67]);
  assign t[44] = ~(t[51] & t[53]);
  assign t[45] = t[64] ? t[41] : t[44];
  assign t[46] = t[64] ? t[52] : t[54];
  assign t[47] = ~(x[4] & t[55]);
  assign t[48] = ~(t[67] & t[56]);
  assign t[49] = ~(t[36] | t[64]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(x[4] | t[65]);
  assign t[51] = x[4] & t[65];
  assign t[52] = ~(t[56] & t[53]);
  assign t[53] = ~(t[67]);
  assign t[54] = ~(x[4] & t[57]);
  assign t[55] = ~(t[65] | t[67]);
  assign t[56] = ~(x[4] | t[58]);
  assign t[57] = ~(t[65] | t[53]);
  assign t[58] = ~(t[65]);
  assign t[59] = t[70] ^ x[2];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[8];
  assign t[61] = t[72] ^ x[13];
  assign t[62] = t[73] ^ x[16];
  assign t[63] = t[74] ^ x[19];
  assign t[64] = t[75] ^ x[22];
  assign t[65] = t[76] ^ x[25];
  assign t[66] = t[77] ^ x[28];
  assign t[67] = t[78] ^ x[31];
  assign t[68] = t[79] ^ x[34];
  assign t[69] = t[80] ^ x[37];
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[0] & x[1]);
  assign t[71] = (x[6] & x[7]);
  assign t[72] = (x[11] & x[12]);
  assign t[73] = (x[14] & x[15]);
  assign t[74] = (x[17] & x[18]);
  assign t[75] = (x[20] & x[21]);
  assign t[76] = (x[23] & x[24]);
  assign t[77] = (x[26] & x[27]);
  assign t[78] = (x[29] & x[30]);
  assign t[79] = (x[32] & x[33]);
  assign t[7] = ~(t[60] ^ t[13]);
  assign t[80] = (x[35] & x[36]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[59];
endmodule

module R1ind178(x, y);
 input [37:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[18] ? x[21] : x[22];
  assign t[12] = ~(t[21] ^ t[14]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] ^ t[25]);
  assign t[15] = t[26] ^ x[2];
  assign t[16] = t[27] ^ x[8];
  assign t[17] = t[28] ^ x[11];
  assign t[18] = t[29] ^ x[14];
  assign t[19] = t[30] ^ x[17];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[20];
  assign t[21] = t[32] ^ x[25];
  assign t[22] = t[33] ^ x[28];
  assign t[23] = t[34] ^ x[31];
  assign t[24] = t[35] ^ x[34];
  assign t[25] = t[36] ^ x[37];
  assign t[26] = (x[0] & x[1]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[29] = (x[12] & x[13]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[15] & x[16]);
  assign t[31] = (x[18] & x[19]);
  assign t[32] = (x[23] & x[24]);
  assign t[33] = (x[26] & x[27]);
  assign t[34] = (x[29] & x[30]);
  assign t[35] = (x[32] & x[33]);
  assign t[36] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[16] & t[17]);
  assign t[7] = ~(t[18] & t[19]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[20] ^ t[13]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind179(x, y);
 input [37:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[18] ? x[21] : x[22];
  assign t[12] = ~(t[21] ^ t[14]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] ^ t[25]);
  assign t[15] = t[26] ^ x[2];
  assign t[16] = t[27] ^ x[8];
  assign t[17] = t[28] ^ x[11];
  assign t[18] = t[29] ^ x[14];
  assign t[19] = t[30] ^ x[17];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[20];
  assign t[21] = t[32] ^ x[25];
  assign t[22] = t[33] ^ x[28];
  assign t[23] = t[34] ^ x[31];
  assign t[24] = t[35] ^ x[34];
  assign t[25] = t[36] ^ x[37];
  assign t[26] = (x[0] & x[1]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[29] = (x[12] & x[13]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[15] & x[16]);
  assign t[31] = (x[18] & x[19]);
  assign t[32] = (x[23] & x[24]);
  assign t[33] = (x[26] & x[27]);
  assign t[34] = (x[29] & x[30]);
  assign t[35] = (x[32] & x[33]);
  assign t[36] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[16] & t[17]);
  assign t[7] = ~(t[18] & t[19]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[20] ^ t[13]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind180(x, y);
 input [37:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[18] ? x[21] : x[22];
  assign t[12] = ~(t[21] ^ t[14]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] ^ t[25]);
  assign t[15] = t[26] ^ x[2];
  assign t[16] = t[27] ^ x[8];
  assign t[17] = t[28] ^ x[11];
  assign t[18] = t[29] ^ x[14];
  assign t[19] = t[30] ^ x[17];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[20];
  assign t[21] = t[32] ^ x[25];
  assign t[22] = t[33] ^ x[28];
  assign t[23] = t[34] ^ x[31];
  assign t[24] = t[35] ^ x[34];
  assign t[25] = t[36] ^ x[37];
  assign t[26] = (x[0] & x[1]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[29] = (x[12] & x[13]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[15] & x[16]);
  assign t[31] = (x[18] & x[19]);
  assign t[32] = (x[23] & x[24]);
  assign t[33] = (x[26] & x[27]);
  assign t[34] = (x[29] & x[30]);
  assign t[35] = (x[32] & x[33]);
  assign t[36] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[16] & t[17]);
  assign t[7] = ~(t[18] & t[19]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[20] ^ t[13]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind181(x, y);
 input [37:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = ~(t[56] ^ t[14]);
  assign t[12] = ~(t[15] ^ t[16]);
  assign t[13] = ~(t[57] ^ t[58]);
  assign t[14] = ~(t[59] ^ t[60]);
  assign t[15] = t[17] ? x[21] : x[22];
  assign t[16] = ~(t[18] & t[19]);
  assign t[17] = ~(t[20]);
  assign t[18] = ~(t[21] | t[22]);
  assign t[19] = ~(t[23]);
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = ~(t[53]);
  assign t[21] = ~(t[24] & t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[28] | t[29]);
  assign t[24] = ~(t[30] & t[31]);
  assign t[25] = ~(t[32] & t[33]);
  assign t[26] = ~(t[34]);
  assign t[27] = t[35] | t[36];
  assign t[28] = ~(t[35]);
  assign t[29] = t[51] ? t[38] : t[37];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[35] | t[51]);
  assign t[31] = ~(t[39] & t[40]);
  assign t[32] = ~(t[52] | t[41]);
  assign t[33] = t[28] & t[51];
  assign t[34] = ~(t[35] | t[42]);
  assign t[35] = ~(t[53]);
  assign t[36] = t[51] ? t[44] : t[43];
  assign t[37] = ~(t[45] & t[54]);
  assign t[38] = ~(t[46] & t[41]);
  assign t[39] = ~(t[54] & t[47]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(x[4] & t[32]);
  assign t[41] = ~(t[54]);
  assign t[42] = t[51] ? t[43] : t[44];
  assign t[43] = ~(t[47] & t[41]);
  assign t[44] = ~(x[4] & t[48]);
  assign t[45] = x[4] & t[52];
  assign t[46] = ~(x[4] | t[52]);
  assign t[47] = ~(x[4] | t[49]);
  assign t[48] = ~(t[52] | t[54]);
  assign t[49] = ~(t[52]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[61] ^ x[2];
  assign t[51] = t[62] ^ x[8];
  assign t[52] = t[63] ^ x[11];
  assign t[53] = t[64] ^ x[14];
  assign t[54] = t[65] ^ x[17];
  assign t[55] = t[66] ^ x[20];
  assign t[56] = t[67] ^ x[25];
  assign t[57] = t[68] ^ x[28];
  assign t[58] = t[69] ^ x[31];
  assign t[59] = t[70] ^ x[34];
  assign t[5] = t[10] ^ x[5];
  assign t[60] = t[71] ^ x[37];
  assign t[61] = (x[0] & x[1]);
  assign t[62] = (x[6] & x[7]);
  assign t[63] = (x[9] & x[10]);
  assign t[64] = (x[12] & x[13]);
  assign t[65] = (x[15] & x[16]);
  assign t[66] = (x[18] & x[19]);
  assign t[67] = (x[23] & x[24]);
  assign t[68] = (x[26] & x[27]);
  assign t[69] = (x[29] & x[30]);
  assign t[6] = ~(t[51] & t[52]);
  assign t[70] = (x[32] & x[33]);
  assign t[71] = (x[35] & x[36]);
  assign t[7] = ~(t[53] & t[54]);
  assign t[8] = ~(t[11] ^ t[12]);
  assign t[9] = ~(t[55] ^ t[13]);
  assign y = t[0] ? t[1] : t[50];
endmodule

module R1ind182(x, y);
 input [28:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[16] ? x[21] : x[22];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[13] = t[21] ^ x[2];
  assign t[14] = t[22] ^ x[8];
  assign t[15] = t[23] ^ x[11];
  assign t[16] = t[24] ^ x[14];
  assign t[17] = t[25] ^ x[17];
  assign t[18] = t[26] ^ x[20];
  assign t[19] = t[27] ^ x[25];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[28] ^ x[28];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[6] & x[7]);
  assign t[23] = (x[9] & x[10]);
  assign t[24] = (x[12] & x[13]);
  assign t[25] = (x[15] & x[16]);
  assign t[26] = (x[18] & x[19]);
  assign t[27] = (x[23] & x[24]);
  assign t[28] = (x[26] & x[27]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[14] & t[15]);
  assign t[7] = ~(t[16] & t[17]);
  assign t[8] = t[11] ^ t[9];
  assign t[9] = ~(t[18] ^ t[12]);
  assign y = t[0] ? t[1] : t[13];
endmodule

module R1ind183(x, y);
 input [28:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[16] ? x[21] : x[22];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[13] = t[21] ^ x[2];
  assign t[14] = t[22] ^ x[8];
  assign t[15] = t[23] ^ x[11];
  assign t[16] = t[24] ^ x[14];
  assign t[17] = t[25] ^ x[17];
  assign t[18] = t[26] ^ x[20];
  assign t[19] = t[27] ^ x[25];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[28] ^ x[28];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[6] & x[7]);
  assign t[23] = (x[9] & x[10]);
  assign t[24] = (x[12] & x[13]);
  assign t[25] = (x[15] & x[16]);
  assign t[26] = (x[18] & x[19]);
  assign t[27] = (x[23] & x[24]);
  assign t[28] = (x[26] & x[27]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[14] & t[15]);
  assign t[7] = ~(t[16] & t[17]);
  assign t[8] = t[11] ^ t[9];
  assign t[9] = ~(t[18] ^ t[12]);
  assign y = t[0] ? t[1] : t[13];
endmodule

module R1ind184(x, y);
 input [28:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[16] ? x[22] : x[21];
  assign t[12] = ~(t[19] ^ t[20]);
  assign t[13] = t[21] ^ x[2];
  assign t[14] = t[22] ^ x[8];
  assign t[15] = t[23] ^ x[11];
  assign t[16] = t[24] ^ x[14];
  assign t[17] = t[25] ^ x[17];
  assign t[18] = t[26] ^ x[20];
  assign t[19] = t[27] ^ x[25];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[28] ^ x[28];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[6] & x[7]);
  assign t[23] = (x[9] & x[10]);
  assign t[24] = (x[12] & x[13]);
  assign t[25] = (x[15] & x[16]);
  assign t[26] = (x[18] & x[19]);
  assign t[27] = (x[23] & x[24]);
  assign t[28] = (x[26] & x[27]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[14] & t[15]);
  assign t[7] = ~(t[16] & t[17]);
  assign t[8] = t[11] ^ t[9];
  assign t[9] = ~(t[18] ^ t[12]);
  assign y = t[0] ? t[1] : t[13];
endmodule

module R1ind185(x, y);
 input [28:0] x;
 output y;

 wire [63:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = ~(t[13] ^ t[14]);
  assign t[12] = ~(t[54] ^ t[55]);
  assign t[13] = t[51] ? x[22] : x[21];
  assign t[14] = t[15] | t[16];
  assign t[15] = ~(t[17] & t[18]);
  assign t[16] = ~(t[19] & t[20]);
  assign t[17] = ~(t[21] & t[22]);
  assign t[18] = ~(t[23] & t[24]);
  assign t[19] = ~(t[25] | t[26]);
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = ~(t[27] | t[28]);
  assign t[21] = ~(t[29] | t[49]);
  assign t[22] = ~(t[30] & t[31]);
  assign t[23] = ~(t[50] | t[32]);
  assign t[24] = t[33] & t[49];
  assign t[25] = ~(t[33] | t[34]);
  assign t[26] = ~(t[33] | t[35]);
  assign t[27] = ~(t[33] | t[36]);
  assign t[28] = ~(t[33] | t[37]);
  assign t[29] = ~(t[51]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = ~(t[52] & t[38]);
  assign t[31] = ~(x[4] & t[23]);
  assign t[32] = ~(t[52]);
  assign t[33] = ~(t[29]);
  assign t[34] = t[49] ? t[40] : t[39];
  assign t[35] = t[49] ? t[42] : t[41];
  assign t[36] = t[49] ? t[43] : t[30];
  assign t[37] = t[49] ? t[41] : t[42];
  assign t[38] = ~(x[4] | t[44]);
  assign t[39] = ~(t[45] & t[52]);
  assign t[3] = ~(x[3]);
  assign t[40] = ~(t[46] & t[32]);
  assign t[41] = ~(t[45] & t[32]);
  assign t[42] = ~(t[46] & t[52]);
  assign t[43] = ~(x[4] & t[47]);
  assign t[44] = ~(t[50]);
  assign t[45] = x[4] & t[50];
  assign t[46] = ~(x[4] | t[50]);
  assign t[47] = ~(t[50] | t[52]);
  assign t[48] = t[56] ^ x[2];
  assign t[49] = t[57] ^ x[8];
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[50] = t[58] ^ x[11];
  assign t[51] = t[59] ^ x[14];
  assign t[52] = t[60] ^ x[17];
  assign t[53] = t[61] ^ x[20];
  assign t[54] = t[62] ^ x[25];
  assign t[55] = t[63] ^ x[28];
  assign t[56] = (x[0] & x[1]);
  assign t[57] = (x[6] & x[7]);
  assign t[58] = (x[9] & x[10]);
  assign t[59] = (x[12] & x[13]);
  assign t[5] = t[10] ^ x[5];
  assign t[60] = (x[15] & x[16]);
  assign t[61] = (x[18] & x[19]);
  assign t[62] = (x[23] & x[24]);
  assign t[63] = (x[26] & x[27]);
  assign t[6] = ~(t[49] & t[50]);
  assign t[7] = ~(t[51] & t[52]);
  assign t[8] = ~(t[9] ^ t[11]);
  assign t[9] = ~(t[53] ^ t[12]);
  assign y = t[0] ? t[1] : t[48];
endmodule

module R1ind186(x, y);
 input [37:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[14] ? x[22] : x[21];
  assign t[12] = ~(t[23] ^ t[15]);
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[26] ^ t[27]);
  assign t[16] = ~(t[20]);
  assign t[17] = t[28] ^ x[2];
  assign t[18] = t[29] ^ x[8];
  assign t[19] = t[30] ^ x[11];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[14];
  assign t[21] = t[32] ^ x[17];
  assign t[22] = t[33] ^ x[20];
  assign t[23] = t[34] ^ x[25];
  assign t[24] = t[35] ^ x[28];
  assign t[25] = t[36] ^ x[31];
  assign t[26] = t[37] ^ x[34];
  assign t[27] = t[38] ^ x[37];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[23] & x[24]);
  assign t[35] = (x[26] & x[27]);
  assign t[36] = (x[29] & x[30]);
  assign t[37] = (x[32] & x[33]);
  assign t[38] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[22] ^ t[13]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind187(x, y);
 input [37:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[14] ? x[21] : x[22];
  assign t[12] = ~(t[23] ^ t[15]);
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[26] ^ t[27]);
  assign t[16] = ~(t[20]);
  assign t[17] = t[28] ^ x[2];
  assign t[18] = t[29] ^ x[8];
  assign t[19] = t[30] ^ x[11];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[14];
  assign t[21] = t[32] ^ x[17];
  assign t[22] = t[33] ^ x[20];
  assign t[23] = t[34] ^ x[25];
  assign t[24] = t[35] ^ x[28];
  assign t[25] = t[36] ^ x[31];
  assign t[26] = t[37] ^ x[34];
  assign t[27] = t[38] ^ x[37];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[23] & x[24]);
  assign t[35] = (x[26] & x[27]);
  assign t[36] = (x[29] & x[30]);
  assign t[37] = (x[32] & x[33]);
  assign t[38] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[22] ^ t[13]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind188(x, y);
 input [37:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[14] ? x[21] : x[22];
  assign t[12] = ~(t[23] ^ t[15]);
  assign t[13] = ~(t[24] ^ t[25]);
  assign t[14] = ~(t[16]);
  assign t[15] = ~(t[26] ^ t[27]);
  assign t[16] = ~(t[20]);
  assign t[17] = t[28] ^ x[2];
  assign t[18] = t[29] ^ x[8];
  assign t[19] = t[30] ^ x[11];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[14];
  assign t[21] = t[32] ^ x[17];
  assign t[22] = t[33] ^ x[20];
  assign t[23] = t[34] ^ x[25];
  assign t[24] = t[35] ^ x[28];
  assign t[25] = t[36] ^ x[31];
  assign t[26] = t[37] ^ x[34];
  assign t[27] = t[38] ^ x[37];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[12] & x[13]);
  assign t[32] = (x[15] & x[16]);
  assign t[33] = (x[18] & x[19]);
  assign t[34] = (x[23] & x[24]);
  assign t[35] = (x[26] & x[27]);
  assign t[36] = (x[29] & x[30]);
  assign t[37] = (x[32] & x[33]);
  assign t[38] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[18] & t[19]);
  assign t[7] = ~(t[20] & t[21]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[22] ^ t[13]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind189(x, y);
 input [37:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[60] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[61] ^ t[62]);
  assign t[14] = ~(t[63] & t[64]);
  assign t[15] = ~(t[65] & t[66]);
  assign t[16] = ~(t[67] ^ t[68]);
  assign t[17] = t[65] ? x[9] : x[10];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[21] | t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[27] & t[28]);
  assign t[23] = ~(t[29] | t[30]);
  assign t[24] = t[31] | t[32];
  assign t[25] = ~(t[29]);
  assign t[26] = t[63] ? t[34] : t[33];
  assign t[27] = ~(t[35] | t[36]);
  assign t[28] = ~(t[37] & t[38]);
  assign t[29] = ~(t[65]);
  assign t[2] = ~(t[5]);
  assign t[30] = t[63] ? t[40] : t[39];
  assign t[31] = ~(t[25] | t[41]);
  assign t[32] = ~(t[42]);
  assign t[33] = ~(t[43] & t[66]);
  assign t[34] = ~(t[44] & t[45]);
  assign t[35] = ~(t[25] | t[46]);
  assign t[36] = ~(t[25] | t[47]);
  assign t[37] = t[66] & t[48];
  assign t[38] = t[44] | t[43];
  assign t[39] = ~(x[4] & t[49]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[50] & t[45]);
  assign t[41] = t[63] ? t[52] : t[51];
  assign t[42] = ~(t[48] & t[53]);
  assign t[43] = x[4] & t[64];
  assign t[44] = ~(x[4] | t[64]);
  assign t[45] = ~(t[66]);
  assign t[46] = t[63] ? t[33] : t[34];
  assign t[47] = t[63] ? t[39] : t[54];
  assign t[48] = ~(t[29] | t[63]);
  assign t[49] = ~(t[64] | t[66]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(x[4] | t[55]);
  assign t[51] = ~(t[43] & t[45]);
  assign t[52] = ~(t[44] & t[66]);
  assign t[53] = ~(t[54] & t[56]);
  assign t[54] = ~(t[66] & t[50]);
  assign t[55] = ~(t[64]);
  assign t[56] = ~(x[4] & t[57]);
  assign t[57] = ~(t[64] | t[45]);
  assign t[58] = t[69] ^ x[2];
  assign t[59] = t[70] ^ x[8];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[13];
  assign t[61] = t[72] ^ x[16];
  assign t[62] = t[73] ^ x[19];
  assign t[63] = t[74] ^ x[22];
  assign t[64] = t[75] ^ x[25];
  assign t[65] = t[76] ^ x[28];
  assign t[66] = t[77] ^ x[31];
  assign t[67] = t[78] ^ x[34];
  assign t[68] = t[79] ^ x[37];
  assign t[69] = (x[0] & x[1]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[6] & x[7]);
  assign t[71] = (x[11] & x[12]);
  assign t[72] = (x[14] & x[15]);
  assign t[73] = (x[17] & x[18]);
  assign t[74] = (x[20] & x[21]);
  assign t[75] = (x[23] & x[24]);
  assign t[76] = (x[26] & x[27]);
  assign t[77] = (x[29] & x[30]);
  assign t[78] = (x[32] & x[33]);
  assign t[79] = (x[35] & x[36]);
  assign t[7] = ~(t[59] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[58];
endmodule

module R1ind190(x, y);
 input [37:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[18] ? x[21] : x[22];
  assign t[12] = ~(t[21] ^ t[14]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] ^ t[25]);
  assign t[15] = t[26] ^ x[2];
  assign t[16] = t[27] ^ x[8];
  assign t[17] = t[28] ^ x[11];
  assign t[18] = t[29] ^ x[14];
  assign t[19] = t[30] ^ x[17];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[20];
  assign t[21] = t[32] ^ x[25];
  assign t[22] = t[33] ^ x[28];
  assign t[23] = t[34] ^ x[31];
  assign t[24] = t[35] ^ x[34];
  assign t[25] = t[36] ^ x[37];
  assign t[26] = (x[0] & x[1]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[29] = (x[12] & x[13]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[15] & x[16]);
  assign t[31] = (x[18] & x[19]);
  assign t[32] = (x[23] & x[24]);
  assign t[33] = (x[26] & x[27]);
  assign t[34] = (x[29] & x[30]);
  assign t[35] = (x[32] & x[33]);
  assign t[36] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[16] & t[17]);
  assign t[7] = ~(t[18] & t[19]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[20] ^ t[13]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind191(x, y);
 input [37:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = t[19] ? x[9] : x[10];
  assign t[12] = ~(t[20] ^ t[16]);
  assign t[13] = ~(t[21] ^ t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[19] & t[25]);
  assign t[16] = ~(t[26] ^ t[27]);
  assign t[17] = t[28] ^ x[2];
  assign t[18] = t[29] ^ x[8];
  assign t[19] = t[30] ^ x[13];
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = t[31] ^ x[16];
  assign t[21] = t[32] ^ x[19];
  assign t[22] = t[33] ^ x[22];
  assign t[23] = t[34] ^ x[25];
  assign t[24] = t[35] ^ x[28];
  assign t[25] = t[36] ^ x[31];
  assign t[26] = t[37] ^ x[34];
  assign t[27] = t[38] ^ x[37];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[5]);
  assign t[30] = (x[11] & x[12]);
  assign t[31] = (x[14] & x[15]);
  assign t[32] = (x[17] & x[18]);
  assign t[33] = (x[20] & x[21]);
  assign t[34] = (x[23] & x[24]);
  assign t[35] = (x[26] & x[27]);
  assign t[36] = (x[29] & x[30]);
  assign t[37] = (x[32] & x[33]);
  assign t[38] = (x[35] & x[36]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[4] = t[8] ^ x[5];
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = t[11] ^ t[12];
  assign t[7] = ~(t[18] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[17];
endmodule

module R1ind192(x, y);
 input [37:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = x[21] ^ x[22];
  assign t[11] = t[18] ? x[21] : x[22];
  assign t[12] = ~(t[21] ^ t[14]);
  assign t[13] = ~(t[22] ^ t[23]);
  assign t[14] = ~(t[24] ^ t[25]);
  assign t[15] = t[26] ^ x[2];
  assign t[16] = t[27] ^ x[8];
  assign t[17] = t[28] ^ x[11];
  assign t[18] = t[29] ^ x[14];
  assign t[19] = t[30] ^ x[17];
  assign t[1] = x[3] ? t[5] : t[4];
  assign t[20] = t[31] ^ x[20];
  assign t[21] = t[32] ^ x[25];
  assign t[22] = t[33] ^ x[28];
  assign t[23] = t[34] ^ x[31];
  assign t[24] = t[35] ^ x[34];
  assign t[25] = t[36] ^ x[37];
  assign t[26] = (x[0] & x[1]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[29] = (x[12] & x[13]);
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = (x[15] & x[16]);
  assign t[31] = (x[18] & x[19]);
  assign t[32] = (x[23] & x[24]);
  assign t[33] = (x[26] & x[27]);
  assign t[34] = (x[29] & x[30]);
  assign t[35] = (x[32] & x[33]);
  assign t[36] = (x[35] & x[36]);
  assign t[3] = ~(x[3]);
  assign t[4] = x[4] ? t[9] : t[8];
  assign t[5] = t[10] ^ x[5];
  assign t[6] = ~(t[16] & t[17]);
  assign t[7] = ~(t[18] & t[19]);
  assign t[8] = t[11] ^ t[12];
  assign t[9] = ~(t[20] ^ t[13]);
  assign y = t[0] ? t[1] : t[15];
endmodule

module R1ind193(x, y);
 input [37:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(x[3]);
  assign t[11] = ~(t[56] ^ t[16]);
  assign t[12] = ~(t[17] ^ t[18]);
  assign t[13] = ~(t[57] ^ t[58]);
  assign t[14] = ~(t[59] & t[60]);
  assign t[15] = ~(t[61] & t[62]);
  assign t[16] = ~(t[63] ^ t[64]);
  assign t[17] = t[61] ? x[9] : x[10];
  assign t[18] = ~(t[19] & t[20]);
  assign t[19] = ~(t[21] | t[22]);
  assign t[1] = x[3] ? t[4] : t[3];
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[27] & t[28]);
  assign t[23] = ~(t[25] | t[29]);
  assign t[24] = ~(t[25] | t[30]);
  assign t[25] = ~(t[31]);
  assign t[26] = t[59] ? t[33] : t[32];
  assign t[27] = ~(t[34] | t[35]);
  assign t[28] = ~(t[36] & t[37]);
  assign t[29] = t[59] ? t[39] : t[38];
  assign t[2] = ~(t[5]);
  assign t[30] = t[59] ? t[41] : t[40];
  assign t[31] = ~(t[61]);
  assign t[32] = ~(t[42] & t[62]);
  assign t[33] = ~(t[43] & t[44]);
  assign t[34] = ~(t[25] | t[45]);
  assign t[35] = ~(t[25] | t[46]);
  assign t[36] = t[62] & t[47];
  assign t[37] = t[43] | t[42];
  assign t[38] = ~(t[48] & t[44]);
  assign t[39] = ~(x[4] & t[49]);
  assign t[3] = x[4] ? t[7] : t[6];
  assign t[40] = ~(t[43] & t[62]);
  assign t[41] = ~(t[42] & t[44]);
  assign t[42] = x[4] & t[60];
  assign t[43] = ~(x[4] | t[60]);
  assign t[44] = ~(t[62]);
  assign t[45] = t[59] ? t[32] : t[33];
  assign t[46] = t[59] ? t[51] : t[50];
  assign t[47] = ~(t[31] | t[59]);
  assign t[48] = ~(x[4] | t[52]);
  assign t[49] = ~(t[60] | t[44]);
  assign t[4] = t[8] ^ x[5];
  assign t[50] = ~(t[62] & t[48]);
  assign t[51] = ~(x[4] & t[53]);
  assign t[52] = ~(t[60]);
  assign t[53] = ~(t[60] | t[62]);
  assign t[54] = t[65] ^ x[2];
  assign t[55] = t[66] ^ x[8];
  assign t[56] = t[67] ^ x[13];
  assign t[57] = t[68] ^ x[16];
  assign t[58] = t[69] ^ x[19];
  assign t[59] = t[70] ^ x[22];
  assign t[5] = ~(t[9] & t[10]);
  assign t[60] = t[71] ^ x[25];
  assign t[61] = t[72] ^ x[28];
  assign t[62] = t[73] ^ x[31];
  assign t[63] = t[74] ^ x[34];
  assign t[64] = t[75] ^ x[37];
  assign t[65] = (x[0] & x[1]);
  assign t[66] = (x[6] & x[7]);
  assign t[67] = (x[11] & x[12]);
  assign t[68] = (x[14] & x[15]);
  assign t[69] = (x[17] & x[18]);
  assign t[6] = ~(t[11] ^ t[12]);
  assign t[70] = (x[20] & x[21]);
  assign t[71] = (x[23] & x[24]);
  assign t[72] = (x[26] & x[27]);
  assign t[73] = (x[29] & x[30]);
  assign t[74] = (x[32] & x[33]);
  assign t[75] = (x[35] & x[36]);
  assign t[7] = ~(t[55] ^ t[13]);
  assign t[8] = x[9] ^ x[10];
  assign t[9] = ~(t[14] | t[15]);
  assign y = t[0] ? t[1] : t[54];
endmodule

module R1ind194(x, y);
 input [12:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[10] ^ t[1];
  assign t[10] = t[14] ^ x[3];
  assign t[11] = t[15] ^ x[6];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[12];
  assign t[14] = (x[1] & x[2]);
  assign t[15] = (x[4] & x[5]);
  assign t[16] = (x[7] & x[8]);
  assign t[17] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[11]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[3] = ~(t[12]);
  assign t[4] = ~(t[5] & t[13]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[11] & t[10]);
  assign t[9] = ~(t[13] & t[12]);
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind195(x, y);
 input [12:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = ~(t[9] ^ t[1]);
  assign t[10] = t[14] ^ x[6];
  assign t[11] = t[15] ^ x[9];
  assign t[12] = t[16] ^ x[12];
  assign t[13] = (x[1] & x[2]);
  assign t[14] = (x[4] & x[5]);
  assign t[15] = (x[7] & x[8]);
  assign t[16] = (x[10] & x[11]);
  assign t[1] = ~(t[2] | t[3]);
  assign t[2] = ~(t[10]);
  assign t[3] = ~(t[4] & t[11]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[6] = ~(x[0]);
  assign t[7] = ~(t[9] & t[12]);
  assign t[8] = ~(t[11] & t[10]);
  assign t[9] = t[13] ^ x[3];
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind196(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = t[7] ^ t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & x[2]);
  assign t[12] = (x[4] & x[5]);
  assign t[13] = (x[7] & x[8]);
  assign t[14] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[8]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = ~(t[8] & t[7]);
  assign t[7] = t[11] ^ x[3];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[9];
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind197(x, y);
 input [12:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[6] ^ t[1]);
  assign t[10] = (x[1] & x[2]);
  assign t[11] = (x[4] & x[5]);
  assign t[12] = (x[7] & x[8]);
  assign t[13] = (x[10] & x[11]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(x[0]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[6] & t[9]);
  assign t[6] = t[10] ^ x[3];
  assign t[7] = t[11] ^ x[6];
  assign t[8] = t[12] ^ x[9];
  assign t[9] = t[13] ^ x[12];
  assign y = ~(x[0] | t[0]);
endmodule

module R1ind198(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind199(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind200(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind201(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind202(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind203(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind204(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind205(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind206(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind207(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind208(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind209(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind210(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind211(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind212(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind213(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind214(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind215(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind216(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind217(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind218(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind219(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind220(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind221(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind222(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind223(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind224(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind225(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind226(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind227(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind228(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind229(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind230(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind231(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind232(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind233(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind234(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind235(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind236(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind237(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind238(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind239(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind240(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind241(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind242(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind243(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind244(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind245(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind246(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind247(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind248(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind249(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind250(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind251(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind252(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind253(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind254(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind255(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind256(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind257(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind258(x, y);
 input [8:0] x;
 output y;

 wire [13:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = (x[0] & x[1]);
  assign t[11] = (x[0] & x[3]);
  assign t[12] = (x[0] & x[5]);
  assign t[13] = (x[0] & x[7]);
  assign t[1] = t[4] | t[6];
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[5] | t[2]);
  assign t[5] = ~(t[9]);
  assign t[6] = t[10] ^ x[2];
  assign t[7] = t[11] ^ x[4];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind259(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[4] & t[7]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind260(x, y);
 input [6:0] x;
 output y;

 wire [10:0] t;
  assign t[0] = ~(t[5] & t[2]);
  assign t[10] = (x[0] & x[5]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[2] = ~(t[7]);
  assign t[3] = ~(t[7] & t[4]);
  assign t[4] = ~(t[5]);
  assign t[5] = t[8] ^ x[2];
  assign t[6] = t[9] ^ x[4];
  assign t[7] = t[10] ^ x[6];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[0] & x[3]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind261(x, y);
 input [8:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[14] ^ x[8];
  assign t[11] = (x[0] & x[1]);
  assign t[12] = (x[0] & x[3]);
  assign t[13] = (x[0] & x[5]);
  assign t[14] = (x[0] & x[7]);
  assign t[1] = ~(t[7] | t[4]);
  assign t[2] = ~(t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind262(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind263(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind264(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind265(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind266(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind267(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind268(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind269(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind270(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind271(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind272(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind273(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind274(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind275(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind276(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind277(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind278(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind279(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind280(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind281(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind282(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind283(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind284(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind285(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind286(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind287(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind288(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind289(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind290(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind291(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind292(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind293(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind294(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind295(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind296(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind297(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind298(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind299(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind300(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind301(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind302(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind303(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind304(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind305(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind306(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind307(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind308(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind309(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind310(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind311(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind312(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind313(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind314(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind315(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind316(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind317(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind318(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind319(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind320(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind321(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind322(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind323(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind324(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind325(x, y);
 input [6:0] x;
 output y;

 wire [3:0] t;
  assign t[0] = t[2] ^ x[3];
  assign t[1] = t[3] ^ x[6];
  assign t[2] = (x[1] & x[2]);
  assign t[3] = (x[4] & x[5]);
  assign y = x[0] ? t[1] : t[0];
endmodule

module R1ind326(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind327(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind328(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind329(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind330(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind331(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind332(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind333(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind334(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind335(x, y);
 input [17:0] x;
 output y;

 wire [50:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] & t[17]);
  assign t[11] = ~(t[42]);
  assign t[12] = t[43] ? t[19] : t[18];
  assign t[13] = t[43] ? t[21] : t[20];
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = ~(t[11] & t[24]);
  assign t[16] = ~(t[25] & t[26]);
  assign t[17] = t[11] | t[27];
  assign t[18] = ~(t[28] & t[29]);
  assign t[19] = ~(t[30] & t[29]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(x[11] & t[31]);
  assign t[21] = ~(t[32] & t[29]);
  assign t[22] = ~(t[11] | t[33]);
  assign t[23] = ~(t[34] | t[35]);
  assign t[24] = ~(t[20] & t[36]);
  assign t[25] = t[44] & t[37];
  assign t[26] = t[28] | t[30];
  assign t[27] = t[43] ? t[20] : t[21];
  assign t[28] = ~(x[11] | t[45]);
  assign t[29] = ~(t[44]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = x[11] & t[45];
  assign t[31] = ~(t[45] | t[44]);
  assign t[32] = ~(x[11] | t[38]);
  assign t[33] = t[43] ? t[18] : t[19];
  assign t[34] = ~(t[11]);
  assign t[35] = t[43] ? t[21] : t[39];
  assign t[36] = ~(t[44] & t[32]);
  assign t[37] = ~(t[11] | t[43]);
  assign t[38] = ~(t[45]);
  assign t[39] = ~(x[11] & t[40]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[45] | t[29]);
  assign t[41] = t[46] ^ x[2];
  assign t[42] = t[47] ^ x[7];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = t[49] ^ x[14];
  assign t[45] = t[50] ^ x[17];
  assign t[46] = (x[0] & x[1]);
  assign t[47] = (x[5] & x[6]);
  assign t[48] = (x[8] & x[9]);
  assign t[49] = (x[12] & x[13]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[50] = (x[15] & x[16]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[42]);
  assign t[7] = ~(t[11] | t[12]);
  assign t[8] = ~(t[11] | t[13]);
  assign t[9] = ~(t[14] & t[15]);
  assign y = ~(t[41] ^ t[0]);
endmodule

module R1ind336(x, y);
 input [17:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[36] ? t[18] : t[17];
  assign t[13] = t[36] ? t[20] : t[19];
  assign t[14] = ~(t[16] | t[36]);
  assign t[15] = ~(t[21] | t[22]);
  assign t[16] = ~(t[34]);
  assign t[17] = ~(t[35] & t[23]);
  assign t[18] = ~(x[14] & t[24]);
  assign t[19] = ~(t[25] & t[35]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[26] & t[27]);
  assign t[21] = ~(t[16] | t[28]);
  assign t[22] = ~(t[16] | t[29]);
  assign t[23] = ~(x[14] | t[30]);
  assign t[24] = ~(t[37] | t[35]);
  assign t[25] = ~(x[14] | t[37]);
  assign t[26] = x[14] & t[37];
  assign t[27] = ~(t[35]);
  assign t[28] = t[36] ? t[20] : t[31];
  assign t[29] = t[36] ? t[32] : t[18];
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = ~(t[37]);
  assign t[31] = ~(t[25] & t[27]);
  assign t[32] = ~(t[23] & t[27]);
  assign t[33] = t[38] ^ x[2];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[10];
  assign t[36] = t[41] ^ x[13];
  assign t[37] = t[42] ^ x[17];
  assign t[38] = (x[0] & x[1]);
  assign t[39] = (x[5] & x[6]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[8] & x[9]);
  assign t[41] = (x[11] & x[12]);
  assign t[42] = (x[15] & x[16]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[34]);
  assign t[7] = ~(t[11] | t[12]);
  assign t[8] = ~(t[11] | t[13]);
  assign t[9] = t[35] & t[14];
  assign y = ~(t[33] ^ t[0]);
endmodule

module R1ind337(x, y);
 input [17:0] x;
 output y;

 wire [53:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[15]);
  assign t[11] = t[46] ? t[17] : t[16];
  assign t[12] = ~(t[18] | t[19]);
  assign t[13] = ~(t[20] | t[21]);
  assign t[14] = t[46] ? t[23] : t[22];
  assign t[15] = ~(t[45]);
  assign t[16] = ~(t[24] & t[25]);
  assign t[17] = ~(x[11] & t[26]);
  assign t[18] = ~(t[10] | t[27]);
  assign t[19] = ~(t[28] & t[29]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[15] | t[30]);
  assign t[21] = ~(t[15] | t[31]);
  assign t[22] = ~(t[32] & t[47]);
  assign t[23] = ~(t[33] & t[25]);
  assign t[24] = ~(x[11] | t[34]);
  assign t[25] = ~(t[47]);
  assign t[26] = ~(t[48] | t[25]);
  assign t[27] = t[46] ? t[22] : t[23];
  assign t[28] = ~(t[35] | t[36]);
  assign t[29] = ~(t[15] & t[37]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = t[46] ? t[38] : t[23];
  assign t[31] = t[46] ? t[16] : t[39];
  assign t[32] = x[11] & t[48];
  assign t[33] = ~(x[11] | t[48]);
  assign t[34] = ~(t[48]);
  assign t[35] = ~(t[15] | t[40]);
  assign t[36] = ~(t[10] | t[41]);
  assign t[37] = ~(t[39] & t[42]);
  assign t[38] = ~(t[32] & t[25]);
  assign t[39] = ~(x[11] & t[43]);
  assign t[3] = ~(t[6]);
  assign t[40] = t[46] ? t[23] : t[38];
  assign t[41] = t[46] ? t[16] : t[17];
  assign t[42] = ~(t[47] & t[24]);
  assign t[43] = ~(t[48] | t[47]);
  assign t[44] = t[49] ^ x[2];
  assign t[45] = t[50] ^ x[7];
  assign t[46] = t[51] ^ x[10];
  assign t[47] = t[52] ^ x[14];
  assign t[48] = t[53] ^ x[17];
  assign t[49] = (x[0] & x[1]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[50] = (x[5] & x[6]);
  assign t[51] = (x[8] & x[9]);
  assign t[52] = (x[12] & x[13]);
  assign t[53] = (x[15] & x[16]);
  assign t[5] = ~(t[9]);
  assign t[6] = ~(t[45]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[12] & t[13]);
  assign t[9] = ~(t[10] | t[14]);
  assign y = ~(t[44] ^ t[0]);
endmodule

module R1ind338(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind339(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind340(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind341(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind342(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind343(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind344(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind345(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind346(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind347(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind348(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind349(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind350(x, y);
 input [17:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[16] | t[17];
  assign t[11] = ~(t[15] & t[18]);
  assign t[12] = ~(t[19] & t[20]);
  assign t[13] = ~(t[21] | t[22]);
  assign t[14] = ~(t[21] | t[23]);
  assign t[15] = ~(t[24] | t[37]);
  assign t[16] = ~(x[14] | t[38]);
  assign t[17] = x[14] & t[38];
  assign t[18] = ~(t[25] & t[26]);
  assign t[19] = ~(t[38] | t[27]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = t[21] & t[37];
  assign t[21] = ~(t[24]);
  assign t[22] = t[37] ? t[25] : t[28];
  assign t[23] = t[37] ? t[30] : t[29];
  assign t[24] = ~(t[35]);
  assign t[25] = ~(t[36] & t[31]);
  assign t[26] = ~(x[14] & t[19]);
  assign t[27] = ~(t[36]);
  assign t[28] = ~(x[14] & t[32]);
  assign t[29] = ~(t[17] & t[27]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = ~(t[16] & t[36]);
  assign t[31] = ~(x[14] | t[33]);
  assign t[32] = ~(t[38] | t[36]);
  assign t[33] = ~(t[38]);
  assign t[34] = t[39] ^ x[2];
  assign t[35] = t[40] ^ x[7];
  assign t[36] = t[41] ^ x[10];
  assign t[37] = t[42] ^ x[13];
  assign t[38] = t[43] ^ x[17];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[5] & x[6]);
  assign t[41] = (x[8] & x[9]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[15] & x[16]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = ~(t[35]);
  assign t[7] = ~(t[11] & t[12]);
  assign t[8] = t[13] | t[14];
  assign t[9] = t[36] & t[15];
  assign y = ~(t[34] ^ t[0]);
endmodule

module R1ind351(x, y);
 input [17:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(t[36]);
  assign t[12] = t[37] ? t[18] : t[17];
  assign t[13] = t[37] ? t[20] : t[19];
  assign t[14] = ~(t[21] | t[22]);
  assign t[15] = ~(t[11]);
  assign t[16] = t[37] ? t[23] : t[19];
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[25]);
  assign t[19] = ~(x[11] & t[27]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[28] & t[25]);
  assign t[21] = ~(t[15] | t[29]);
  assign t[22] = ~(t[15] | t[30]);
  assign t[23] = ~(t[38] & t[28]);
  assign t[24] = x[11] & t[39];
  assign t[25] = ~(t[38]);
  assign t[26] = ~(x[11] | t[39]);
  assign t[27] = ~(t[39] | t[38]);
  assign t[28] = ~(x[11] | t[31]);
  assign t[29] = t[37] ? t[32] : t[20];
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = t[37] ? t[17] : t[33];
  assign t[31] = ~(t[39]);
  assign t[32] = ~(x[11] & t[34]);
  assign t[33] = ~(t[26] & t[38]);
  assign t[34] = ~(t[39] | t[25]);
  assign t[35] = t[40] ^ x[2];
  assign t[36] = t[41] ^ x[7];
  assign t[37] = t[42] ^ x[10];
  assign t[38] = t[43] ^ x[14];
  assign t[39] = t[44] ^ x[17];
  assign t[3] = ~(t[6]);
  assign t[40] = (x[0] & x[1]);
  assign t[41] = (x[5] & x[6]);
  assign t[42] = (x[8] & x[9]);
  assign t[43] = (x[12] & x[13]);
  assign t[44] = (x[15] & x[16]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[36]);
  assign t[7] = ~(t[11] | t[12]);
  assign t[8] = ~(t[11] | t[13]);
  assign t[9] = ~(t[14]);
  assign y = ~(t[35] ^ t[0]);
endmodule

module R1ind352(x, y);
 input [17:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[31] ? t[17] : t[16];
  assign t[11] = ~(t[15] | t[18]);
  assign t[12] = ~(t[15] | t[19]);
  assign t[13] = ~(t[32] | t[20]);
  assign t[14] = t[9] & t[31];
  assign t[15] = ~(t[30]);
  assign t[16] = ~(x[14] & t[21]);
  assign t[17] = ~(t[33] & t[22]);
  assign t[18] = t[31] ? t[24] : t[23];
  assign t[19] = t[31] ? t[25] : t[16];
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[32] | t[33]);
  assign t[22] = ~(x[14] | t[26]);
  assign t[23] = ~(t[27] & t[20]);
  assign t[24] = ~(t[28] & t[20]);
  assign t[25] = ~(t[22] & t[20]);
  assign t[26] = ~(t[32]);
  assign t[27] = ~(x[14] | t[32]);
  assign t[28] = x[14] & t[32];
  assign t[29] = t[34] ^ x[2];
  assign t[2] = t[4] | t[5];
  assign t[30] = t[35] ^ x[7];
  assign t[31] = t[36] ^ x[10];
  assign t[32] = t[37] ^ x[13];
  assign t[33] = t[38] ^ x[17];
  assign t[34] = (x[0] & x[1]);
  assign t[35] = (x[5] & x[6]);
  assign t[36] = (x[8] & x[9]);
  assign t[37] = (x[11] & x[12]);
  assign t[38] = (x[15] & x[16]);
  assign t[3] = ~(t[6]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[30]);
  assign t[7] = ~(t[11] | t[12]);
  assign t[8] = ~(t[13] & t[14]);
  assign t[9] = ~(t[15]);
  assign y = ~(t[29] ^ t[0]);
endmodule

module R1ind353(x, y);
 input [17:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[14]);
  assign t[11] = t[36] ? t[16] : t[15];
  assign t[12] = ~(t[17] | t[18]);
  assign t[13] = t[36] ? t[20] : t[19];
  assign t[14] = ~(t[35]);
  assign t[15] = ~(t[21] & t[22]);
  assign t[16] = ~(t[23] & t[37]);
  assign t[17] = ~(t[10] | t[24]);
  assign t[18] = ~(t[10] | t[25]);
  assign t[19] = ~(x[14] & t[26]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[37] & t[27]);
  assign t[21] = ~(x[14] | t[38]);
  assign t[22] = ~(t[37]);
  assign t[23] = x[14] & t[38];
  assign t[24] = t[36] ? t[29] : t[28];
  assign t[25] = t[36] ? t[31] : t[30];
  assign t[26] = ~(t[38] | t[37]);
  assign t[27] = ~(x[14] | t[32]);
  assign t[28] = ~(t[27] & t[22]);
  assign t[29] = ~(x[14] & t[33]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = ~(t[21] & t[37]);
  assign t[31] = ~(t[23] & t[22]);
  assign t[32] = ~(t[38]);
  assign t[33] = ~(t[38] | t[22]);
  assign t[34] = t[39] ^ x[2];
  assign t[35] = t[40] ^ x[7];
  assign t[36] = t[41] ^ x[10];
  assign t[37] = t[42] ^ x[13];
  assign t[38] = t[43] ^ x[17];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[5] & x[6]);
  assign t[41] = (x[8] & x[9]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[15] & x[16]);
  assign t[4] = ~(t[7]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[6] = ~(t[35]);
  assign t[7] = ~(t[10] | t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[10] | t[13]);
  assign y = ~(t[34] ^ t[0]);
endmodule

module R1ind354(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind355(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind356(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind357(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind358(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind359(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind360(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind361(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind362(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind363(x, y);
 input [17:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[40] ? t[17] : t[16];
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = t[40] ? t[23] : t[22];
  assign t[14] = t[40] ? t[25] : t[24];
  assign t[15] = ~(t[39]);
  assign t[16] = ~(t[26] & t[41]);
  assign t[17] = ~(t[27] & t[28]);
  assign t[18] = ~(t[9] | t[29]);
  assign t[19] = ~(t[9] | t[30]);
  assign t[1] = t[39] ? x[7] : x[6];
  assign t[20] = t[41] & t[31];
  assign t[21] = t[27] | t[26];
  assign t[22] = ~(t[32] & t[28]);
  assign t[23] = ~(x[14] & t[33]);
  assign t[24] = ~(t[27] & t[41]);
  assign t[25] = ~(t[26] & t[28]);
  assign t[26] = x[14] & t[42];
  assign t[27] = ~(x[14] | t[42]);
  assign t[28] = ~(t[41]);
  assign t[29] = t[40] ? t[16] : t[17];
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = t[40] ? t[35] : t[34];
  assign t[31] = ~(t[15] | t[40]);
  assign t[32] = ~(x[14] | t[36]);
  assign t[33] = ~(t[42] | t[28]);
  assign t[34] = ~(t[41] & t[32]);
  assign t[35] = ~(x[14] & t[37]);
  assign t[36] = ~(t[42]);
  assign t[37] = ~(t[42] | t[41]);
  assign t[38] = t[43] ^ x[2];
  assign t[39] = t[44] ^ x[5];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[45] ^ x[10];
  assign t[41] = t[46] ^ x[13];
  assign t[42] = t[47] ^ x[17];
  assign t[43] = (x[0] & x[1]);
  assign t[44] = (x[3] & x[4]);
  assign t[45] = (x[8] & x[9]);
  assign t[46] = (x[11] & x[12]);
  assign t[47] = (x[15] & x[16]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[11] & t[12]);
  assign t[7] = ~(t[9] | t[13]);
  assign t[8] = ~(t[9] | t[14]);
  assign t[9] = ~(t[15]);
  assign y = ~(t[38] ^ t[0]);
endmodule

module R1ind364(x, y);
 input [17:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] & t[17]);
  assign t[11] = ~(t[18] & t[19]);
  assign t[12] = ~(t[20]);
  assign t[13] = t[21] | t[22];
  assign t[14] = ~(t[21]);
  assign t[15] = t[38] ? t[24] : t[23];
  assign t[16] = ~(t[21] | t[38]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(t[39] | t[27]);
  assign t[19] = t[14] & t[38];
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[21] | t[28]);
  assign t[21] = ~(t[37]);
  assign t[22] = t[38] ? t[30] : t[29];
  assign t[23] = ~(t[31] & t[40]);
  assign t[24] = ~(t[32] & t[27]);
  assign t[25] = ~(t[40] & t[33]);
  assign t[26] = ~(x[17] & t[18]);
  assign t[27] = ~(t[40]);
  assign t[28] = t[38] ? t[29] : t[30];
  assign t[29] = ~(t[33] & t[27]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = ~(x[17] & t[34]);
  assign t[31] = x[17] & t[39];
  assign t[32] = ~(x[17] | t[39]);
  assign t[33] = ~(x[17] | t[35]);
  assign t[34] = ~(t[39] | t[40]);
  assign t[35] = ~(t[39]);
  assign t[36] = t[41] ^ x[2];
  assign t[37] = t[42] ^ x[7];
  assign t[38] = t[43] ^ x[10];
  assign t[39] = t[44] ^ x[13];
  assign t[3] = ~(t[6]);
  assign t[40] = t[45] ^ x[16];
  assign t[41] = (x[0] & x[1]);
  assign t[42] = (x[5] & x[6]);
  assign t[43] = (x[8] & x[9]);
  assign t[44] = (x[11] & x[12]);
  assign t[45] = (x[14] & x[15]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[5] = ~(t[9]);
  assign t[6] = ~(t[37]);
  assign t[7] = ~(t[10] & t[11]);
  assign t[8] = ~(t[12] & t[13]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = ~(t[36] ^ t[0]);
endmodule

module R1ind365(x, y);
 input [17:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[18] & t[19]);
  assign t[11] = ~(t[39] | t[20]);
  assign t[12] = t[21] & t[38];
  assign t[13] = ~(t[21] | t[22]);
  assign t[14] = ~(t[21] | t[23]);
  assign t[15] = ~(t[21] | t[24]);
  assign t[16] = ~(t[21] | t[25]);
  assign t[17] = ~(t[37]);
  assign t[18] = ~(t[40] & t[26]);
  assign t[19] = ~(x[17] & t[11]);
  assign t[1] = t[37] ? x[7] : x[6];
  assign t[20] = ~(t[40]);
  assign t[21] = ~(t[17]);
  assign t[22] = t[38] ? t[28] : t[27];
  assign t[23] = t[38] ? t[30] : t[29];
  assign t[24] = t[38] ? t[31] : t[18];
  assign t[25] = t[38] ? t[29] : t[30];
  assign t[26] = ~(x[17] | t[32]);
  assign t[27] = ~(t[33] & t[40]);
  assign t[28] = ~(t[34] & t[20]);
  assign t[29] = ~(t[33] & t[20]);
  assign t[2] = t[3] | t[4];
  assign t[30] = ~(t[34] & t[40]);
  assign t[31] = ~(x[17] & t[35]);
  assign t[32] = ~(t[39]);
  assign t[33] = x[17] & t[39];
  assign t[34] = ~(x[17] | t[39]);
  assign t[35] = ~(t[39] | t[40]);
  assign t[36] = t[41] ^ x[2];
  assign t[37] = t[42] ^ x[5];
  assign t[38] = t[43] ^ x[10];
  assign t[39] = t[44] ^ x[13];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[45] ^ x[16];
  assign t[41] = (x[0] & x[1]);
  assign t[42] = (x[3] & x[4]);
  assign t[43] = (x[8] & x[9]);
  assign t[44] = (x[11] & x[12]);
  assign t[45] = (x[14] & x[15]);
  assign t[4] = ~(t[7] & t[8]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = ~(t[11] & t[12]);
  assign t[7] = ~(t[13] | t[14]);
  assign t[8] = ~(t[15] | t[16]);
  assign t[9] = ~(t[17] | t[38]);
  assign y = ~(t[36] ^ t[0]);
endmodule

module R1ind366(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind367(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind368(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind369(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind370(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind371(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind372(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind373(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind374(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind375(x, y);
 input [17:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] & t[17]);
  assign t[11] = ~(t[18]);
  assign t[12] = t[50] ? t[20] : t[19];
  assign t[13] = t[50] ? t[22] : t[21];
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = ~(t[11] | t[25]);
  assign t[16] = ~(t[26] | t[27]);
  assign t[17] = t[18] | t[28];
  assign t[18] = ~(t[49]);
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[31] & t[51]);
  assign t[21] = ~(t[51] & t[32]);
  assign t[22] = ~(x[14] & t[33]);
  assign t[23] = ~(t[34] | t[35]);
  assign t[24] = ~(t[36] & t[37]);
  assign t[25] = t[50] ? t[21] : t[22];
  assign t[26] = ~(t[38]);
  assign t[27] = ~(t[11] | t[39]);
  assign t[28] = t[50] ? t[22] : t[40];
  assign t[29] = ~(x[14] | t[52]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = ~(t[51]);
  assign t[31] = x[14] & t[52];
  assign t[32] = ~(x[14] | t[41]);
  assign t[33] = ~(t[52] | t[51]);
  assign t[34] = ~(t[18] | t[42]);
  assign t[35] = ~(t[18] | t[43]);
  assign t[36] = ~(t[52] | t[30]);
  assign t[37] = t[11] & t[50];
  assign t[38] = ~(t[44] & t[45]);
  assign t[39] = t[50] ? t[46] : t[40];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[32] & t[30]);
  assign t[41] = ~(t[52]);
  assign t[42] = t[50] ? t[47] : t[19];
  assign t[43] = t[50] ? t[40] : t[22];
  assign t[44] = ~(t[18] | t[50]);
  assign t[45] = ~(t[21] & t[46]);
  assign t[46] = ~(x[14] & t[36]);
  assign t[47] = ~(t[31] & t[30]);
  assign t[48] = t[53] ^ x[2];
  assign t[49] = t[54] ^ x[7];
  assign t[4] = ~(t[7] | t[8]);
  assign t[50] = t[55] ^ x[10];
  assign t[51] = t[56] ^ x[13];
  assign t[52] = t[57] ^ x[17];
  assign t[53] = (x[0] & x[1]);
  assign t[54] = (x[5] & x[6]);
  assign t[55] = (x[8] & x[9]);
  assign t[56] = (x[11] & x[12]);
  assign t[57] = (x[15] & x[16]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[49]);
  assign t[7] = ~(t[11] | t[12]);
  assign t[8] = ~(t[11] | t[13]);
  assign t[9] = t[14] | t[15];
  assign y = ~(t[48] ^ t[0]);
endmodule

module R1ind376(x, y);
 input [17:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] & t[17]);
  assign t[11] = ~(t[38]);
  assign t[12] = t[39] ? t[19] : t[18];
  assign t[13] = ~(t[11]);
  assign t[14] = t[39] ? t[21] : t[20];
  assign t[15] = t[39] ? t[22] : t[18];
  assign t[16] = ~(t[23] | t[24]);
  assign t[17] = t[11] | t[25];
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[28] & t[27]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(x[11] & t[29]);
  assign t[21] = ~(t[30] & t[27]);
  assign t[22] = ~(t[28] & t[40]);
  assign t[23] = ~(t[13] | t[31]);
  assign t[24] = ~(t[13] | t[32]);
  assign t[25] = t[39] ? t[33] : t[21];
  assign t[26] = x[11] & t[41];
  assign t[27] = ~(t[40]);
  assign t[28] = ~(x[11] | t[41]);
  assign t[29] = ~(t[41] | t[27]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = ~(x[11] | t[34]);
  assign t[31] = t[39] ? t[35] : t[19];
  assign t[32] = t[39] ? t[18] : t[22];
  assign t[33] = ~(x[11] & t[36]);
  assign t[34] = ~(t[41]);
  assign t[35] = ~(t[26] & t[40]);
  assign t[36] = ~(t[41] | t[40]);
  assign t[37] = t[42] ^ x[2];
  assign t[38] = t[43] ^ x[7];
  assign t[39] = t[44] ^ x[10];
  assign t[3] = ~(t[6]);
  assign t[40] = t[45] ^ x[14];
  assign t[41] = t[46] ^ x[17];
  assign t[42] = (x[0] & x[1]);
  assign t[43] = (x[5] & x[6]);
  assign t[44] = (x[8] & x[9]);
  assign t[45] = (x[12] & x[13]);
  assign t[46] = (x[15] & x[16]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[38]);
  assign t[7] = ~(t[11] | t[12]);
  assign t[8] = ~(t[13] | t[14]);
  assign t[9] = ~(t[13] | t[15]);
  assign y = ~(t[37] ^ t[0]);
endmodule

module R1ind377(x, y);
 input [17:0] x;
 output y;

 wire [52:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[15] | t[17]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = t[20] | t[24];
  assign t[15] = ~(t[20]);
  assign t[16] = t[45] ? t[26] : t[25];
  assign t[17] = t[45] ? t[28] : t[27];
  assign t[18] = ~(t[20] | t[29]);
  assign t[19] = ~(t[15] | t[30]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[44]);
  assign t[21] = ~(t[31] & t[32]);
  assign t[22] = t[46] & t[33];
  assign t[23] = t[34] | t[35];
  assign t[24] = t[45] ? t[31] : t[36];
  assign t[25] = ~(t[34] & t[37]);
  assign t[26] = ~(t[35] & t[46]);
  assign t[27] = ~(t[34] & t[46]);
  assign t[28] = ~(t[35] & t[37]);
  assign t[29] = t[45] ? t[25] : t[28];
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = t[45] ? t[36] : t[38];
  assign t[31] = ~(x[14] & t[39]);
  assign t[32] = ~(t[46] & t[40]);
  assign t[33] = ~(t[20] | t[45]);
  assign t[34] = ~(x[14] | t[47]);
  assign t[35] = x[14] & t[47];
  assign t[36] = ~(t[40] & t[37]);
  assign t[37] = ~(t[46]);
  assign t[38] = ~(x[14] & t[41]);
  assign t[39] = ~(t[47] | t[46]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(x[14] | t[42]);
  assign t[41] = ~(t[47] | t[37]);
  assign t[42] = ~(t[47]);
  assign t[43] = t[48] ^ x[2];
  assign t[44] = t[49] ^ x[7];
  assign t[45] = t[50] ^ x[10];
  assign t[46] = t[51] ^ x[13];
  assign t[47] = t[52] ^ x[17];
  assign t[48] = (x[0] & x[1]);
  assign t[49] = (x[5] & x[6]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[50] = (x[8] & x[9]);
  assign t[51] = (x[11] & x[12]);
  assign t[52] = (x[15] & x[16]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[44]);
  assign t[7] = ~(t[11] & t[12]);
  assign t[8] = ~(t[13] & t[14]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = ~(t[43] ^ t[0]);
endmodule

module R1ind378(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind379(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind380(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind381(x, y);
 input [17:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[11] & t[37];
  assign t[11] = ~(t[16]);
  assign t[12] = t[37] ? t[18] : t[17];
  assign t[13] = ~(t[19] | t[20]);
  assign t[14] = ~(t[16] & t[21]);
  assign t[15] = ~(t[38]);
  assign t[16] = ~(t[35]);
  assign t[17] = ~(t[22] & t[15]);
  assign t[18] = ~(t[23] & t[38]);
  assign t[19] = ~(t[16] | t[24]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[11] | t[25]);
  assign t[21] = ~(t[26] & t[27]);
  assign t[22] = ~(x[17] | t[36]);
  assign t[23] = x[17] & t[36];
  assign t[24] = t[37] ? t[17] : t[28];
  assign t[25] = t[37] ? t[30] : t[29];
  assign t[26] = ~(x[17] & t[31]);
  assign t[27] = ~(t[38] & t[32]);
  assign t[28] = ~(t[23] & t[15]);
  assign t[29] = ~(x[17] & t[9]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = ~(t[32] & t[15]);
  assign t[31] = ~(t[36] | t[38]);
  assign t[32] = ~(x[17] | t[33]);
  assign t[33] = ~(t[36]);
  assign t[34] = t[39] ^ x[2];
  assign t[35] = t[40] ^ x[7];
  assign t[36] = t[41] ^ x[10];
  assign t[37] = t[42] ^ x[13];
  assign t[38] = t[43] ^ x[16];
  assign t[39] = (x[0] & x[1]);
  assign t[3] = ~(t[6]);
  assign t[40] = (x[5] & x[6]);
  assign t[41] = (x[8] & x[9]);
  assign t[42] = (x[11] & x[12]);
  assign t[43] = (x[14] & x[15]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[5] = ~(t[9] & t[10]);
  assign t[6] = ~(t[35]);
  assign t[7] = ~(t[11] | t[12]);
  assign t[8] = ~(t[13] & t[14]);
  assign t[9] = ~(t[36] | t[15]);
  assign y = ~(t[34] ^ t[0]);
endmodule

module R1ind382(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind383(x, y);
 input [7:0] x;
 output y;

 wire [4:0] t;
  assign t[0] = t[2] ? x[7] : x[6];
  assign t[1] = t[3] ^ x[2];
  assign t[2] = t[4] ^ x[5];
  assign t[3] = (x[0] & x[1]);
  assign t[4] = (x[3] & x[4]);
  assign y = t[0] ^ t[1];
endmodule

module R1ind384(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind385(x, y);
 input [17:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = ~(t[16] & t[17]);
  assign t[11] = ~(t[14]);
  assign t[12] = t[38] ? t[19] : t[18];
  assign t[13] = t[38] ? t[21] : t[20];
  assign t[14] = ~(t[37]);
  assign t[15] = t[38] ? t[19] : t[20];
  assign t[16] = ~(t[22] | t[23]);
  assign t[17] = ~(t[24] & t[25]);
  assign t[18] = ~(t[26] & t[39]);
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = t[3] ? x[4] : x[3];
  assign t[20] = ~(t[26] & t[28]);
  assign t[21] = ~(t[27] & t[39]);
  assign t[22] = ~(t[14] | t[29]);
  assign t[23] = ~(t[14] | t[30]);
  assign t[24] = ~(t[40] | t[28]);
  assign t[25] = t[11] & t[38];
  assign t[26] = x[17] & t[40];
  assign t[27] = ~(x[17] | t[40]);
  assign t[28] = ~(t[39]);
  assign t[29] = t[38] ? t[20] : t[19];
  assign t[2] = ~(t[4] & t[5]);
  assign t[30] = t[38] ? t[32] : t[31];
  assign t[31] = ~(x[17] & t[33]);
  assign t[32] = ~(t[34] & t[28]);
  assign t[33] = ~(t[40] | t[39]);
  assign t[34] = ~(x[17] | t[35]);
  assign t[35] = ~(t[40]);
  assign t[36] = t[41] ^ x[2];
  assign t[37] = t[42] ^ x[7];
  assign t[38] = t[43] ^ x[10];
  assign t[39] = t[44] ^ x[13];
  assign t[3] = ~(t[6]);
  assign t[40] = t[45] ^ x[16];
  assign t[41] = (x[0] & x[1]);
  assign t[42] = (x[5] & x[6]);
  assign t[43] = (x[8] & x[9]);
  assign t[44] = (x[11] & x[12]);
  assign t[45] = (x[14] & x[15]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[37]);
  assign t[7] = ~(t[11] | t[12]);
  assign t[8] = ~(t[11] | t[13]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = ~(t[36] ^ t[0]);
endmodule

module R1ind386(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind387(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind388(x, y);
 input [7:0] x;
 output y;

 wire [6:0] t;
  assign t[0] = t[1] ? x[4] : x[3];
  assign t[1] = ~(t[2]);
  assign t[2] = ~(t[4]);
  assign t[3] = t[5] ^ x[2];
  assign t[4] = t[6] ^ x[7];
  assign t[5] = (x[0] & x[1]);
  assign t[6] = (x[5] & x[6]);
  assign y = t[0] ^ t[3];
endmodule

module R1ind389(x, y);
 input [17:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] ^ t[2]);
  assign t[10] = t[44] ? t[18] : t[17];
  assign t[11] = ~(t[19] | t[20]);
  assign t[12] = ~(t[21] & t[22]);
  assign t[13] = ~(t[43]);
  assign t[14] = t[44] ? t[24] : t[23];
  assign t[15] = ~(t[9] | t[25]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[27] & t[45]);
  assign t[18] = ~(t[28] & t[29]);
  assign t[19] = ~(t[9] | t[30]);
  assign t[1] = t[43] ? x[7] : x[6];
  assign t[20] = ~(t[9] | t[31]);
  assign t[21] = t[45] & t[32];
  assign t[22] = t[28] | t[27];
  assign t[23] = ~(x[14] & t[33]);
  assign t[24] = ~(t[34] & t[29]);
  assign t[25] = t[44] ? t[36] : t[35];
  assign t[26] = ~(t[32] & t[37]);
  assign t[27] = x[14] & t[46];
  assign t[28] = ~(x[14] | t[46]);
  assign t[29] = ~(t[45]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = t[44] ? t[17] : t[18];
  assign t[31] = t[44] ? t[23] : t[38];
  assign t[32] = ~(t[13] | t[44]);
  assign t[33] = ~(t[46] | t[45]);
  assign t[34] = ~(x[14] | t[39]);
  assign t[35] = ~(t[27] & t[29]);
  assign t[36] = ~(t[28] & t[45]);
  assign t[37] = ~(t[38] & t[40]);
  assign t[38] = ~(t[45] & t[34]);
  assign t[39] = ~(t[46]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = ~(x[14] & t[41]);
  assign t[41] = ~(t[46] | t[29]);
  assign t[42] = t[47] ^ x[2];
  assign t[43] = t[48] ^ x[5];
  assign t[44] = t[49] ^ x[10];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[17];
  assign t[47] = (x[0] & x[1]);
  assign t[48] = (x[3] & x[4]);
  assign t[49] = (x[8] & x[9]);
  assign t[4] = ~(t[7] | t[8]);
  assign t[50] = (x[11] & x[12]);
  assign t[51] = (x[15] & x[16]);
  assign t[5] = ~(t[9] | t[10]);
  assign t[6] = ~(t[11] & t[12]);
  assign t[7] = ~(t[13] | t[14]);
  assign t[8] = t[15] | t[16];
  assign t[9] = ~(t[13]);
  assign y = ~(t[42] ^ t[0]);
endmodule

module R1_ind(x, y);
 input [928:0] x;
 output [389:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[7], x[6], x[3]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[9], x[8], x[3]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[11], x[10], x[3]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[14], x[13], x[12]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[16], x[15], x[12]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[18], x[17], x[12]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[20], x[19], x[12]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[23], x[22], x[21]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[25], x[24], x[21]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[27], x[26], x[21]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[29], x[28], x[21]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[32], x[31], x[30]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[34], x[33], x[30]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[36], x[35], x[30]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[38], x[37], x[30]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[41], x[40], x[39]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[43], x[42], x[39]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[45], x[44], x[39]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[47], x[46], x[39]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[50], x[49], x[48]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[52], x[51], x[48]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[54], x[53], x[48]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[56], x[55], x[48]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[59], x[58], x[57]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[61], x[60], x[57]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[63], x[62], x[57]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[65], x[64], x[57]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[68], x[67], x[66]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[70], x[69], x[66]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[72], x[71], x[66]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[74], x[73], x[66]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[77], x[76], x[75]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[79], x[78], x[75]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[81], x[80], x[75]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[83], x[82], x[75]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[86], x[85], x[84]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[88], x[87], x[84]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[90], x[89], x[84]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[92], x[91], x[84]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[95], x[94], x[93]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[97], x[96], x[93]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[99], x[98], x[93]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[101], x[100], x[93]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[104], x[103], x[102]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[106], x[105], x[102]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[108], x[107], x[102]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[110], x[109], x[102]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[113], x[112], x[111]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[115], x[114], x[111]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[117], x[116], x[111]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[119], x[118], x[111]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[122], x[121], x[120]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[124], x[123], x[120]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[126], x[125], x[120]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[128], x[127], x[120]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[131], x[130], x[129]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[133], x[132], x[129]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[135], x[134], x[129]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[137], x[136], x[129]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[140], x[139], x[138]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[142], x[141], x[138]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[144], x[143], x[138]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[146], x[145], x[138]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[151], x[150], x[149], x[148], x[147]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[155], x[154], x[153], x[152], x[147]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[159], x[158], x[157], x[156], x[147]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[163], x[162], x[161], x[160], x[147]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[168], x[167], x[166], x[165], x[164]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[172], x[171], x[170], x[169], x[164]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[176], x[175], x[174], x[173], x[164]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[180], x[179], x[178], x[177], x[164]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[185], x[184], x[183], x[182], x[181]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[189], x[188], x[187], x[186], x[181]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[193], x[192], x[191], x[190], x[181]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[197], x[196], x[195], x[194], x[181]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[202], x[201], x[200], x[199], x[198]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[206], x[205], x[204], x[203], x[198]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[210], x[209], x[208], x[207], x[198]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[214], x[213], x[212], x[211], x[198]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[219], x[218], x[217], x[216], x[215]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[223], x[222], x[221], x[220], x[215]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[227], x[226], x[225], x[224], x[215]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[231], x[230], x[229], x[228], x[215]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[236], x[235], x[234], x[233], x[232]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[240], x[239], x[238], x[237], x[232]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[244], x[243], x[242], x[241], x[232]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[248], x[247], x[246], x[245], x[232]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[253], x[252], x[251], x[250], x[249]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[257], x[256], x[255], x[254], x[249]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[261], x[260], x[259], x[258], x[249]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[265], x[264], x[263], x[262], x[249]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[270], x[269], x[268], x[267], x[266]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[274], x[273], x[272], x[271], x[266]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[278], x[277], x[276], x[275], x[266]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[282], x[281], x[280], x[279], x[266]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[287], x[286], x[285], x[284], x[283]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[291], x[290], x[289], x[288], x[283]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[295], x[294], x[293], x[292], x[283]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[299], x[298], x[297], x[296], x[283]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[304], x[303], x[302], x[301], x[300]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[308], x[307], x[306], x[305], x[300]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[312], x[311], x[310], x[309], x[300]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[316], x[315], x[314], x[313], x[300]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[321], x[320], x[319], x[318], x[317]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[325], x[324], x[323], x[322], x[317]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[329], x[328], x[327], x[326], x[317]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[333], x[332], x[331], x[330], x[317]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[338], x[337], x[336], x[335], x[334]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[342], x[341], x[340], x[339], x[334]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[346], x[345], x[344], x[343], x[334]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[350], x[349], x[348], x[347], x[334]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[355], x[354], x[353], x[352], x[351]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[359], x[358], x[357], x[356], x[351]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[363], x[362], x[361], x[360], x[351]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[367], x[366], x[365], x[364], x[351]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[372], x[371], x[370], x[369], x[368]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[376], x[375], x[374], x[373], x[368]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[380], x[379], x[378], x[377], x[368]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[384], x[383], x[382], x[381], x[368]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[389], x[388], x[387], x[386], x[385]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[393], x[392], x[391], x[390], x[385]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[397], x[396], x[395], x[394], x[385]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[401], x[400], x[399], x[398], x[385]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[406], x[405], x[404], x[403], x[402]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[410], x[409], x[408], x[407], x[402]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[414], x[413], x[412], x[411], x[402]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[418], x[417], x[416], x[415], x[402]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[445], x[444], x[443], x[442], x[441], x[440], x[151], x[150], x[439], x[438], x[437], x[436], x[435], x[434], x[433], x[432], x[431]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[454], x[453], x[443], x[452], x[451], x[440], x[155], x[154], x[450], x[449], x[437], x[448], x[435], x[434], x[447], x[446], x[431]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[463], x[462], x[443], x[461], x[460], x[440], x[159], x[158], x[459], x[458], x[437], x[457], x[435], x[434], x[456], x[455], x[431]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[472], x[471], x[440], x[470], x[469], x[443], x[163], x[162], x[468], x[467], x[437], x[466], x[435], x[434], x[465], x[464], x[431]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[445], x[444], x[443], x[442], x[441], x[440], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[488], x[487], x[486], x[485], x[484], x[483], x[482], x[481], x[480], x[168], x[167], x[479], x[478], x[477], x[476], x[435], x[434], x[475], x[474], x[473]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[454], x[453], x[443], x[452], x[451], x[440], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[499], x[498], x[486], x[497], x[496], x[483], x[495], x[494], x[480], x[172], x[171], x[493], x[492], x[477], x[491], x[435], x[434], x[490], x[489], x[473]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[463], x[462], x[443], x[461], x[460], x[440], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[510], x[509], x[483], x[508], x[507], x[486], x[506], x[505], x[480], x[176], x[175], x[504], x[503], x[477], x[502], x[435], x[434], x[501], x[500], x[473]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[472], x[471], x[440], x[470], x[469], x[443], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[521], x[520], x[486], x[519], x[518], x[483], x[517], x[516], x[480], x[180], x[179], x[515], x[514], x[477], x[513], x[435], x[434], x[512], x[511], x[473]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[439], x[438], x[437], x[482], x[481], x[480], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[534], x[533], x[532], x[531], x[530], x[529], x[442], x[441], x[440], x[185], x[184], x[528], x[527], x[526], x[525], x[435], x[434], x[524], x[523], x[522]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[450], x[449], x[437], x[495], x[494], x[480], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[543], x[542], x[532], x[541], x[540], x[529], x[452], x[451], x[440], x[189], x[188], x[539], x[538], x[526], x[537], x[435], x[434], x[536], x[535], x[522]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[506], x[505], x[480], x[459], x[458], x[437], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[552], x[551], x[529], x[550], x[549], x[532], x[461], x[460], x[440], x[193], x[192], x[548], x[547], x[526], x[546], x[435], x[434], x[545], x[544], x[522]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[468], x[467], x[437], x[517], x[516], x[480], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[561], x[560], x[532], x[559], x[558], x[529], x[472], x[471], x[440], x[197], x[196], x[557], x[556], x[526], x[555], x[435], x[434], x[554], x[553], x[522]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[439], x[438], x[437], x[482], x[481], x[480], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[574], x[573], x[572], x[571], x[570], x[569], x[445], x[444], x[443], x[202], x[201], x[568], x[567], x[566], x[565], x[435], x[434], x[564], x[563], x[562]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[450], x[449], x[437], x[495], x[494], x[480], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[583], x[582], x[572], x[581], x[580], x[569], x[454], x[453], x[443], x[206], x[205], x[579], x[578], x[566], x[577], x[435], x[434], x[576], x[575], x[562]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[506], x[505], x[480], x[459], x[458], x[437], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[592], x[591], x[572], x[590], x[589], x[569], x[463], x[462], x[443], x[210], x[209], x[588], x[587], x[566], x[586], x[435], x[434], x[585], x[584], x[562]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[468], x[467], x[437], x[517], x[516], x[480], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[601], x[600], x[569], x[599], x[598], x[572], x[470], x[469], x[443], x[214], x[213], x[597], x[596], x[566], x[595], x[435], x[434], x[594], x[593], x[562]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[479], x[478], x[477], x[608], x[607], x[606], x[488], x[487], x[486], x[219], x[218], x[485], x[484], x[483], x[605], x[435], x[434], x[604], x[603], x[602]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[493], x[492], x[477], x[613], x[612], x[606], x[499], x[498], x[486], x[223], x[222], x[497], x[496], x[483], x[611], x[435], x[434], x[610], x[609], x[602]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[504], x[503], x[477], x[618], x[617], x[606], x[508], x[507], x[486], x[227], x[226], x[510], x[509], x[483], x[616], x[435], x[434], x[615], x[614], x[602]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[623], x[622], x[606], x[515], x[514], x[477], x[521], x[520], x[486], x[231], x[230], x[519], x[518], x[483], x[621], x[435], x[434], x[620], x[619], x[602]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[479], x[478], x[477], x[608], x[607], x[606], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[439], x[438], x[437], x[482], x[481], x[480], x[485], x[484], x[483], x[236], x[235], x[442], x[441], x[440], x[627], x[435], x[434], x[626], x[625], x[624]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[493], x[492], x[477], x[613], x[612], x[606], x[450], x[449], x[437], x[495], x[494], x[480], x[497], x[496], x[483], x[240], x[239], x[452], x[451], x[440], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[630], x[435], x[434], x[629], x[628], x[624]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[504], x[503], x[477], x[618], x[617], x[606], x[506], x[505], x[480], x[459], x[458], x[437], x[510], x[509], x[483], x[244], x[243], x[461], x[460], x[440], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[633], x[435], x[434], x[632], x[631], x[624]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[623], x[622], x[606], x[515], x[514], x[477], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[468], x[467], x[437], x[517], x[516], x[480], x[519], x[518], x[483], x[248], x[247], x[472], x[471], x[440], x[636], x[435], x[434], x[635], x[634], x[624]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[488], x[487], x[486], x[485], x[484], x[483], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[643], x[642], x[641], x[568], x[567], x[566], x[608], x[607], x[606], x[253], x[252], x[574], x[573], x[572], x[640], x[435], x[434], x[639], x[638], x[637]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[499], x[498], x[486], x[497], x[496], x[483], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[648], x[647], x[641], x[579], x[578], x[566], x[613], x[612], x[606], x[257], x[256], x[583], x[582], x[572], x[646], x[435], x[434], x[645], x[644], x[637]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[510], x[509], x[483], x[508], x[507], x[486], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[588], x[587], x[566], x[653], x[652], x[641], x[618], x[617], x[606], x[261], x[260], x[592], x[591], x[572], x[651], x[435], x[434], x[650], x[649], x[637]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[521], x[520], x[486], x[519], x[518], x[483], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[658], x[657], x[641], x[597], x[596], x[566], x[623], x[622], x[606], x[265], x[264], x[599], x[598], x[572], x[656], x[435], x[434], x[655], x[654], x[637]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[488], x[487], x[486], x[485], x[484], x[483], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[665], x[664], x[663], x[528], x[527], x[526], x[479], x[478], x[477], x[270], x[269], x[534], x[533], x[532], x[662], x[435], x[434], x[661], x[660], x[659]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[499], x[498], x[486], x[497], x[496], x[483], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[670], x[669], x[663], x[539], x[538], x[526], x[493], x[492], x[477], x[274], x[273], x[543], x[542], x[532], x[668], x[435], x[434], x[667], x[666], x[659]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[510], x[509], x[483], x[508], x[507], x[486], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[675], x[674], x[663], x[548], x[547], x[526], x[504], x[503], x[477], x[278], x[277], x[550], x[549], x[532], x[673], x[435], x[434], x[672], x[671], x[659]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[521], x[520], x[486], x[519], x[518], x[483], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[557], x[556], x[526], x[680], x[679], x[663], x[515], x[514], x[477], x[282], x[281], x[561], x[560], x[532], x[678], x[435], x[434], x[677], x[676], x[659]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[574], x[573], x[572], x[571], x[570], x[569], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[534], x[533], x[532], x[531], x[530], x[529], x[643], x[642], x[641], x[287], x[286], x[665], x[664], x[663], x[684], x[435], x[434], x[683], x[682], x[681]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[583], x[582], x[572], x[581], x[580], x[569], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[543], x[542], x[532], x[541], x[540], x[529], x[648], x[647], x[641], x[291], x[290], x[670], x[669], x[663], x[687], x[435], x[434], x[686], x[685], x[681]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[592], x[591], x[572], x[590], x[589], x[569], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[552], x[551], x[529], x[550], x[549], x[532], x[653], x[652], x[641], x[295], x[294], x[675], x[674], x[663], x[690], x[435], x[434], x[689], x[688], x[681]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[601], x[600], x[569], x[599], x[598], x[572], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[561], x[560], x[532], x[559], x[558], x[529], x[658], x[657], x[641], x[299], x[298], x[680], x[679], x[663], x[693], x[435], x[434], x[692], x[691], x[681]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[574], x[573], x[572], x[571], x[570], x[569], x[568], x[567], x[566], x[304], x[303], x[643], x[642], x[641], x[697], x[435], x[434], x[696], x[695], x[694]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[430], x[429], x[428], x[424], x[423], x[422], x[421], x[420], x[419], x[583], x[582], x[572], x[581], x[580], x[569], x[579], x[578], x[566], x[427], x[426], x[425], x[308], x[307], x[648], x[647], x[641], x[700], x[435], x[434], x[699], x[698], x[694]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[592], x[591], x[572], x[590], x[589], x[569], x[588], x[587], x[566], x[312], x[311], x[653], x[652], x[641], x[703], x[435], x[434], x[702], x[701], x[694]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[601], x[600], x[569], x[599], x[598], x[572], x[597], x[596], x[566], x[316], x[315], x[658], x[657], x[641], x[706], x[435], x[434], x[705], x[704], x[694]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[643], x[642], x[641], x[568], x[567], x[566], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[445], x[444], x[443], x[442], x[441], x[440], x[571], x[570], x[569], x[321], x[320], x[482], x[481], x[480], x[710], x[435], x[434], x[709], x[708], x[707]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[648], x[647], x[641], x[579], x[578], x[566], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[454], x[453], x[443], x[452], x[451], x[440], x[581], x[580], x[569], x[325], x[324], x[495], x[494], x[480], x[713], x[435], x[434], x[712], x[711], x[707]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[588], x[587], x[566], x[653], x[652], x[641], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[463], x[462], x[443], x[461], x[460], x[440], x[590], x[589], x[569], x[329], x[328], x[506], x[505], x[480], x[716], x[435], x[434], x[715], x[714], x[707]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[658], x[657], x[641], x[597], x[596], x[566], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[472], x[471], x[440], x[470], x[469], x[443], x[601], x[600], x[569], x[333], x[332], x[517], x[516], x[480], x[719], x[435], x[434], x[718], x[717], x[707]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[643], x[642], x[641], x[568], x[567], x[566], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[488], x[487], x[486], x[485], x[484], x[483], x[574], x[573], x[572], x[338], x[337], x[608], x[607], x[606], x[723], x[435], x[434], x[722], x[721], x[720]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[648], x[647], x[641], x[579], x[578], x[566], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[499], x[498], x[486], x[497], x[496], x[483], x[583], x[582], x[572], x[342], x[341], x[613], x[612], x[606], x[726], x[435], x[434], x[725], x[724], x[720]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[588], x[587], x[566], x[653], x[652], x[641], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[510], x[509], x[483], x[508], x[507], x[486], x[592], x[591], x[572], x[346], x[345], x[618], x[617], x[606], x[729], x[435], x[434], x[728], x[727], x[720]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[658], x[657], x[641], x[597], x[596], x[566], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[521], x[520], x[486], x[519], x[518], x[483], x[599], x[598], x[572], x[350], x[349], x[623], x[622], x[606], x[732], x[435], x[434], x[731], x[730], x[720]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[665], x[664], x[663], x[528], x[527], x[526], x[643], x[642], x[641], x[568], x[567], x[566], x[534], x[533], x[532], x[355], x[354], x[571], x[570], x[569], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[736], x[435], x[434], x[735], x[734], x[733]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[670], x[669], x[663], x[539], x[538], x[526], x[648], x[647], x[641], x[579], x[578], x[566], x[543], x[542], x[532], x[359], x[358], x[581], x[580], x[569], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[739], x[435], x[434], x[738], x[737], x[733]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[675], x[674], x[663], x[548], x[547], x[526], x[588], x[587], x[566], x[653], x[652], x[641], x[550], x[549], x[532], x[363], x[362], x[590], x[589], x[569], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[742], x[435], x[434], x[741], x[740], x[733]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[557], x[556], x[526], x[680], x[679], x[663], x[658], x[657], x[641], x[597], x[596], x[566], x[561], x[560], x[532], x[367], x[366], x[601], x[600], x[569], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[745], x[435], x[434], x[744], x[743], x[733]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[665], x[664], x[663], x[528], x[527], x[526], x[372], x[371], x[531], x[530], x[529], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[749], x[435], x[434], x[748], x[747], x[746]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[670], x[669], x[663], x[539], x[538], x[526], x[376], x[375], x[541], x[540], x[529], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[752], x[435], x[434], x[751], x[750], x[746]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[675], x[674], x[663], x[548], x[547], x[526], x[380], x[379], x[552], x[551], x[529], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[755], x[435], x[434], x[754], x[753], x[746]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[557], x[556], x[526], x[680], x[679], x[663], x[384], x[383], x[559], x[558], x[529], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[758], x[435], x[434], x[757], x[756], x[746]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[534], x[533], x[532], x[531], x[530], x[529], x[479], x[478], x[477], x[608], x[607], x[606], x[528], x[527], x[526], x[389], x[388], x[488], x[487], x[486], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[762], x[435], x[434], x[761], x[760], x[759]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[543], x[542], x[532], x[541], x[540], x[529], x[493], x[492], x[477], x[613], x[612], x[606], x[539], x[538], x[526], x[393], x[392], x[499], x[498], x[486], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[765], x[435], x[434], x[764], x[763], x[759]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[552], x[551], x[529], x[550], x[549], x[532], x[504], x[503], x[477], x[618], x[617], x[606], x[548], x[547], x[526], x[397], x[396], x[508], x[507], x[486], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[768], x[435], x[434], x[767], x[766], x[759]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[561], x[560], x[532], x[559], x[558], x[529], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[623], x[622], x[606], x[515], x[514], x[477], x[557], x[556], x[526], x[401], x[400], x[521], x[520], x[486], x[771], x[435], x[434], x[770], x[769], x[759]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[534], x[533], x[532], x[531], x[530], x[529], x[439], x[438], x[437], x[482], x[481], x[480], x[665], x[664], x[663], x[406], x[405], x[445], x[444], x[443], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[775], x[435], x[434], x[774], x[773], x[772]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[543], x[542], x[532], x[541], x[540], x[529], x[430], x[429], x[428], x[424], x[423], x[422], x[421], x[420], x[419], x[450], x[449], x[437], x[495], x[494], x[480], x[670], x[669], x[663], x[427], x[426], x[425], x[410], x[409], x[454], x[453], x[443], x[778], x[435], x[434], x[777], x[776], x[772]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[552], x[551], x[529], x[550], x[549], x[532], x[506], x[505], x[480], x[459], x[458], x[437], x[675], x[674], x[663], x[414], x[413], x[463], x[462], x[443], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[781], x[435], x[434], x[780], x[779], x[772]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[561], x[560], x[532], x[559], x[558], x[529], x[430], x[429], x[428], x[427], x[426], x[425], x[424], x[423], x[422], x[421], x[420], x[419], x[468], x[467], x[437], x[517], x[516], x[480], x[680], x[679], x[663], x[418], x[417], x[470], x[469], x[443], x[784], x[435], x[434], x[783], x[782], x[772]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[427], x[426], x[425], x[430], x[429], x[428], x[421], x[420], x[419], x[424], x[423], x[422], x[434]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[424], x[423], x[422], x[427], x[426], x[425], x[430], x[429], x[428], x[421], x[420], x[419], x[434]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[424], x[423], x[422], x[421], x[420], x[419], x[427], x[426], x[425], x[430], x[429], x[428], x[434]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[430], x[429], x[428], x[424], x[423], x[422], x[421], x[420], x[419], x[427], x[426], x[425], x[434]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[447], x[446], x[465], x[464], x[433], x[432], x[456], x[455], x[431]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[447], x[446], x[465], x[464], x[433], x[432], x[456], x[455], x[431]}), .y(y[199]));
  R1ind200 R1ind200_inst(.x({x[433], x[432], x[465], x[464], x[447], x[446], x[431]}), .y(y[200]));
  R1ind201 R1ind201_inst(.x({x[465], x[464], x[433], x[432], x[447], x[446], x[456], x[455], x[431]}), .y(y[201]));
  R1ind202 R1ind202_inst(.x({x[490], x[489], x[512], x[511], x[475], x[474], x[501], x[500], x[473]}), .y(y[202]));
  R1ind203 R1ind203_inst(.x({x[490], x[489], x[512], x[511], x[475], x[474], x[501], x[500], x[473]}), .y(y[203]));
  R1ind204 R1ind204_inst(.x({x[475], x[474], x[512], x[511], x[490], x[489], x[473]}), .y(y[204]));
  R1ind205 R1ind205_inst(.x({x[512], x[511], x[475], x[474], x[490], x[489], x[501], x[500], x[473]}), .y(y[205]));
  R1ind206 R1ind206_inst(.x({x[536], x[535], x[554], x[553], x[524], x[523], x[545], x[544], x[522]}), .y(y[206]));
  R1ind207 R1ind207_inst(.x({x[536], x[535], x[554], x[553], x[524], x[523], x[545], x[544], x[522]}), .y(y[207]));
  R1ind208 R1ind208_inst(.x({x[524], x[523], x[554], x[553], x[536], x[535], x[522]}), .y(y[208]));
  R1ind209 R1ind209_inst(.x({x[554], x[553], x[524], x[523], x[536], x[535], x[545], x[544], x[522]}), .y(y[209]));
  R1ind210 R1ind210_inst(.x({x[576], x[575], x[594], x[593], x[564], x[563], x[585], x[584], x[562]}), .y(y[210]));
  R1ind211 R1ind211_inst(.x({x[576], x[575], x[594], x[593], x[564], x[563], x[585], x[584], x[562]}), .y(y[211]));
  R1ind212 R1ind212_inst(.x({x[564], x[563], x[594], x[593], x[576], x[575], x[562]}), .y(y[212]));
  R1ind213 R1ind213_inst(.x({x[594], x[593], x[564], x[563], x[576], x[575], x[585], x[584], x[562]}), .y(y[213]));
  R1ind214 R1ind214_inst(.x({x[610], x[609], x[620], x[619], x[604], x[603], x[615], x[614], x[602]}), .y(y[214]));
  R1ind215 R1ind215_inst(.x({x[610], x[609], x[620], x[619], x[604], x[603], x[615], x[614], x[602]}), .y(y[215]));
  R1ind216 R1ind216_inst(.x({x[604], x[603], x[620], x[619], x[610], x[609], x[602]}), .y(y[216]));
  R1ind217 R1ind217_inst(.x({x[620], x[619], x[604], x[603], x[610], x[609], x[615], x[614], x[602]}), .y(y[217]));
  R1ind218 R1ind218_inst(.x({x[629], x[628], x[635], x[634], x[626], x[625], x[632], x[631], x[624]}), .y(y[218]));
  R1ind219 R1ind219_inst(.x({x[629], x[628], x[635], x[634], x[626], x[625], x[632], x[631], x[624]}), .y(y[219]));
  R1ind220 R1ind220_inst(.x({x[626], x[625], x[635], x[634], x[629], x[628], x[624]}), .y(y[220]));
  R1ind221 R1ind221_inst(.x({x[635], x[634], x[626], x[625], x[629], x[628], x[632], x[631], x[624]}), .y(y[221]));
  R1ind222 R1ind222_inst(.x({x[645], x[644], x[655], x[654], x[639], x[638], x[650], x[649], x[637]}), .y(y[222]));
  R1ind223 R1ind223_inst(.x({x[645], x[644], x[655], x[654], x[639], x[638], x[650], x[649], x[637]}), .y(y[223]));
  R1ind224 R1ind224_inst(.x({x[639], x[638], x[655], x[654], x[645], x[644], x[637]}), .y(y[224]));
  R1ind225 R1ind225_inst(.x({x[655], x[654], x[639], x[638], x[645], x[644], x[650], x[649], x[637]}), .y(y[225]));
  R1ind226 R1ind226_inst(.x({x[667], x[666], x[677], x[676], x[661], x[660], x[672], x[671], x[659]}), .y(y[226]));
  R1ind227 R1ind227_inst(.x({x[667], x[666], x[677], x[676], x[661], x[660], x[672], x[671], x[659]}), .y(y[227]));
  R1ind228 R1ind228_inst(.x({x[661], x[660], x[677], x[676], x[667], x[666], x[659]}), .y(y[228]));
  R1ind229 R1ind229_inst(.x({x[677], x[676], x[661], x[660], x[667], x[666], x[672], x[671], x[659]}), .y(y[229]));
  R1ind230 R1ind230_inst(.x({x[686], x[685], x[692], x[691], x[683], x[682], x[689], x[688], x[681]}), .y(y[230]));
  R1ind231 R1ind231_inst(.x({x[686], x[685], x[692], x[691], x[683], x[682], x[689], x[688], x[681]}), .y(y[231]));
  R1ind232 R1ind232_inst(.x({x[683], x[682], x[692], x[691], x[686], x[685], x[681]}), .y(y[232]));
  R1ind233 R1ind233_inst(.x({x[692], x[691], x[683], x[682], x[686], x[685], x[689], x[688], x[681]}), .y(y[233]));
  R1ind234 R1ind234_inst(.x({x[699], x[698], x[705], x[704], x[696], x[695], x[702], x[701], x[694]}), .y(y[234]));
  R1ind235 R1ind235_inst(.x({x[699], x[698], x[705], x[704], x[696], x[695], x[702], x[701], x[694]}), .y(y[235]));
  R1ind236 R1ind236_inst(.x({x[696], x[695], x[705], x[704], x[699], x[698], x[694]}), .y(y[236]));
  R1ind237 R1ind237_inst(.x({x[705], x[704], x[696], x[695], x[699], x[698], x[702], x[701], x[694]}), .y(y[237]));
  R1ind238 R1ind238_inst(.x({x[712], x[711], x[718], x[717], x[709], x[708], x[715], x[714], x[707]}), .y(y[238]));
  R1ind239 R1ind239_inst(.x({x[712], x[711], x[718], x[717], x[709], x[708], x[715], x[714], x[707]}), .y(y[239]));
  R1ind240 R1ind240_inst(.x({x[709], x[708], x[718], x[717], x[712], x[711], x[707]}), .y(y[240]));
  R1ind241 R1ind241_inst(.x({x[718], x[717], x[709], x[708], x[712], x[711], x[715], x[714], x[707]}), .y(y[241]));
  R1ind242 R1ind242_inst(.x({x[725], x[724], x[731], x[730], x[722], x[721], x[728], x[727], x[720]}), .y(y[242]));
  R1ind243 R1ind243_inst(.x({x[725], x[724], x[731], x[730], x[722], x[721], x[728], x[727], x[720]}), .y(y[243]));
  R1ind244 R1ind244_inst(.x({x[722], x[721], x[731], x[730], x[725], x[724], x[720]}), .y(y[244]));
  R1ind245 R1ind245_inst(.x({x[731], x[730], x[722], x[721], x[725], x[724], x[728], x[727], x[720]}), .y(y[245]));
  R1ind246 R1ind246_inst(.x({x[738], x[737], x[744], x[743], x[735], x[734], x[741], x[740], x[733]}), .y(y[246]));
  R1ind247 R1ind247_inst(.x({x[738], x[737], x[744], x[743], x[735], x[734], x[741], x[740], x[733]}), .y(y[247]));
  R1ind248 R1ind248_inst(.x({x[735], x[734], x[744], x[743], x[738], x[737], x[733]}), .y(y[248]));
  R1ind249 R1ind249_inst(.x({x[744], x[743], x[735], x[734], x[738], x[737], x[741], x[740], x[733]}), .y(y[249]));
  R1ind250 R1ind250_inst(.x({x[751], x[750], x[757], x[756], x[748], x[747], x[754], x[753], x[746]}), .y(y[250]));
  R1ind251 R1ind251_inst(.x({x[751], x[750], x[757], x[756], x[748], x[747], x[754], x[753], x[746]}), .y(y[251]));
  R1ind252 R1ind252_inst(.x({x[748], x[747], x[757], x[756], x[751], x[750], x[746]}), .y(y[252]));
  R1ind253 R1ind253_inst(.x({x[757], x[756], x[748], x[747], x[751], x[750], x[754], x[753], x[746]}), .y(y[253]));
  R1ind254 R1ind254_inst(.x({x[764], x[763], x[770], x[769], x[761], x[760], x[767], x[766], x[759]}), .y(y[254]));
  R1ind255 R1ind255_inst(.x({x[764], x[763], x[770], x[769], x[761], x[760], x[767], x[766], x[759]}), .y(y[255]));
  R1ind256 R1ind256_inst(.x({x[761], x[760], x[770], x[769], x[764], x[763], x[759]}), .y(y[256]));
  R1ind257 R1ind257_inst(.x({x[770], x[769], x[761], x[760], x[764], x[763], x[767], x[766], x[759]}), .y(y[257]));
  R1ind258 R1ind258_inst(.x({x[777], x[776], x[783], x[782], x[774], x[773], x[780], x[779], x[772]}), .y(y[258]));
  R1ind259 R1ind259_inst(.x({x[777], x[776], x[783], x[782], x[774], x[773], x[780], x[779], x[772]}), .y(y[259]));
  R1ind260 R1ind260_inst(.x({x[774], x[773], x[783], x[782], x[777], x[776], x[772]}), .y(y[260]));
  R1ind261 R1ind261_inst(.x({x[783], x[782], x[774], x[773], x[777], x[776], x[780], x[779], x[772]}), .y(y[261]));
  R1ind262 R1ind262_inst(.x({x[787], x[786], x[785], x[319], x[318], x[317], x[435]}), .y(y[262]));
  R1ind263 R1ind263_inst(.x({x[790], x[789], x[788], x[404], x[403], x[402], x[435]}), .y(y[263]));
  R1ind264 R1ind264_inst(.x({x[793], x[792], x[791], x[234], x[233], x[232], x[435]}), .y(y[264]));
  R1ind265 R1ind265_inst(.x({x[795], x[794], x[785], x[323], x[322], x[317], x[435]}), .y(y[265]));
  R1ind266 R1ind266_inst(.x({x[797], x[796], x[788], x[408], x[407], x[402], x[435]}), .y(y[266]));
  R1ind267 R1ind267_inst(.x({x[799], x[798], x[791], x[238], x[237], x[232], x[435]}), .y(y[267]));
  R1ind268 R1ind268_inst(.x({x[801], x[800], x[785], x[327], x[326], x[317], x[435]}), .y(y[268]));
  R1ind269 R1ind269_inst(.x({x[803], x[802], x[788], x[412], x[411], x[402], x[435]}), .y(y[269]));
  R1ind270 R1ind270_inst(.x({x[805], x[804], x[791], x[242], x[241], x[232], x[435]}), .y(y[270]));
  R1ind271 R1ind271_inst(.x({x[807], x[806], x[785], x[331], x[330], x[317], x[435]}), .y(y[271]));
  R1ind272 R1ind272_inst(.x({x[809], x[808], x[791], x[246], x[245], x[232], x[435]}), .y(y[272]));
  R1ind273 R1ind273_inst(.x({x[811], x[810], x[788], x[416], x[415], x[402], x[435]}), .y(y[273]));
  R1ind274 R1ind274_inst(.x({x[814], x[813], x[812], x[336], x[335], x[334], x[435]}), .y(y[274]));
  R1ind275 R1ind275_inst(.x({x[817], x[816], x[815], x[149], x[148], x[147], x[435]}), .y(y[275]));
  R1ind276 R1ind276_inst(.x({x[820], x[819], x[818], x[387], x[386], x[385], x[435]}), .y(y[276]));
  R1ind277 R1ind277_inst(.x({x[823], x[822], x[821], x[217], x[216], x[215], x[435]}), .y(y[277]));
  R1ind278 R1ind278_inst(.x({x[825], x[824], x[812], x[340], x[339], x[334], x[435]}), .y(y[278]));
  R1ind279 R1ind279_inst(.x({x[827], x[826], x[815], x[153], x[152], x[147], x[435]}), .y(y[279]));
  R1ind280 R1ind280_inst(.x({x[829], x[828], x[818], x[391], x[390], x[385], x[435]}), .y(y[280]));
  R1ind281 R1ind281_inst(.x({x[831], x[830], x[821], x[221], x[220], x[215], x[435]}), .y(y[281]));
  R1ind282 R1ind282_inst(.x({x[833], x[832], x[812], x[344], x[343], x[334], x[435]}), .y(y[282]));
  R1ind283 R1ind283_inst(.x({x[835], x[834], x[815], x[157], x[156], x[147], x[435]}), .y(y[283]));
  R1ind284 R1ind284_inst(.x({x[837], x[836], x[821], x[225], x[224], x[215], x[435]}), .y(y[284]));
  R1ind285 R1ind285_inst(.x({x[839], x[838], x[818], x[395], x[394], x[385], x[435]}), .y(y[285]));
  R1ind286 R1ind286_inst(.x({x[841], x[840], x[812], x[348], x[347], x[334], x[435]}), .y(y[286]));
  R1ind287 R1ind287_inst(.x({x[843], x[842], x[815], x[161], x[160], x[147], x[435]}), .y(y[287]));
  R1ind288 R1ind288_inst(.x({x[845], x[844], x[818], x[399], x[398], x[385], x[435]}), .y(y[288]));
  R1ind289 R1ind289_inst(.x({x[847], x[846], x[821], x[229], x[228], x[215], x[435]}), .y(y[289]));
  R1ind290 R1ind290_inst(.x({x[850], x[849], x[848], x[285], x[284], x[283], x[435]}), .y(y[290]));
  R1ind291 R1ind291_inst(.x({x[853], x[852], x[851], x[268], x[267], x[266], x[435]}), .y(y[291]));
  R1ind292 R1ind292_inst(.x({x[856], x[855], x[854], x[370], x[369], x[368], x[435]}), .y(y[292]));
  R1ind293 R1ind293_inst(.x({x[858], x[857], x[848], x[289], x[288], x[283], x[435]}), .y(y[293]));
  R1ind294 R1ind294_inst(.x({x[860], x[859], x[851], x[272], x[271], x[266], x[435]}), .y(y[294]));
  R1ind295 R1ind295_inst(.x({x[862], x[861], x[854], x[374], x[373], x[368], x[435]}), .y(y[295]));
  R1ind296 R1ind296_inst(.x({x[864], x[863], x[848], x[293], x[292], x[283], x[435]}), .y(y[296]));
  R1ind297 R1ind297_inst(.x({x[866], x[865], x[854], x[378], x[377], x[368], x[435]}), .y(y[297]));
  R1ind298 R1ind298_inst(.x({x[868], x[867], x[851], x[276], x[275], x[266], x[435]}), .y(y[298]));
  R1ind299 R1ind299_inst(.x({x[870], x[869], x[848], x[297], x[296], x[283], x[435]}), .y(y[299]));
  R1ind300 R1ind300_inst(.x({x[872], x[871], x[851], x[280], x[279], x[266], x[435]}), .y(y[300]));
  R1ind301 R1ind301_inst(.x({x[874], x[873], x[854], x[382], x[381], x[368], x[435]}), .y(y[301]));
  R1ind302 R1ind302_inst(.x({x[877], x[876], x[875], x[302], x[301], x[300], x[435]}), .y(y[302]));
  R1ind303 R1ind303_inst(.x({x[880], x[879], x[878], x[251], x[250], x[249], x[435]}), .y(y[303]));
  R1ind304 R1ind304_inst(.x({x[883], x[882], x[881], x[353], x[352], x[351], x[435]}), .y(y[304]));
  R1ind305 R1ind305_inst(.x({x[885], x[884], x[875], x[306], x[305], x[300], x[435]}), .y(y[305]));
  R1ind306 R1ind306_inst(.x({x[887], x[886], x[878], x[255], x[254], x[249], x[435]}), .y(y[306]));
  R1ind307 R1ind307_inst(.x({x[889], x[888], x[881], x[357], x[356], x[351], x[435]}), .y(y[307]));
  R1ind308 R1ind308_inst(.x({x[891], x[890], x[875], x[310], x[309], x[300], x[435]}), .y(y[308]));
  R1ind309 R1ind309_inst(.x({x[893], x[892], x[878], x[259], x[258], x[249], x[435]}), .y(y[309]));
  R1ind310 R1ind310_inst(.x({x[895], x[894], x[881], x[361], x[360], x[351], x[435]}), .y(y[310]));
  R1ind311 R1ind311_inst(.x({x[897], x[896], x[875], x[314], x[313], x[300], x[435]}), .y(y[311]));
  R1ind312 R1ind312_inst(.x({x[899], x[898], x[881], x[365], x[364], x[351], x[435]}), .y(y[312]));
  R1ind313 R1ind313_inst(.x({x[901], x[900], x[878], x[263], x[262], x[249], x[435]}), .y(y[313]));
  R1ind314 R1ind314_inst(.x({x[904], x[903], x[902], x[166], x[165], x[164], x[435]}), .y(y[314]));
  R1ind315 R1ind315_inst(.x({x[906], x[905], x[902], x[170], x[169], x[164], x[435]}), .y(y[315]));
  R1ind316 R1ind316_inst(.x({x[908], x[907], x[902], x[174], x[173], x[164], x[435]}), .y(y[316]));
  R1ind317 R1ind317_inst(.x({x[910], x[909], x[902], x[178], x[177], x[164], x[435]}), .y(y[317]));
  R1ind318 R1ind318_inst(.x({x[913], x[912], x[911], x[200], x[199], x[198], x[435]}), .y(y[318]));
  R1ind319 R1ind319_inst(.x({x[915], x[914], x[911], x[204], x[203], x[198], x[435]}), .y(y[319]));
  R1ind320 R1ind320_inst(.x({x[917], x[916], x[911], x[208], x[207], x[198], x[435]}), .y(y[320]));
  R1ind321 R1ind321_inst(.x({x[919], x[918], x[911], x[212], x[211], x[198], x[435]}), .y(y[321]));
  R1ind322 R1ind322_inst(.x({x[922], x[921], x[920], x[183], x[182], x[181], x[435]}), .y(y[322]));
  R1ind323 R1ind323_inst(.x({x[924], x[923], x[920], x[187], x[186], x[181], x[435]}), .y(y[323]));
  R1ind324 R1ind324_inst(.x({x[926], x[925], x[920], x[191], x[190], x[181], x[435]}), .y(y[324]));
  R1ind325 R1ind325_inst(.x({x[928], x[927], x[920], x[195], x[194], x[181], x[435]}), .y(y[325]));
  R1ind326 R1ind326_inst(.x({x[427], x[426], x[425], x[168], x[167], x[166], x[165], x[164]}), .y(y[326]));
  R1ind327 R1ind327_inst(.x({x[427], x[426], x[425], x[202], x[201], x[200], x[199], x[198]}), .y(y[327]));
  R1ind328 R1ind328_inst(.x({x[427], x[426], x[425], x[185], x[184], x[183], x[182], x[181]}), .y(y[328]));
  R1ind329 R1ind329_inst(.x({x[427], x[426], x[425], x[172], x[171], x[170], x[169], x[164]}), .y(y[329]));
  R1ind330 R1ind330_inst(.x({x[427], x[426], x[425], x[206], x[205], x[204], x[203], x[198]}), .y(y[330]));
  R1ind331 R1ind331_inst(.x({x[427], x[426], x[425], x[189], x[188], x[187], x[186], x[181]}), .y(y[331]));
  R1ind332 R1ind332_inst(.x({x[427], x[426], x[425], x[176], x[175], x[174], x[173], x[164]}), .y(y[332]));
  R1ind333 R1ind333_inst(.x({x[427], x[426], x[425], x[210], x[209], x[208], x[207], x[198]}), .y(y[333]));
  R1ind334 R1ind334_inst(.x({x[427], x[426], x[425], x[193], x[192], x[191], x[190], x[181]}), .y(y[334]));
  R1ind335 R1ind335_inst(.x({x[424], x[423], x[422], x[430], x[429], x[428], x[435], x[421], x[420], x[419], x[427], x[426], x[425], x[180], x[179], x[178], x[177], x[164]}), .y(y[335]));
  R1ind336 R1ind336_inst(.x({x[424], x[423], x[422], x[435], x[421], x[420], x[419], x[430], x[429], x[428], x[427], x[426], x[425], x[197], x[196], x[195], x[194], x[181]}), .y(y[336]));
  R1ind337 R1ind337_inst(.x({x[424], x[423], x[422], x[430], x[429], x[428], x[435], x[421], x[420], x[419], x[427], x[426], x[425], x[214], x[213], x[212], x[211], x[198]}), .y(y[337]));
  R1ind338 R1ind338_inst(.x({x[427], x[426], x[425], x[253], x[252], x[251], x[250], x[249]}), .y(y[338]));
  R1ind339 R1ind339_inst(.x({x[427], x[426], x[425], x[151], x[150], x[149], x[148], x[147]}), .y(y[339]));
  R1ind340 R1ind340_inst(.x({x[427], x[426], x[425], x[219], x[218], x[217], x[216], x[215]}), .y(y[340]));
  R1ind341 R1ind341_inst(.x({x[427], x[426], x[425], x[236], x[235], x[234], x[233], x[232]}), .y(y[341]));
  R1ind342 R1ind342_inst(.x({x[427], x[426], x[425], x[257], x[256], x[255], x[254], x[249]}), .y(y[342]));
  R1ind343 R1ind343_inst(.x({x[427], x[426], x[425], x[155], x[154], x[153], x[152], x[147]}), .y(y[343]));
  R1ind344 R1ind344_inst(.x({x[427], x[426], x[425], x[223], x[222], x[221], x[220], x[215]}), .y(y[344]));
  R1ind345 R1ind345_inst(.x({x[427], x[426], x[425], x[240], x[239], x[238], x[237], x[232]}), .y(y[345]));
  R1ind346 R1ind346_inst(.x({x[427], x[426], x[425], x[261], x[260], x[259], x[258], x[249]}), .y(y[346]));
  R1ind347 R1ind347_inst(.x({x[427], x[426], x[425], x[159], x[158], x[157], x[156], x[147]}), .y(y[347]));
  R1ind348 R1ind348_inst(.x({x[427], x[426], x[425], x[244], x[243], x[242], x[241], x[232]}), .y(y[348]));
  R1ind349 R1ind349_inst(.x({x[427], x[426], x[425], x[227], x[226], x[225], x[224], x[215]}), .y(y[349]));
  R1ind350 R1ind350_inst(.x({x[424], x[423], x[422], x[435], x[421], x[420], x[419], x[430], x[429], x[428], x[427], x[426], x[425], x[265], x[264], x[263], x[262], x[249]}), .y(y[350]));
  R1ind351 R1ind351_inst(.x({x[424], x[423], x[422], x[430], x[429], x[428], x[435], x[421], x[420], x[419], x[427], x[426], x[425], x[163], x[162], x[161], x[160], x[147]}), .y(y[351]));
  R1ind352 R1ind352_inst(.x({x[430], x[429], x[428], x[435], x[424], x[423], x[422], x[421], x[420], x[419], x[427], x[426], x[425], x[231], x[230], x[229], x[228], x[215]}), .y(y[352]));
  R1ind353 R1ind353_inst(.x({x[424], x[423], x[422], x[435], x[430], x[429], x[428], x[421], x[420], x[419], x[427], x[426], x[425], x[248], x[247], x[246], x[245], x[232]}), .y(y[353]));
  R1ind354 R1ind354_inst(.x({x[405], x[406], x[427], x[426], x[425], x[404], x[403], x[402]}), .y(y[354]));
  R1ind355 R1ind355_inst(.x({x[354], x[355], x[427], x[426], x[425], x[353], x[352], x[351]}), .y(y[355]));
  R1ind356 R1ind356_inst(.x({x[371], x[372], x[427], x[426], x[425], x[370], x[369], x[368]}), .y(y[356]));
  R1ind357 R1ind357_inst(.x({x[409], x[410], x[427], x[426], x[425], x[408], x[407], x[402]}), .y(y[357]));
  R1ind358 R1ind358_inst(.x({x[358], x[359], x[427], x[426], x[425], x[357], x[356], x[351]}), .y(y[358]));
  R1ind359 R1ind359_inst(.x({x[375], x[376], x[427], x[426], x[425], x[374], x[373], x[368]}), .y(y[359]));
  R1ind360 R1ind360_inst(.x({x[413], x[414], x[427], x[426], x[425], x[412], x[411], x[402]}), .y(y[360]));
  R1ind361 R1ind361_inst(.x({x[380], x[379], x[427], x[426], x[425], x[378], x[377], x[368]}), .y(y[361]));
  R1ind362 R1ind362_inst(.x({x[362], x[363], x[427], x[426], x[425], x[361], x[360], x[351]}), .y(y[362]));
  R1ind363 R1ind363_inst(.x({x[424], x[423], x[422], x[435], x[430], x[429], x[428], x[421], x[420], x[419], x[417], x[418], x[427], x[426], x[425], x[416], x[415], x[402]}), .y(y[363]));
  R1ind364 R1ind364_inst(.x({x[435], x[430], x[429], x[428], x[424], x[423], x[422], x[421], x[420], x[419], x[427], x[426], x[425], x[366], x[367], x[365], x[364], x[351]}), .y(y[364]));
  R1ind365 R1ind365_inst(.x({x[435], x[430], x[429], x[428], x[424], x[423], x[422], x[421], x[420], x[419], x[384], x[383], x[427], x[426], x[425], x[382], x[381], x[368]}), .y(y[365]));
  R1ind366 R1ind366_inst(.x({x[427], x[426], x[425], x[286], x[287], x[285], x[284], x[283]}), .y(y[366]));
  R1ind367 R1ind367_inst(.x({x[427], x[426], x[425], x[337], x[338], x[336], x[335], x[334]}), .y(y[367]));
  R1ind368 R1ind368_inst(.x({x[427], x[426], x[425], x[320], x[321], x[319], x[318], x[317]}), .y(y[368]));
  R1ind369 R1ind369_inst(.x({x[427], x[426], x[425], x[290], x[291], x[289], x[288], x[283]}), .y(y[369]));
  R1ind370 R1ind370_inst(.x({x[427], x[426], x[425], x[341], x[342], x[340], x[339], x[334]}), .y(y[370]));
  R1ind371 R1ind371_inst(.x({x[427], x[426], x[425], x[324], x[325], x[323], x[322], x[317]}), .y(y[371]));
  R1ind372 R1ind372_inst(.x({x[427], x[426], x[425], x[294], x[295], x[293], x[292], x[283]}), .y(y[372]));
  R1ind373 R1ind373_inst(.x({x[427], x[426], x[425], x[345], x[346], x[344], x[343], x[334]}), .y(y[373]));
  R1ind374 R1ind374_inst(.x({x[427], x[426], x[425], x[328], x[329], x[327], x[326], x[317]}), .y(y[374]));
  R1ind375 R1ind375_inst(.x({x[424], x[423], x[422], x[435], x[430], x[429], x[428], x[421], x[420], x[419], x[427], x[426], x[425], x[298], x[299], x[297], x[296], x[283]}), .y(y[375]));
  R1ind376 R1ind376_inst(.x({x[424], x[423], x[422], x[430], x[429], x[428], x[435], x[421], x[420], x[419], x[427], x[426], x[425], x[332], x[333], x[331], x[330], x[317]}), .y(y[376]));
  R1ind377 R1ind377_inst(.x({x[424], x[423], x[422], x[435], x[430], x[429], x[428], x[421], x[420], x[419], x[427], x[426], x[425], x[349], x[350], x[348], x[347], x[334]}), .y(y[377]));
  R1ind378 R1ind378_inst(.x({x[427], x[426], x[425], x[269], x[270], x[268], x[267], x[266]}), .y(y[378]));
  R1ind379 R1ind379_inst(.x({x[427], x[426], x[425], x[273], x[274], x[272], x[271], x[266]}), .y(y[379]));
  R1ind380 R1ind380_inst(.x({x[427], x[426], x[425], x[277], x[278], x[276], x[275], x[266]}), .y(y[380]));
  R1ind381 R1ind381_inst(.x({x[435], x[430], x[429], x[428], x[421], x[420], x[419], x[424], x[423], x[422], x[427], x[426], x[425], x[281], x[282], x[280], x[279], x[266]}), .y(y[381]));
  R1ind382 R1ind382_inst(.x({x[427], x[426], x[425], x[303], x[304], x[302], x[301], x[300]}), .y(y[382]));
  R1ind383 R1ind383_inst(.x({x[307], x[308], x[427], x[426], x[425], x[306], x[305], x[300]}), .y(y[383]));
  R1ind384 R1ind384_inst(.x({x[427], x[426], x[425], x[311], x[312], x[310], x[309], x[300]}), .y(y[384]));
  R1ind385 R1ind385_inst(.x({x[435], x[424], x[423], x[422], x[430], x[429], x[428], x[421], x[420], x[419], x[427], x[426], x[425], x[315], x[316], x[314], x[313], x[300]}), .y(y[385]));
  R1ind386 R1ind386_inst(.x({x[427], x[426], x[425], x[389], x[388], x[387], x[386], x[385]}), .y(y[386]));
  R1ind387 R1ind387_inst(.x({x[427], x[426], x[425], x[392], x[393], x[391], x[390], x[385]}), .y(y[387]));
  R1ind388 R1ind388_inst(.x({x[427], x[426], x[425], x[396], x[397], x[395], x[394], x[385]}), .y(y[388]));
  R1ind389 R1ind389_inst(.x({x[424], x[423], x[422], x[435], x[430], x[429], x[428], x[421], x[420], x[419], x[400], x[401], x[427], x[426], x[425], x[399], x[398], x[385]}), .y(y[389]));
endmodule

module R2ind0(x, y);
 input [5:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = t[1] ^ x[5];
  assign t[10] = (1'b0);
  assign t[11] = (x[0]);
  assign t[1] = (t[2] & ~t[3] & ~t[4] & ~t[5] & ~t[6]);
  assign t[2] = t[7] ^ x[5];
  assign t[3] = t[8] ^ x[1];
  assign t[4] = t[9] ^ x[2];
  assign t[5] = t[10] ^ x[3];
  assign t[6] = t[11] ^ x[4];
  assign t[7] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = (1'b0);
  assign t[9] = (1'b0);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind3(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (1'b0);
  assign y = t[0];
endmodule

module R2ind4(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind5(x, y);
 input [11:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[14] ^ x[11];
  assign t[11] = (~t[15] & t[16]);
  assign t[12] = (~t[17] & t[18]);
  assign t[13] = (~t[19] & t[20]);
  assign t[14] = (~t[21] & t[22]);
  assign t[15] = t[23] ^ x[1];
  assign t[16] = t[24] ^ x[2];
  assign t[17] = t[25] ^ x[4];
  assign t[18] = t[26] ^ x[5];
  assign t[19] = t[27] ^ x[7];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[28] ^ x[8];
  assign t[21] = t[29] ^ x[10];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[24] = (x[0]);
  assign t[25] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[26] = (x[3]);
  assign t[27] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[6]);
  assign t[29] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (x[9]);
  assign t[3] = (t[7]);
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind6(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind7(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind8(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind9(x, y);
 input [11:0] x;
 output y;

 wire [30:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[14] ^ x[11];
  assign t[11] = (~t[15] & t[16]);
  assign t[12] = (~t[17] & t[18]);
  assign t[13] = (~t[19] & t[20]);
  assign t[14] = (~t[21] & t[22]);
  assign t[15] = t[23] ^ x[1];
  assign t[16] = t[24] ^ x[2];
  assign t[17] = t[25] ^ x[4];
  assign t[18] = t[26] ^ x[5];
  assign t[19] = t[27] ^ x[7];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[28] ^ x[8];
  assign t[21] = t[29] ^ x[10];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = (x[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[0] & 1'b0 & ~1'b0 & ~1'b0) | (~x[0] & ~1'b0 & 1'b0 & ~1'b0) | (~x[0] & ~1'b0 & ~1'b0 & 1'b0) | (x[0] & 1'b0 & 1'b0 & ~1'b0) | (x[0] & 1'b0 & ~1'b0 & 1'b0) | (x[0] & ~1'b0 & 1'b0 & 1'b0) | (~x[0] & 1'b0 & 1'b0 & 1'b0);
  assign t[24] = (x[0]);
  assign t[25] = (x[3] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[3] & 1'b0 & ~1'b0 & ~1'b0) | (~x[3] & ~1'b0 & 1'b0 & ~1'b0) | (~x[3] & ~1'b0 & ~1'b0 & 1'b0) | (x[3] & 1'b0 & 1'b0 & ~1'b0) | (x[3] & 1'b0 & ~1'b0 & 1'b0) | (x[3] & ~1'b0 & 1'b0 & 1'b0) | (~x[3] & 1'b0 & 1'b0 & 1'b0);
  assign t[26] = (x[3]);
  assign t[27] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[6]);
  assign t[29] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (x[9]);
  assign t[3] = (t[7]);
  assign t[4] = (t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = t[11] ^ x[2];
  assign t[8] = t[12] ^ x[5];
  assign t[9] = t[13] ^ x[8];
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [12:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = ~(t[14] & t[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[3];
  assign t[16] = t[20] ^ x[6];
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[12];
  assign t[19] = (~t[23] & t[24]);
  assign t[1] = t[11] ^ t[2];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[3];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[6];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[3] & t[12]);
  assign t[30] = t[38] ^ x[12];
  assign t[31] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[1]);
  assign t[33] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[4]);
  assign t[35] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[7]);
  assign t[37] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[13]);
  assign t[5] = ~(t[6] & t[14]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(x[0]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind11(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind12(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind13(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind14(x, y);
 input [12:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = ~(t[14] & t[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[3];
  assign t[16] = t[20] ^ x[6];
  assign t[17] = t[21] ^ x[9];
  assign t[18] = t[22] ^ x[12];
  assign t[19] = (~t[23] & t[24]);
  assign t[1] = t[11] ^ t[2];
  assign t[20] = (~t[25] & t[26]);
  assign t[21] = (~t[27] & t[28]);
  assign t[22] = (~t[29] & t[30]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[3];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[6];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[9];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[3] & t[12]);
  assign t[30] = t[38] ^ x[12];
  assign t[31] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[1]);
  assign t[33] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[4]);
  assign t[35] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[36] = (x[7]);
  assign t[37] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[38] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[13]);
  assign t[5] = ~(t[6] & t[14]);
  assign t[6] = ~(t[7] & t[8]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(x[0]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [12:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[3];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[12];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = ~(t[10] ^ t[2]);
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[1]);
  assign t[32] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[4]);
  assign t[34] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[7]);
  assign t[36] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[10]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[5] & t[12]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[10] & t[13]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind16(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind17(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind18(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind19(x, y);
 input [12:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[3];
  assign t[15] = t[19] ^ x[6];
  assign t[16] = t[20] ^ x[9];
  assign t[17] = t[21] ^ x[12];
  assign t[18] = (~t[22] & t[23]);
  assign t[19] = (~t[24] & t[25]);
  assign t[1] = ~(t[10] ^ t[2]);
  assign t[20] = (~t[26] & t[27]);
  assign t[21] = (~t[28] & t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[3];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[6];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[9];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[12];
  assign t[2] = ~(t[3] | t[4]);
  assign t[30] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[1]);
  assign t[32] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[4]);
  assign t[34] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[7]);
  assign t[36] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[37] = (x[10]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[5] & t[12]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[10] & t[13]);
  assign t[9] = ~(t[12] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [12:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[3];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[9];
  assign t[15] = t[19] ^ x[12];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[8] ^ t[2];
  assign t[20] = t[28] ^ x[2];
  assign t[21] = t[29] ^ x[3];
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[6];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[9];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[29] = (x[1]);
  assign t[2] = ~(t[3] & t[9]);
  assign t[30] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[4]);
  assign t[32] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[7]);
  assign t[34] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[10]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[7] = ~(t[9] & t[8]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind21(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind22(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind23(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind24(x, y);
 input [12:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[3];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[9];
  assign t[15] = t[19] ^ x[12];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[22] & t[23]);
  assign t[18] = (~t[24] & t[25]);
  assign t[19] = (~t[26] & t[27]);
  assign t[1] = t[8] ^ t[2];
  assign t[20] = t[28] ^ x[2];
  assign t[21] = t[29] ^ x[3];
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[6];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[9];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[29] = (x[1]);
  assign t[2] = ~(t[3] & t[9]);
  assign t[30] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[31] = (x[4]);
  assign t[32] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[33] = (x[7]);
  assign t[34] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[35] = (x[10]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[7] = ~(t[9] & t[8]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [12:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[3];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[21] & t[22]);
  assign t[17] = (~t[23] & t[24]);
  assign t[18] = (~t[25] & t[26]);
  assign t[19] = t[27] ^ x[2];
  assign t[1] = ~(t[7] ^ t[2]);
  assign t[20] = t[28] ^ x[3];
  assign t[21] = t[29] ^ x[5];
  assign t[22] = t[30] ^ x[6];
  assign t[23] = t[31] ^ x[8];
  assign t[24] = t[32] ^ x[9];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[12];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[1]);
  assign t[29] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[31] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[7]);
  assign t[33] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[10]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[6] = ~(t[7] & t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~1'b0 & ~1'b0 & ~1'b0) | (~t[0] & 1'b0 & ~1'b0 & ~1'b0) | (~t[0] & ~1'b0 & 1'b0 & ~1'b0) | (~t[0] & ~1'b0 & ~1'b0 & 1'b0) | (t[0] & 1'b0 & 1'b0 & ~1'b0) | (t[0] & 1'b0 & ~1'b0 & 1'b0) | (t[0] & ~1'b0 & 1'b0 & 1'b0) | (~t[0] & 1'b0 & 1'b0 & 1'b0);
endmodule

module R2ind26(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind27(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind28(y);
 output y;

  assign y = (1'b0);
endmodule

module R2ind29(x, y);
 input [12:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = ~(x[0] | t[1]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[3];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[9];
  assign t[14] = t[18] ^ x[12];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[21] & t[22]);
  assign t[17] = (~t[23] & t[24]);
  assign t[18] = (~t[25] & t[26]);
  assign t[19] = t[27] ^ x[2];
  assign t[1] = ~(t[7] ^ t[2]);
  assign t[20] = t[28] ^ x[3];
  assign t[21] = t[29] ^ x[5];
  assign t[22] = t[30] ^ x[6];
  assign t[23] = t[31] ^ x[8];
  assign t[24] = t[32] ^ x[9];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[12];
  assign t[27] = (x[1] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[1] & 1'b0 & ~1'b0 & ~1'b0) | (~x[1] & ~1'b0 & 1'b0 & ~1'b0) | (~x[1] & ~1'b0 & ~1'b0 & 1'b0) | (x[1] & 1'b0 & 1'b0 & ~1'b0) | (x[1] & 1'b0 & ~1'b0 & 1'b0) | (x[1] & ~1'b0 & 1'b0 & 1'b0) | (~x[1] & 1'b0 & 1'b0 & 1'b0);
  assign t[28] = (x[1]);
  assign t[29] = (x[4] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[4] & 1'b0 & ~1'b0 & ~1'b0) | (~x[4] & ~1'b0 & 1'b0 & ~1'b0) | (~x[4] & ~1'b0 & ~1'b0 & 1'b0) | (x[4] & 1'b0 & 1'b0 & ~1'b0) | (x[4] & 1'b0 & ~1'b0 & 1'b0) | (x[4] & ~1'b0 & 1'b0 & 1'b0) | (~x[4] & 1'b0 & 1'b0 & 1'b0);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (x[4]);
  assign t[31] = (x[7] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[7] & 1'b0 & ~1'b0 & ~1'b0) | (~x[7] & ~1'b0 & 1'b0 & ~1'b0) | (~x[7] & ~1'b0 & ~1'b0 & 1'b0) | (x[7] & 1'b0 & 1'b0 & ~1'b0) | (x[7] & 1'b0 & ~1'b0 & 1'b0) | (x[7] & ~1'b0 & 1'b0 & 1'b0) | (~x[7] & 1'b0 & 1'b0 & 1'b0);
  assign t[32] = (x[7]);
  assign t[33] = (x[10] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[10] & 1'b0 & ~1'b0 & ~1'b0) | (~x[10] & ~1'b0 & 1'b0 & ~1'b0) | (~x[10] & ~1'b0 & ~1'b0 & 1'b0) | (x[10] & 1'b0 & 1'b0 & ~1'b0) | (x[10] & 1'b0 & ~1'b0 & 1'b0) | (x[10] & ~1'b0 & 1'b0 & 1'b0) | (~x[10] & 1'b0 & 1'b0 & 1'b0);
  assign t[34] = (x[10]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[4] = ~(x[0]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[6] = ~(t[7] & t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind31(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind32(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind33(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind34(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind36(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind37(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind38(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind39(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind41(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind46(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind51(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind56(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind61(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind66(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind71(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind76(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind81(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind86(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind91(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind96(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind101(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [16:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = t[1] ^ t[8];
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[8];
  assign t[14] = t[18] ^ x[11];
  assign t[15] = t[19] ^ x[14];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = x[6] ^ x[7];
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[8];
  assign t[23] = t[28] ^ x[11];
  assign t[24] = t[29] ^ x[14];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[0]);
  assign t[27] = (x[1]);
  assign t[28] = (x[2]);
  assign t[29] = (x[3]);
  assign t[2] = t[3] ^ t[9];
  assign t[3] = x[9] ^ x[10];
  assign t[4] = t[5] ^ t[10];
  assign t[5] = x[12] ^ x[13];
  assign t[6] = t[7] ^ t[11];
  assign t[7] = x[15] ^ x[16];
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0] & ~t[2] & ~t[4] & ~t[6]) | (~t[0] & t[2] & ~t[4] & ~t[6]) | (~t[0] & ~t[2] & t[4] & ~t[6]) | (~t[0] & ~t[2] & ~t[4] & t[6]) | (t[0] & t[2] & t[4] & ~t[6]) | (t[0] & t[2] & ~t[4] & t[6]) | (t[0] & ~t[2] & t[4] & t[6]) | (~t[0] & t[2] & t[4] & t[6]);
endmodule

module R2ind106(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[3]);
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[2]);
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[1]);
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [7:0] x;
 output y;

 wire [8:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[1] = x[6] ^ x[7];
  assign t[2] = (t[3]);
  assign t[3] = t[4] ^ x[5];
  assign t[4] = (~t[5] & t[6]);
  assign t[5] = t[7] ^ x[4];
  assign t[6] = t[8] ^ x[5];
  assign t[7] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [88:0] x;
 output y;

 wire [269:0] t;
  assign t[0] = t[1] ? t[2] : t[88];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[5];
  assign t[121] = t[153] ^ x[14];
  assign t[122] = t[154] ^ x[22];
  assign t[123] = t[155] ^ x[28];
  assign t[124] = t[156] ^ x[34];
  assign t[125] = t[157] ^ x[37];
  assign t[126] = t[158] ^ x[40];
  assign t[127] = t[159] ^ x[43];
  assign t[128] = t[160] ^ x[46];
  assign t[129] = t[161] ^ x[52];
  assign t[12] = ~(t[90] ^ t[17]);
  assign t[130] = t[162] ^ x[58];
  assign t[131] = t[163] ^ x[59];
  assign t[132] = t[164] ^ x[61];
  assign t[133] = t[165] ^ x[64];
  assign t[134] = t[166] ^ x[65];
  assign t[135] = t[167] ^ x[66];
  assign t[136] = t[168] ^ x[67];
  assign t[137] = t[169] ^ x[68];
  assign t[138] = t[170] ^ x[69];
  assign t[139] = t[171] ^ x[71];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[74];
  assign t[141] = t[173] ^ x[75];
  assign t[142] = t[174] ^ x[76];
  assign t[143] = t[175] ^ x[77];
  assign t[144] = t[176] ^ x[78];
  assign t[145] = t[177] ^ x[79];
  assign t[146] = t[178] ^ x[81];
  assign t[147] = t[179] ^ x[84];
  assign t[148] = t[180] ^ x[85];
  assign t[149] = t[181] ^ x[86];
  assign t[14] = ~(t[91] ^ t[92]);
  assign t[150] = t[182] ^ x[87];
  assign t[151] = t[183] ^ x[88];
  assign t[152] = (~t[184] & t[185]);
  assign t[153] = (~t[186] & t[187]);
  assign t[154] = (~t[188] & t[189]);
  assign t[155] = (~t[190] & t[191]);
  assign t[156] = (~t[192] & t[193]);
  assign t[157] = (~t[194] & t[195]);
  assign t[158] = (~t[196] & t[197]);
  assign t[159] = (~t[198] & t[199]);
  assign t[15] = ~(t[93] & t[94]);
  assign t[160] = (~t[200] & t[201]);
  assign t[161] = (~t[202] & t[203]);
  assign t[162] = (~t[204] & t[205]);
  assign t[163] = (~t[184] & t[206]);
  assign t[164] = (~t[186] & t[207]);
  assign t[165] = (~t[188] & t[208]);
  assign t[166] = (~t[192] & t[209]);
  assign t[167] = (~t[190] & t[210]);
  assign t[168] = (~t[204] & t[211]);
  assign t[169] = (~t[202] & t[212]);
  assign t[16] = ~(t[95] & t[96]);
  assign t[170] = (~t[184] & t[213]);
  assign t[171] = (~t[186] & t[214]);
  assign t[172] = (~t[188] & t[215]);
  assign t[173] = (~t[190] & t[216]);
  assign t[174] = (~t[192] & t[217]);
  assign t[175] = (~t[202] & t[218]);
  assign t[176] = (~t[204] & t[219]);
  assign t[177] = (~t[184] & t[220]);
  assign t[178] = (~t[186] & t[221]);
  assign t[179] = (~t[188] & t[222]);
  assign t[17] = ~(t[97] ^ t[98]);
  assign t[180] = (~t[190] & t[223]);
  assign t[181] = (~t[192] & t[224]);
  assign t[182] = (~t[202] & t[225]);
  assign t[183] = (~t[204] & t[226]);
  assign t[184] = t[227] ^ x[4];
  assign t[185] = t[228] ^ x[5];
  assign t[186] = t[229] ^ x[13];
  assign t[187] = t[230] ^ x[14];
  assign t[188] = t[231] ^ x[21];
  assign t[189] = t[232] ^ x[22];
  assign t[18] = t[95] ? x[15] : x[16];
  assign t[190] = t[233] ^ x[27];
  assign t[191] = t[234] ^ x[28];
  assign t[192] = t[235] ^ x[33];
  assign t[193] = t[236] ^ x[34];
  assign t[194] = t[237] ^ x[36];
  assign t[195] = t[238] ^ x[37];
  assign t[196] = t[239] ^ x[39];
  assign t[197] = t[240] ^ x[40];
  assign t[198] = t[241] ^ x[42];
  assign t[199] = t[242] ^ x[43];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[45];
  assign t[201] = t[244] ^ x[46];
  assign t[202] = t[245] ^ x[51];
  assign t[203] = t[246] ^ x[52];
  assign t[204] = t[247] ^ x[57];
  assign t[205] = t[248] ^ x[58];
  assign t[206] = t[249] ^ x[59];
  assign t[207] = t[250] ^ x[61];
  assign t[208] = t[251] ^ x[64];
  assign t[209] = t[252] ^ x[65];
  assign t[20] = ~(t[22] | t[23]);
  assign t[210] = t[253] ^ x[66];
  assign t[211] = t[254] ^ x[67];
  assign t[212] = t[255] ^ x[68];
  assign t[213] = t[256] ^ x[69];
  assign t[214] = t[257] ^ x[71];
  assign t[215] = t[258] ^ x[74];
  assign t[216] = t[259] ^ x[75];
  assign t[217] = t[260] ^ x[76];
  assign t[218] = t[261] ^ x[77];
  assign t[219] = t[262] ^ x[78];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[79];
  assign t[221] = t[264] ^ x[81];
  assign t[222] = t[265] ^ x[84];
  assign t[223] = t[266] ^ x[85];
  assign t[224] = t[267] ^ x[86];
  assign t[225] = t[268] ^ x[87];
  assign t[226] = t[269] ^ x[88];
  assign t[227] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[228] = (x[0]);
  assign t[229] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[230] = (x[9]);
  assign t[231] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[232] = (x[17]);
  assign t[233] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[234] = (x[23]);
  assign t[235] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[236] = (x[29]);
  assign t[237] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[238] = (x[35]);
  assign t[239] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[23] = ~(t[28] & t[29]);
  assign t[240] = (x[38]);
  assign t[241] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[242] = (x[41]);
  assign t[243] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[244] = (x[44]);
  assign t[245] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[246] = (x[47]);
  assign t[247] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[248] = (x[53]);
  assign t[249] = (x[1]);
  assign t[24] = ~(t[26] | t[30]);
  assign t[250] = (x[10]);
  assign t[251] = (x[18]);
  assign t[252] = (x[30]);
  assign t[253] = (x[24]);
  assign t[254] = (x[54]);
  assign t[255] = (x[48]);
  assign t[256] = (x[2]);
  assign t[257] = (x[11]);
  assign t[258] = (x[19]);
  assign t[259] = (x[25]);
  assign t[25] = ~(t[26] | t[31]);
  assign t[260] = (x[31]);
  assign t[261] = (x[49]);
  assign t[262] = (x[55]);
  assign t[263] = (x[3]);
  assign t[264] = (x[12]);
  assign t[265] = (x[20]);
  assign t[266] = (x[26]);
  assign t[267] = (x[32]);
  assign t[268] = (x[50]);
  assign t[269] = (x[56]);
  assign t[26] = ~(t[32]);
  assign t[27] = t[93] ? t[34] : t[33];
  assign t[28] = ~(t[35] | t[36]);
  assign t[29] = ~(t[37] & t[38]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[93] ? t[40] : t[39];
  assign t[31] = t[93] ? t[42] : t[41];
  assign t[32] = ~(t[95]);
  assign t[33] = ~(t[43] & t[96]);
  assign t[34] = ~(t[44] & t[45]);
  assign t[35] = ~(t[26] | t[46]);
  assign t[36] = ~(t[26] | t[47]);
  assign t[37] = t[96] & t[48];
  assign t[38] = t[44] | t[43];
  assign t[39] = ~(t[49] & t[45]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(x[7] & t[50]);
  assign t[41] = ~(t[44] & t[96]);
  assign t[42] = ~(t[43] & t[45]);
  assign t[43] = x[7] & t[94];
  assign t[44] = ~(x[7] | t[94]);
  assign t[45] = ~(t[96]);
  assign t[46] = t[93] ? t[33] : t[34];
  assign t[47] = t[93] ? t[52] : t[51];
  assign t[48] = ~(t[32] | t[93]);
  assign t[49] = ~(x[7] | t[53]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[94] | t[45]);
  assign t[51] = ~(t[96] & t[49]);
  assign t[52] = ~(x[7] & t[54]);
  assign t[53] = ~(t[94]);
  assign t[54] = ~(t[94] | t[96]);
  assign t[55] = t[6] ? t[56] : t[99];
  assign t[56] = x[6] ? t[58] : t[57];
  assign t[57] = x[7] ? t[60] : t[59];
  assign t[58] = t[61] ^ x[60];
  assign t[59] = t[62] ^ t[63];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[100] ^ t[64]);
  assign t[61] = x[62] ^ x[63];
  assign t[62] = t[95] ? x[62] : x[63];
  assign t[63] = ~(t[101] ^ t[65]);
  assign t[64] = ~(t[102] ^ t[103]);
  assign t[65] = ~(t[104] ^ t[105]);
  assign t[66] = t[1] ? t[67] : t[106];
  assign t[67] = x[6] ? t[69] : t[68];
  assign t[68] = x[7] ? t[71] : t[70];
  assign t[69] = t[72] ^ x[70];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[73] ^ t[74];
  assign t[71] = ~(t[107] ^ t[75]);
  assign t[72] = x[72] ^ x[73];
  assign t[73] = t[95] ? x[72] : x[73];
  assign t[74] = ~(t[108] ^ t[76]);
  assign t[75] = ~(t[109] ^ t[110]);
  assign t[76] = ~(t[111] ^ t[112]);
  assign t[77] = t[6] ? t[78] : t[113];
  assign t[78] = x[6] ? t[80] : t[79];
  assign t[79] = x[7] ? t[82] : t[81];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[83] ^ x[80];
  assign t[81] = t[84] ^ t[85];
  assign t[82] = ~(t[114] ^ t[86]);
  assign t[83] = x[82] ^ x[83];
  assign t[84] = t[95] ? x[82] : x[83];
  assign t[85] = ~(t[115] ^ t[87]);
  assign t[86] = ~(t[116] ^ t[117]);
  assign t[87] = ~(t[118] ^ t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[89] ^ t[14]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[55] & ~t[66] & ~t[77]) | (~t[0] & t[55] & ~t[66] & ~t[77]) | (~t[0] & ~t[55] & t[66] & ~t[77]) | (~t[0] & ~t[55] & ~t[66] & t[77]) | (t[0] & t[55] & t[66] & ~t[77]) | (t[0] & t[55] & ~t[66] & t[77]) | (t[0] & ~t[55] & t[66] & t[77]) | (~t[0] & t[55] & t[66] & t[77]);
endmodule

module R2ind111(x, y);
 input [58:0] x;
 output y;

 wire [92:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[21] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[19] ? x[27] : x[28];
  assign t[13] = ~(t[22] ^ t[15]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] ^ t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[11];
  assign t[29] = t[40] ^ x[14];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[17];
  assign t[31] = t[42] ^ x[20];
  assign t[32] = t[43] ^ x[26];
  assign t[33] = t[44] ^ x[34];
  assign t[34] = t[45] ^ x[40];
  assign t[35] = t[46] ^ x[46];
  assign t[36] = t[47] ^ x[52];
  assign t[37] = t[48] ^ x[58];
  assign t[38] = (~t[49] & t[50]);
  assign t[39] = (~t[51] & t[52]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[53] & t[54]);
  assign t[41] = (~t[55] & t[56]);
  assign t[42] = (~t[57] & t[58]);
  assign t[43] = (~t[59] & t[60]);
  assign t[44] = (~t[61] & t[62]);
  assign t[45] = (~t[63] & t[64]);
  assign t[46] = (~t[65] & t[66]);
  assign t[47] = (~t[67] & t[68]);
  assign t[48] = (~t[69] & t[70]);
  assign t[49] = t[71] ^ x[4];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[5];
  assign t[51] = t[73] ^ x[10];
  assign t[52] = t[74] ^ x[11];
  assign t[53] = t[75] ^ x[13];
  assign t[54] = t[76] ^ x[14];
  assign t[55] = t[77] ^ x[16];
  assign t[56] = t[78] ^ x[17];
  assign t[57] = t[79] ^ x[19];
  assign t[58] = t[80] ^ x[20];
  assign t[59] = t[81] ^ x[25];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[26];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[39];
  assign t[64] = t[86] ^ x[40];
  assign t[65] = t[87] ^ x[45];
  assign t[66] = t[88] ^ x[46];
  assign t[67] = t[89] ^ x[51];
  assign t[68] = t[90] ^ x[52];
  assign t[69] = t[91] ^ x[57];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[58];
  assign t[71] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[72] = (x[3]);
  assign t[73] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[9]);
  assign t[75] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[12]);
  assign t[77] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[15]);
  assign t[79] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[17] & t[18]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[86] = (x[38]);
  assign t[87] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[88] = (x[44]);
  assign t[89] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[8] = ~(t[19] & t[20]);
  assign t[90] = (x[50]);
  assign t[91] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[92] = (x[56]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [58:0] x;
 output y;

 wire [94:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[20] ? x[15] : x[16];
  assign t[13] = ~(t[21] ^ t[17]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[20] & t[26]);
  assign t[17] = ~(t[27] ^ t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = t[40] ^ x[5];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[41] ^ x[14];
  assign t[31] = t[42] ^ x[19];
  assign t[32] = t[43] ^ x[25];
  assign t[33] = t[44] ^ x[31];
  assign t[34] = t[45] ^ x[37];
  assign t[35] = t[46] ^ x[40];
  assign t[36] = t[47] ^ x[43];
  assign t[37] = t[48] ^ x[46];
  assign t[38] = t[49] ^ x[52];
  assign t[39] = t[50] ^ x[58];
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[51] & t[52]);
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = t[73] ^ x[4];
  assign t[52] = t[74] ^ x[5];
  assign t[53] = t[75] ^ x[13];
  assign t[54] = t[76] ^ x[14];
  assign t[55] = t[77] ^ x[18];
  assign t[56] = t[78] ^ x[19];
  assign t[57] = t[79] ^ x[24];
  assign t[58] = t[80] ^ x[25];
  assign t[59] = t[81] ^ x[30];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[31];
  assign t[61] = t[83] ^ x[36];
  assign t[62] = t[84] ^ x[37];
  assign t[63] = t[85] ^ x[39];
  assign t[64] = t[86] ^ x[40];
  assign t[65] = t[87] ^ x[42];
  assign t[66] = t[88] ^ x[43];
  assign t[67] = t[89] ^ x[45];
  assign t[68] = t[90] ^ x[46];
  assign t[69] = t[91] ^ x[51];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[52];
  assign t[71] = t[93] ^ x[57];
  assign t[72] = t[94] ^ x[58];
  assign t[73] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[74] = (x[2]);
  assign t[75] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[76] = (x[11]);
  assign t[77] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[17]);
  assign t[79] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[22]);
  assign t[81] = (x[26] & ~x[27] & ~x[28] & ~x[29]) | (~x[26] & x[27] & ~x[28] & ~x[29]) | (~x[26] & ~x[27] & x[28] & ~x[29]) | (~x[26] & ~x[27] & ~x[28] & x[29]) | (x[26] & x[27] & x[28] & ~x[29]) | (x[26] & x[27] & ~x[28] & x[29]) | (x[26] & ~x[27] & x[28] & x[29]) | (~x[26] & x[27] & x[28] & x[29]);
  assign t[82] = (x[28]);
  assign t[83] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[84] = (x[34]);
  assign t[85] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[38]);
  assign t[87] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[41]);
  assign t[89] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[19] ^ t[14]);
  assign t[90] = (x[44]);
  assign t[91] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[92] = (x[49]);
  assign t[93] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[94] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [58:0] x;
 output y;

 wire [92:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[21] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[19] ? x[27] : x[28];
  assign t[13] = ~(t[22] ^ t[15]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] ^ t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[11];
  assign t[29] = t[40] ^ x[14];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[17];
  assign t[31] = t[42] ^ x[20];
  assign t[32] = t[43] ^ x[26];
  assign t[33] = t[44] ^ x[34];
  assign t[34] = t[45] ^ x[40];
  assign t[35] = t[46] ^ x[46];
  assign t[36] = t[47] ^ x[52];
  assign t[37] = t[48] ^ x[58];
  assign t[38] = (~t[49] & t[50]);
  assign t[39] = (~t[51] & t[52]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[53] & t[54]);
  assign t[41] = (~t[55] & t[56]);
  assign t[42] = (~t[57] & t[58]);
  assign t[43] = (~t[59] & t[60]);
  assign t[44] = (~t[61] & t[62]);
  assign t[45] = (~t[63] & t[64]);
  assign t[46] = (~t[65] & t[66]);
  assign t[47] = (~t[67] & t[68]);
  assign t[48] = (~t[69] & t[70]);
  assign t[49] = t[71] ^ x[4];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[5];
  assign t[51] = t[73] ^ x[10];
  assign t[52] = t[74] ^ x[11];
  assign t[53] = t[75] ^ x[13];
  assign t[54] = t[76] ^ x[14];
  assign t[55] = t[77] ^ x[16];
  assign t[56] = t[78] ^ x[17];
  assign t[57] = t[79] ^ x[19];
  assign t[58] = t[80] ^ x[20];
  assign t[59] = t[81] ^ x[25];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[26];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[39];
  assign t[64] = t[86] ^ x[40];
  assign t[65] = t[87] ^ x[45];
  assign t[66] = t[88] ^ x[46];
  assign t[67] = t[89] ^ x[51];
  assign t[68] = t[90] ^ x[52];
  assign t[69] = t[91] ^ x[57];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[58];
  assign t[71] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[72] = (x[1]);
  assign t[73] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[9]);
  assign t[75] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[12]);
  assign t[77] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[15]);
  assign t[79] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[17] & t[18]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[82] = (x[22]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[86] = (x[36]);
  assign t[87] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[88] = (x[42]);
  assign t[89] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[8] = ~(t[19] & t[20]);
  assign t[90] = (x[48]);
  assign t[91] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[92] = (x[54]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [58:0] x;
 output y;

 wire [131:0] t;
  assign t[0] = t[1] ? t[2] : t[55];
  assign t[100] = t[122] ^ x[39];
  assign t[101] = t[123] ^ x[40];
  assign t[102] = t[124] ^ x[42];
  assign t[103] = t[125] ^ x[43];
  assign t[104] = t[126] ^ x[45];
  assign t[105] = t[127] ^ x[46];
  assign t[106] = t[128] ^ x[51];
  assign t[107] = t[129] ^ x[52];
  assign t[108] = t[130] ^ x[57];
  assign t[109] = t[131] ^ x[58];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[111] = (x[0]);
  assign t[112] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[113] = (x[9]);
  assign t[114] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[115] = (x[17]);
  assign t[116] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[117] = (x[23]);
  assign t[118] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[119] = (x[29]);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[121] = (x[35]);
  assign t[122] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[38]);
  assign t[124] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[41]);
  assign t[126] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[44]);
  assign t[128] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[129] = (x[47]);
  assign t[12] = ~(t[57] ^ t[17]);
  assign t[130] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[131] = (x[53]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[58] ^ t[59]);
  assign t[15] = ~(t[60] & t[61]);
  assign t[16] = ~(t[62] & t[63]);
  assign t[17] = ~(t[64] ^ t[65]);
  assign t[18] = t[62] ? x[15] : x[16];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[22] | t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[28] & t[29]);
  assign t[24] = ~(t[26] | t[30]);
  assign t[25] = ~(t[26] | t[31]);
  assign t[26] = ~(t[32]);
  assign t[27] = t[60] ? t[34] : t[33];
  assign t[28] = ~(t[35] | t[36]);
  assign t[29] = ~(t[37] & t[38]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[60] ? t[40] : t[39];
  assign t[31] = t[60] ? t[42] : t[41];
  assign t[32] = ~(t[62]);
  assign t[33] = ~(t[43] & t[63]);
  assign t[34] = ~(t[44] & t[45]);
  assign t[35] = ~(t[26] | t[46]);
  assign t[36] = ~(t[26] | t[47]);
  assign t[37] = t[63] & t[48];
  assign t[38] = t[44] | t[43];
  assign t[39] = ~(t[49] & t[45]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(x[7] & t[50]);
  assign t[41] = ~(t[44] & t[63]);
  assign t[42] = ~(t[43] & t[45]);
  assign t[43] = x[7] & t[61];
  assign t[44] = ~(x[7] | t[61]);
  assign t[45] = ~(t[63]);
  assign t[46] = t[60] ? t[33] : t[34];
  assign t[47] = t[60] ? t[52] : t[51];
  assign t[48] = ~(t[32] | t[60]);
  assign t[49] = ~(x[7] | t[53]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[61] | t[45]);
  assign t[51] = ~(t[63] & t[49]);
  assign t[52] = ~(x[7] & t[54]);
  assign t[53] = ~(t[61]);
  assign t[54] = ~(t[61] | t[63]);
  assign t[55] = (t[66]);
  assign t[56] = (t[67]);
  assign t[57] = (t[68]);
  assign t[58] = (t[69]);
  assign t[59] = (t[70]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = (t[73]);
  assign t[63] = (t[74]);
  assign t[64] = (t[75]);
  assign t[65] = (t[76]);
  assign t[66] = t[77] ^ x[5];
  assign t[67] = t[78] ^ x[14];
  assign t[68] = t[79] ^ x[22];
  assign t[69] = t[80] ^ x[28];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[81] ^ x[34];
  assign t[71] = t[82] ^ x[37];
  assign t[72] = t[83] ^ x[40];
  assign t[73] = t[84] ^ x[43];
  assign t[74] = t[85] ^ x[46];
  assign t[75] = t[86] ^ x[52];
  assign t[76] = t[87] ^ x[58];
  assign t[77] = (~t[88] & t[89]);
  assign t[78] = (~t[90] & t[91]);
  assign t[79] = (~t[92] & t[93]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[94] & t[95]);
  assign t[81] = (~t[96] & t[97]);
  assign t[82] = (~t[98] & t[99]);
  assign t[83] = (~t[100] & t[101]);
  assign t[84] = (~t[102] & t[103]);
  assign t[85] = (~t[104] & t[105]);
  assign t[86] = (~t[106] & t[107]);
  assign t[87] = (~t[108] & t[109]);
  assign t[88] = t[110] ^ x[4];
  assign t[89] = t[111] ^ x[5];
  assign t[8] = ~(t[56] ^ t[14]);
  assign t[90] = t[112] ^ x[13];
  assign t[91] = t[113] ^ x[14];
  assign t[92] = t[114] ^ x[21];
  assign t[93] = t[115] ^ x[22];
  assign t[94] = t[116] ^ x[27];
  assign t[95] = t[117] ^ x[28];
  assign t[96] = t[118] ^ x[33];
  assign t[97] = t[119] ^ x[34];
  assign t[98] = t[120] ^ x[36];
  assign t[99] = t[121] ^ x[37];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [88:0] x;
 output y;

 wire [277:0] t;
  assign t[0] = t[1] ? t[2] : t[96];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = (t[158]);
  assign t[127] = (t[159]);
  assign t[128] = t[160] ^ x[5];
  assign t[129] = t[161] ^ x[14];
  assign t[12] = ~(t[98] ^ t[17]);
  assign t[130] = t[162] ^ x[22];
  assign t[131] = t[163] ^ x[28];
  assign t[132] = t[164] ^ x[34];
  assign t[133] = t[165] ^ x[37];
  assign t[134] = t[166] ^ x[40];
  assign t[135] = t[167] ^ x[43];
  assign t[136] = t[168] ^ x[46];
  assign t[137] = t[169] ^ x[52];
  assign t[138] = t[170] ^ x[58];
  assign t[139] = t[171] ^ x[59];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[61];
  assign t[141] = t[173] ^ x[64];
  assign t[142] = t[174] ^ x[65];
  assign t[143] = t[175] ^ x[66];
  assign t[144] = t[176] ^ x[67];
  assign t[145] = t[177] ^ x[68];
  assign t[146] = t[178] ^ x[69];
  assign t[147] = t[179] ^ x[71];
  assign t[148] = t[180] ^ x[74];
  assign t[149] = t[181] ^ x[75];
  assign t[14] = ~(t[99] ^ t[100]);
  assign t[150] = t[182] ^ x[76];
  assign t[151] = t[183] ^ x[77];
  assign t[152] = t[184] ^ x[78];
  assign t[153] = t[185] ^ x[79];
  assign t[154] = t[186] ^ x[81];
  assign t[155] = t[187] ^ x[84];
  assign t[156] = t[188] ^ x[85];
  assign t[157] = t[189] ^ x[86];
  assign t[158] = t[190] ^ x[87];
  assign t[159] = t[191] ^ x[88];
  assign t[15] = ~(t[101] & t[102]);
  assign t[160] = (~t[192] & t[193]);
  assign t[161] = (~t[194] & t[195]);
  assign t[162] = (~t[196] & t[197]);
  assign t[163] = (~t[198] & t[199]);
  assign t[164] = (~t[200] & t[201]);
  assign t[165] = (~t[202] & t[203]);
  assign t[166] = (~t[204] & t[205]);
  assign t[167] = (~t[206] & t[207]);
  assign t[168] = (~t[208] & t[209]);
  assign t[169] = (~t[210] & t[211]);
  assign t[16] = ~(t[103] & t[104]);
  assign t[170] = (~t[212] & t[213]);
  assign t[171] = (~t[192] & t[214]);
  assign t[172] = (~t[194] & t[215]);
  assign t[173] = (~t[196] & t[216]);
  assign t[174] = (~t[200] & t[217]);
  assign t[175] = (~t[198] & t[218]);
  assign t[176] = (~t[212] & t[219]);
  assign t[177] = (~t[210] & t[220]);
  assign t[178] = (~t[192] & t[221]);
  assign t[179] = (~t[194] & t[222]);
  assign t[17] = ~(t[105] ^ t[106]);
  assign t[180] = (~t[196] & t[223]);
  assign t[181] = (~t[200] & t[224]);
  assign t[182] = (~t[198] & t[225]);
  assign t[183] = (~t[210] & t[226]);
  assign t[184] = (~t[212] & t[227]);
  assign t[185] = (~t[192] & t[228]);
  assign t[186] = (~t[194] & t[229]);
  assign t[187] = (~t[196] & t[230]);
  assign t[188] = (~t[200] & t[231]);
  assign t[189] = (~t[198] & t[232]);
  assign t[18] = t[103] ? x[15] : x[16];
  assign t[190] = (~t[210] & t[233]);
  assign t[191] = (~t[212] & t[234]);
  assign t[192] = t[235] ^ x[4];
  assign t[193] = t[236] ^ x[5];
  assign t[194] = t[237] ^ x[13];
  assign t[195] = t[238] ^ x[14];
  assign t[196] = t[239] ^ x[21];
  assign t[197] = t[240] ^ x[22];
  assign t[198] = t[241] ^ x[27];
  assign t[199] = t[242] ^ x[28];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[33];
  assign t[201] = t[244] ^ x[34];
  assign t[202] = t[245] ^ x[36];
  assign t[203] = t[246] ^ x[37];
  assign t[204] = t[247] ^ x[39];
  assign t[205] = t[248] ^ x[40];
  assign t[206] = t[249] ^ x[42];
  assign t[207] = t[250] ^ x[43];
  assign t[208] = t[251] ^ x[45];
  assign t[209] = t[252] ^ x[46];
  assign t[20] = ~(t[22] | t[23]);
  assign t[210] = t[253] ^ x[51];
  assign t[211] = t[254] ^ x[52];
  assign t[212] = t[255] ^ x[57];
  assign t[213] = t[256] ^ x[58];
  assign t[214] = t[257] ^ x[59];
  assign t[215] = t[258] ^ x[61];
  assign t[216] = t[259] ^ x[64];
  assign t[217] = t[260] ^ x[65];
  assign t[218] = t[261] ^ x[66];
  assign t[219] = t[262] ^ x[67];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[68];
  assign t[221] = t[264] ^ x[69];
  assign t[222] = t[265] ^ x[71];
  assign t[223] = t[266] ^ x[74];
  assign t[224] = t[267] ^ x[75];
  assign t[225] = t[268] ^ x[76];
  assign t[226] = t[269] ^ x[77];
  assign t[227] = t[270] ^ x[78];
  assign t[228] = t[271] ^ x[79];
  assign t[229] = t[272] ^ x[81];
  assign t[22] = ~(t[26] | t[27]);
  assign t[230] = t[273] ^ x[84];
  assign t[231] = t[274] ^ x[85];
  assign t[232] = t[275] ^ x[86];
  assign t[233] = t[276] ^ x[87];
  assign t[234] = t[277] ^ x[88];
  assign t[235] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[236] = (x[0]);
  assign t[237] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[238] = (x[9]);
  assign t[239] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[23] = ~(t[28] & t[29]);
  assign t[240] = (x[17]);
  assign t[241] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[242] = (x[23]);
  assign t[243] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[244] = (x[29]);
  assign t[245] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[246] = (x[35]);
  assign t[247] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[248] = (x[38]);
  assign t[249] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[24] = ~(t[30] | t[31]);
  assign t[250] = (x[41]);
  assign t[251] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[252] = (x[44]);
  assign t[253] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[254] = (x[47]);
  assign t[255] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[256] = (x[53]);
  assign t[257] = (x[1]);
  assign t[258] = (x[10]);
  assign t[259] = (x[18]);
  assign t[25] = t[32] | t[33];
  assign t[260] = (x[30]);
  assign t[261] = (x[24]);
  assign t[262] = (x[54]);
  assign t[263] = (x[48]);
  assign t[264] = (x[2]);
  assign t[265] = (x[11]);
  assign t[266] = (x[19]);
  assign t[267] = (x[31]);
  assign t[268] = (x[25]);
  assign t[269] = (x[49]);
  assign t[26] = ~(t[30]);
  assign t[270] = (x[55]);
  assign t[271] = (x[3]);
  assign t[272] = (x[12]);
  assign t[273] = (x[20]);
  assign t[274] = (x[32]);
  assign t[275] = (x[26]);
  assign t[276] = (x[50]);
  assign t[277] = (x[56]);
  assign t[27] = t[101] ? t[35] : t[34];
  assign t[28] = ~(t[36] | t[37]);
  assign t[29] = ~(t[38] & t[39]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[103]);
  assign t[31] = t[101] ? t[41] : t[40];
  assign t[32] = ~(t[26] | t[42]);
  assign t[33] = ~(t[43]);
  assign t[34] = ~(t[44] & t[104]);
  assign t[35] = ~(t[45] & t[46]);
  assign t[36] = ~(t[26] | t[47]);
  assign t[37] = ~(t[26] | t[48]);
  assign t[38] = t[104] & t[49];
  assign t[39] = t[45] | t[44];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(x[7] & t[50]);
  assign t[41] = ~(t[51] & t[46]);
  assign t[42] = t[101] ? t[53] : t[52];
  assign t[43] = ~(t[49] & t[54]);
  assign t[44] = x[7] & t[102];
  assign t[45] = ~(x[7] | t[102]);
  assign t[46] = ~(t[104]);
  assign t[47] = t[101] ? t[34] : t[35];
  assign t[48] = t[101] ? t[40] : t[55];
  assign t[49] = ~(t[30] | t[101]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[102] | t[104]);
  assign t[51] = ~(x[7] | t[56]);
  assign t[52] = ~(t[44] & t[46]);
  assign t[53] = ~(t[45] & t[104]);
  assign t[54] = ~(t[55] & t[57]);
  assign t[55] = ~(t[104] & t[51]);
  assign t[56] = ~(t[102]);
  assign t[57] = ~(x[7] & t[58]);
  assign t[58] = ~(t[102] | t[46]);
  assign t[59] = t[6] ? t[60] : t[107];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = x[6] ? t[62] : t[61];
  assign t[61] = x[7] ? t[64] : t[63];
  assign t[62] = t[65] ^ x[60];
  assign t[63] = t[66] ^ t[67];
  assign t[64] = ~(t[108] ^ t[68]);
  assign t[65] = x[62] ^ x[63];
  assign t[66] = t[69] ? x[62] : x[63];
  assign t[67] = ~(t[109] ^ t[70]);
  assign t[68] = ~(t[110] ^ t[111]);
  assign t[69] = ~(t[71]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[112] ^ t[113]);
  assign t[71] = ~(t[103]);
  assign t[72] = t[6] ? t[73] : t[114];
  assign t[73] = x[6] ? t[75] : t[74];
  assign t[74] = x[7] ? t[77] : t[76];
  assign t[75] = t[78] ^ x[70];
  assign t[76] = t[79] ^ t[80];
  assign t[77] = ~(t[115] ^ t[81]);
  assign t[78] = x[72] ^ x[73];
  assign t[79] = t[82] ? x[72] : x[73];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[116] ^ t[83]);
  assign t[81] = ~(t[117] ^ t[118]);
  assign t[82] = ~(t[71]);
  assign t[83] = ~(t[119] ^ t[120]);
  assign t[84] = t[6] ? t[85] : t[121];
  assign t[85] = x[6] ? t[87] : t[86];
  assign t[86] = x[7] ? t[89] : t[88];
  assign t[87] = t[90] ^ x[80];
  assign t[88] = t[91] ^ t[92];
  assign t[89] = ~(t[122] ^ t[93]);
  assign t[8] = ~(t[97] ^ t[14]);
  assign t[90] = x[82] ^ x[83];
  assign t[91] = t[94] ? x[83] : x[82];
  assign t[92] = ~(t[123] ^ t[95]);
  assign t[93] = ~(t[124] ^ t[125]);
  assign t[94] = ~(t[71]);
  assign t[95] = ~(t[126] ^ t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[59] & ~t[72] & ~t[84]) | (~t[0] & t[59] & ~t[72] & ~t[84]) | (~t[0] & ~t[59] & t[72] & ~t[84]) | (~t[0] & ~t[59] & ~t[72] & t[84]) | (t[0] & t[59] & t[72] & ~t[84]) | (t[0] & t[59] & ~t[72] & t[84]) | (t[0] & ~t[59] & t[72] & t[84]) | (~t[0] & t[59] & t[72] & t[84]);
endmodule

module R2ind116(x, y);
 input [58:0] x;
 output y;

 wire [94:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[23] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[15] ? x[28] : x[27];
  assign t[13] = ~(t[24] ^ t[16]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[15] = ~(t[17]);
  assign t[16] = ~(t[27] ^ t[28]);
  assign t[17] = ~(t[21]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = t[40] ^ x[5];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[11];
  assign t[31] = t[42] ^ x[14];
  assign t[32] = t[43] ^ x[17];
  assign t[33] = t[44] ^ x[20];
  assign t[34] = t[45] ^ x[26];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[40];
  assign t[37] = t[48] ^ x[46];
  assign t[38] = t[49] ^ x[52];
  assign t[39] = t[50] ^ x[58];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[51] & t[52]);
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[6]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = t[73] ^ x[4];
  assign t[52] = t[74] ^ x[5];
  assign t[53] = t[75] ^ x[10];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[16];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[19];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[25];
  assign t[62] = t[84] ^ x[26];
  assign t[63] = t[85] ^ x[33];
  assign t[64] = t[86] ^ x[34];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[45];
  assign t[68] = t[90] ^ x[46];
  assign t[69] = t[91] ^ x[51];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[52];
  assign t[71] = t[93] ^ x[57];
  assign t[72] = t[94] ^ x[58];
  assign t[73] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[74] = (x[3]);
  assign t[75] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[9]);
  assign t[77] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[12]);
  assign t[79] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[15]);
  assign t[81] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[18]);
  assign t[83] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[84] = (x[24]);
  assign t[85] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[86] = (x[32]);
  assign t[87] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[44]);
  assign t[91] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[92] = (x[50]);
  assign t[93] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[94] = (x[56]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [58:0] x;
 output y;

 wire [94:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[23] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[15] ? x[27] : x[28];
  assign t[13] = ~(t[24] ^ t[16]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[15] = ~(t[17]);
  assign t[16] = ~(t[27] ^ t[28]);
  assign t[17] = ~(t[21]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = t[40] ^ x[5];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[11];
  assign t[31] = t[42] ^ x[14];
  assign t[32] = t[43] ^ x[17];
  assign t[33] = t[44] ^ x[20];
  assign t[34] = t[45] ^ x[26];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[40];
  assign t[37] = t[48] ^ x[46];
  assign t[38] = t[49] ^ x[52];
  assign t[39] = t[50] ^ x[58];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[51] & t[52]);
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[6]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = t[73] ^ x[4];
  assign t[52] = t[74] ^ x[5];
  assign t[53] = t[75] ^ x[10];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[16];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[19];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[25];
  assign t[62] = t[84] ^ x[26];
  assign t[63] = t[85] ^ x[33];
  assign t[64] = t[86] ^ x[34];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[45];
  assign t[68] = t[90] ^ x[46];
  assign t[69] = t[91] ^ x[51];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[52];
  assign t[71] = t[93] ^ x[57];
  assign t[72] = t[94] ^ x[58];
  assign t[73] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[74] = (x[2]);
  assign t[75] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[9]);
  assign t[77] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[12]);
  assign t[79] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[15]);
  assign t[81] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[18]);
  assign t[83] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[84] = (x[23]);
  assign t[85] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[86] = (x[31]);
  assign t[87] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[88] = (x[37]);
  assign t[89] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[43]);
  assign t[91] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[92] = (x[49]);
  assign t[93] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[94] = (x[55]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [58:0] x;
 output y;

 wire [94:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[23] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[15] ? x[27] : x[28];
  assign t[13] = ~(t[24] ^ t[16]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[15] = ~(t[17]);
  assign t[16] = ~(t[27] ^ t[28]);
  assign t[17] = ~(t[21]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = t[40] ^ x[5];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[11];
  assign t[31] = t[42] ^ x[14];
  assign t[32] = t[43] ^ x[17];
  assign t[33] = t[44] ^ x[20];
  assign t[34] = t[45] ^ x[26];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[40];
  assign t[37] = t[48] ^ x[46];
  assign t[38] = t[49] ^ x[52];
  assign t[39] = t[50] ^ x[58];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[51] & t[52]);
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[6]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = t[73] ^ x[4];
  assign t[52] = t[74] ^ x[5];
  assign t[53] = t[75] ^ x[10];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[16];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[19];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[25];
  assign t[62] = t[84] ^ x[26];
  assign t[63] = t[85] ^ x[33];
  assign t[64] = t[86] ^ x[34];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[45];
  assign t[68] = t[90] ^ x[46];
  assign t[69] = t[91] ^ x[51];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[52];
  assign t[71] = t[93] ^ x[57];
  assign t[72] = t[94] ^ x[58];
  assign t[73] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[74] = (x[1]);
  assign t[75] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[9]);
  assign t[77] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[12]);
  assign t[79] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[15]);
  assign t[81] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[18]);
  assign t[83] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[84] = (x[22]);
  assign t[85] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[86] = (x[30]);
  assign t[87] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[88] = (x[36]);
  assign t[89] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[42]);
  assign t[91] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[92] = (x[48]);
  assign t[93] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[94] = (x[54]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [58:0] x;
 output y;

 wire [135:0] t;
  assign t[0] = t[1] ? t[2] : t[59];
  assign t[100] = t[122] ^ x[33];
  assign t[101] = t[123] ^ x[34];
  assign t[102] = t[124] ^ x[36];
  assign t[103] = t[125] ^ x[37];
  assign t[104] = t[126] ^ x[39];
  assign t[105] = t[127] ^ x[40];
  assign t[106] = t[128] ^ x[42];
  assign t[107] = t[129] ^ x[43];
  assign t[108] = t[130] ^ x[45];
  assign t[109] = t[131] ^ x[46];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[132] ^ x[51];
  assign t[111] = t[133] ^ x[52];
  assign t[112] = t[134] ^ x[57];
  assign t[113] = t[135] ^ x[58];
  assign t[114] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[115] = (x[0]);
  assign t[116] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[117] = (x[9]);
  assign t[118] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[119] = (x[17]);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[121] = (x[23]);
  assign t[122] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[123] = (x[29]);
  assign t[124] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[125] = (x[35]);
  assign t[126] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[38]);
  assign t[128] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[41]);
  assign t[12] = ~(t[61] ^ t[17]);
  assign t[130] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[44]);
  assign t[132] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[133] = (x[47]);
  assign t[134] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[135] = (x[53]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[62] ^ t[63]);
  assign t[15] = ~(t[64] & t[65]);
  assign t[16] = ~(t[66] & t[67]);
  assign t[17] = ~(t[68] ^ t[69]);
  assign t[18] = t[66] ? x[15] : x[16];
  assign t[19] = ~(t[20] & t[21]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[22] | t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[28] & t[29]);
  assign t[24] = ~(t[30] | t[31]);
  assign t[25] = t[32] | t[33];
  assign t[26] = ~(t[30]);
  assign t[27] = t[64] ? t[35] : t[34];
  assign t[28] = ~(t[36] | t[37]);
  assign t[29] = ~(t[38] & t[39]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[66]);
  assign t[31] = t[64] ? t[41] : t[40];
  assign t[32] = ~(t[26] | t[42]);
  assign t[33] = ~(t[43]);
  assign t[34] = ~(t[44] & t[67]);
  assign t[35] = ~(t[45] & t[46]);
  assign t[36] = ~(t[26] | t[47]);
  assign t[37] = ~(t[26] | t[48]);
  assign t[38] = t[67] & t[49];
  assign t[39] = t[45] | t[44];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(x[7] & t[50]);
  assign t[41] = ~(t[51] & t[46]);
  assign t[42] = t[64] ? t[53] : t[52];
  assign t[43] = ~(t[49] & t[54]);
  assign t[44] = x[7] & t[65];
  assign t[45] = ~(x[7] | t[65]);
  assign t[46] = ~(t[67]);
  assign t[47] = t[64] ? t[34] : t[35];
  assign t[48] = t[64] ? t[40] : t[55];
  assign t[49] = ~(t[30] | t[64]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[65] | t[67]);
  assign t[51] = ~(x[7] | t[56]);
  assign t[52] = ~(t[44] & t[46]);
  assign t[53] = ~(t[45] & t[67]);
  assign t[54] = ~(t[55] & t[57]);
  assign t[55] = ~(t[67] & t[51]);
  assign t[56] = ~(t[65]);
  assign t[57] = ~(x[7] & t[58]);
  assign t[58] = ~(t[65] | t[46]);
  assign t[59] = (t[70]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = (t[73]);
  assign t[63] = (t[74]);
  assign t[64] = (t[75]);
  assign t[65] = (t[76]);
  assign t[66] = (t[77]);
  assign t[67] = (t[78]);
  assign t[68] = (t[79]);
  assign t[69] = (t[80]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[81] ^ x[5];
  assign t[71] = t[82] ^ x[14];
  assign t[72] = t[83] ^ x[22];
  assign t[73] = t[84] ^ x[28];
  assign t[74] = t[85] ^ x[34];
  assign t[75] = t[86] ^ x[37];
  assign t[76] = t[87] ^ x[40];
  assign t[77] = t[88] ^ x[43];
  assign t[78] = t[89] ^ x[46];
  assign t[79] = t[90] ^ x[52];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[91] ^ x[58];
  assign t[81] = (~t[92] & t[93]);
  assign t[82] = (~t[94] & t[95]);
  assign t[83] = (~t[96] & t[97]);
  assign t[84] = (~t[98] & t[99]);
  assign t[85] = (~t[100] & t[101]);
  assign t[86] = (~t[102] & t[103]);
  assign t[87] = (~t[104] & t[105]);
  assign t[88] = (~t[106] & t[107]);
  assign t[89] = (~t[108] & t[109]);
  assign t[8] = ~(t[60] ^ t[14]);
  assign t[90] = (~t[110] & t[111]);
  assign t[91] = (~t[112] & t[113]);
  assign t[92] = t[114] ^ x[4];
  assign t[93] = t[115] ^ x[5];
  assign t[94] = t[116] ^ x[13];
  assign t[95] = t[117] ^ x[14];
  assign t[96] = t[118] ^ x[21];
  assign t[97] = t[119] ^ x[22];
  assign t[98] = t[120] ^ x[27];
  assign t[99] = t[121] ^ x[28];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [61:0] x;
 output y;

 wire [191:0] t;
  assign t[0] = t[1] ? t[2] : t[76];
  assign t[100] = t[120] ^ x[20];
  assign t[101] = t[121] ^ x[26];
  assign t[102] = t[122] ^ x[34];
  assign t[103] = t[123] ^ x[40];
  assign t[104] = t[124] ^ x[41];
  assign t[105] = t[125] ^ x[43];
  assign t[106] = t[126] ^ x[46];
  assign t[107] = t[127] ^ x[47];
  assign t[108] = t[128] ^ x[48];
  assign t[109] = t[129] ^ x[50];
  assign t[10] = ~(t[81] ^ t[13]);
  assign t[110] = t[130] ^ x[53];
  assign t[111] = t[131] ^ x[54];
  assign t[112] = t[132] ^ x[55];
  assign t[113] = t[133] ^ x[57];
  assign t[114] = t[134] ^ x[60];
  assign t[115] = t[135] ^ x[61];
  assign t[116] = (~t[136] & t[137]);
  assign t[117] = (~t[138] & t[139]);
  assign t[118] = (~t[140] & t[141]);
  assign t[119] = (~t[142] & t[143]);
  assign t[11] = x[27] ^ x[28];
  assign t[120] = (~t[144] & t[145]);
  assign t[121] = (~t[146] & t[147]);
  assign t[122] = (~t[148] & t[149]);
  assign t[123] = (~t[150] & t[151]);
  assign t[124] = (~t[136] & t[152]);
  assign t[125] = (~t[146] & t[153]);
  assign t[126] = (~t[150] & t[154]);
  assign t[127] = (~t[148] & t[155]);
  assign t[128] = (~t[136] & t[156]);
  assign t[129] = (~t[146] & t[157]);
  assign t[12] = ~(t[14] ^ t[15]);
  assign t[130] = (~t[150] & t[158]);
  assign t[131] = (~t[148] & t[159]);
  assign t[132] = (~t[136] & t[160]);
  assign t[133] = (~t[146] & t[161]);
  assign t[134] = (~t[150] & t[162]);
  assign t[135] = (~t[148] & t[163]);
  assign t[136] = t[164] ^ x[4];
  assign t[137] = t[165] ^ x[5];
  assign t[138] = t[166] ^ x[10];
  assign t[139] = t[167] ^ x[11];
  assign t[13] = ~(t[82] ^ t[83]);
  assign t[140] = t[168] ^ x[13];
  assign t[141] = t[169] ^ x[14];
  assign t[142] = t[170] ^ x[16];
  assign t[143] = t[171] ^ x[17];
  assign t[144] = t[172] ^ x[19];
  assign t[145] = t[173] ^ x[20];
  assign t[146] = t[174] ^ x[25];
  assign t[147] = t[175] ^ x[26];
  assign t[148] = t[176] ^ x[33];
  assign t[149] = t[177] ^ x[34];
  assign t[14] = t[79] ? x[28] : x[27];
  assign t[150] = t[178] ^ x[39];
  assign t[151] = t[179] ^ x[40];
  assign t[152] = t[180] ^ x[41];
  assign t[153] = t[181] ^ x[43];
  assign t[154] = t[182] ^ x[46];
  assign t[155] = t[183] ^ x[47];
  assign t[156] = t[184] ^ x[48];
  assign t[157] = t[185] ^ x[50];
  assign t[158] = t[186] ^ x[53];
  assign t[159] = t[187] ^ x[54];
  assign t[15] = t[16] | t[17];
  assign t[160] = t[188] ^ x[55];
  assign t[161] = t[189] ^ x[57];
  assign t[162] = t[190] ^ x[60];
  assign t[163] = t[191] ^ x[61];
  assign t[164] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[165] = (x[0]);
  assign t[166] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[167] = (x[9]);
  assign t[168] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[169] = (x[12]);
  assign t[16] = ~(t[18] & t[19]);
  assign t[170] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[171] = (x[15]);
  assign t[172] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[173] = (x[18]);
  assign t[174] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[175] = (x[21]);
  assign t[176] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[177] = (x[29]);
  assign t[178] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[179] = (x[35]);
  assign t[17] = ~(t[20] & t[21]);
  assign t[180] = (x[1]);
  assign t[181] = (x[22]);
  assign t[182] = (x[36]);
  assign t[183] = (x[30]);
  assign t[184] = (x[2]);
  assign t[185] = (x[23]);
  assign t[186] = (x[37]);
  assign t[187] = (x[31]);
  assign t[188] = (x[3]);
  assign t[189] = (x[24]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[190] = (x[38]);
  assign t[191] = (x[32]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[26] | t[27]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[30] | t[77]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = ~(t[78] | t[33]);
  assign t[25] = t[34] & t[77];
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[34] | t[36]);
  assign t[28] = ~(t[34] | t[37]);
  assign t[29] = ~(t[34] | t[38]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = ~(t[79]);
  assign t[31] = ~(t[80] & t[39]);
  assign t[32] = ~(x[7] & t[24]);
  assign t[33] = ~(t[80]);
  assign t[34] = ~(t[30]);
  assign t[35] = t[77] ? t[41] : t[40];
  assign t[36] = t[77] ? t[43] : t[42];
  assign t[37] = t[77] ? t[44] : t[31];
  assign t[38] = t[77] ? t[42] : t[43];
  assign t[39] = ~(x[7] | t[45]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[46] & t[80]);
  assign t[41] = ~(t[47] & t[33]);
  assign t[42] = ~(t[46] & t[33]);
  assign t[43] = ~(t[47] & t[80]);
  assign t[44] = ~(x[7] & t[48]);
  assign t[45] = ~(t[78]);
  assign t[46] = x[7] & t[78];
  assign t[47] = ~(x[7] | t[78]);
  assign t[48] = ~(t[78] | t[80]);
  assign t[49] = t[1] ? t[50] : t[84];
  assign t[4] = ~(x[6]);
  assign t[50] = x[6] ? t[52] : t[51];
  assign t[51] = x[7] ? t[54] : t[53];
  assign t[52] = t[55] ^ x[42];
  assign t[53] = t[56] ^ t[54];
  assign t[54] = ~(t[85] ^ t[57]);
  assign t[55] = x[44] ^ x[45];
  assign t[56] = t[79] ? x[45] : x[44];
  assign t[57] = ~(t[86] ^ t[87]);
  assign t[58] = t[1] ? t[59] : t[88];
  assign t[59] = x[6] ? t[61] : t[60];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = x[7] ? t[63] : t[62];
  assign t[61] = t[64] ^ x[49];
  assign t[62] = t[65] ^ t[63];
  assign t[63] = ~(t[89] ^ t[66]);
  assign t[64] = x[51] ^ x[52];
  assign t[65] = t[79] ? x[51] : x[52];
  assign t[66] = ~(t[90] ^ t[91]);
  assign t[67] = t[1] ? t[68] : t[92];
  assign t[68] = x[6] ? t[70] : t[69];
  assign t[69] = x[7] ? t[72] : t[71];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[73] ^ x[56];
  assign t[71] = t[74] ^ t[72];
  assign t[72] = ~(t[93] ^ t[75]);
  assign t[73] = x[58] ^ x[59];
  assign t[74] = t[79] ? x[58] : x[59];
  assign t[75] = ~(t[94] ^ t[95]);
  assign t[76] = (t[96]);
  assign t[77] = (t[97]);
  assign t[78] = (t[98]);
  assign t[79] = (t[99]);
  assign t[7] = ~(t[77] & t[78]);
  assign t[80] = (t[100]);
  assign t[81] = (t[101]);
  assign t[82] = (t[102]);
  assign t[83] = (t[103]);
  assign t[84] = (t[104]);
  assign t[85] = (t[105]);
  assign t[86] = (t[106]);
  assign t[87] = (t[107]);
  assign t[88] = (t[108]);
  assign t[89] = (t[109]);
  assign t[8] = ~(t[79] & t[80]);
  assign t[90] = (t[110]);
  assign t[91] = (t[111]);
  assign t[92] = (t[112]);
  assign t[93] = (t[113]);
  assign t[94] = (t[114]);
  assign t[95] = (t[115]);
  assign t[96] = t[116] ^ x[5];
  assign t[97] = t[117] ^ x[11];
  assign t[98] = t[118] ^ x[14];
  assign t[99] = t[119] ^ x[17];
  assign t[9] = ~(t[10] ^ t[12]);
  assign y = (t[0] & ~t[49] & ~t[58] & ~t[67]) | (~t[0] & t[49] & ~t[58] & ~t[67]) | (~t[0] & ~t[49] & t[58] & ~t[67]) | (~t[0] & ~t[49] & ~t[58] & t[67]) | (t[0] & t[49] & t[58] & ~t[67]) | (t[0] & t[49] & ~t[58] & t[67]) | (t[0] & ~t[49] & t[58] & t[67]) | (~t[0] & t[49] & t[58] & t[67]);
endmodule

module R2ind121(x, y);
 input [40:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = t[1] ? t[2] : t[14];
  assign t[10] = ~(t[19] ^ t[13]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[17] ? x[27] : x[28];
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[11];
  assign t[24] = t[32] ^ x[14];
  assign t[25] = t[33] ^ x[17];
  assign t[26] = t[34] ^ x[20];
  assign t[27] = t[35] ^ x[26];
  assign t[28] = t[36] ^ x[34];
  assign t[29] = t[37] ^ x[40];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = (~t[38] & t[39]);
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = t[54] ^ x[4];
  assign t[39] = t[55] ^ x[5];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[56] ^ x[10];
  assign t[41] = t[57] ^ x[11];
  assign t[42] = t[58] ^ x[13];
  assign t[43] = t[59] ^ x[14];
  assign t[44] = t[60] ^ x[16];
  assign t[45] = t[61] ^ x[17];
  assign t[46] = t[62] ^ x[19];
  assign t[47] = t[63] ^ x[20];
  assign t[48] = t[64] ^ x[25];
  assign t[49] = t[65] ^ x[26];
  assign t[4] = ~(x[6]);
  assign t[50] = t[66] ^ x[33];
  assign t[51] = t[67] ^ x[34];
  assign t[52] = t[68] ^ x[39];
  assign t[53] = t[69] ^ x[40];
  assign t[54] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[55] = (x[3]);
  assign t[56] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[9]);
  assign t[58] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[12]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[15]);
  assign t[62] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[18]);
  assign t[64] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[65] = (x[24]);
  assign t[66] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[67] = (x[32]);
  assign t[68] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[69] = (x[38]);
  assign t[6] = t[11] ^ x[8];
  assign t[7] = ~(t[15] & t[16]);
  assign t[8] = ~(t[17] & t[18]);
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [40:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = t[1] ? t[2] : t[14];
  assign t[10] = ~(t[19] ^ t[13]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[17] ? x[27] : x[28];
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[11];
  assign t[24] = t[32] ^ x[14];
  assign t[25] = t[33] ^ x[17];
  assign t[26] = t[34] ^ x[20];
  assign t[27] = t[35] ^ x[26];
  assign t[28] = t[36] ^ x[34];
  assign t[29] = t[37] ^ x[40];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = (~t[38] & t[39]);
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = t[54] ^ x[4];
  assign t[39] = t[55] ^ x[5];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[56] ^ x[10];
  assign t[41] = t[57] ^ x[11];
  assign t[42] = t[58] ^ x[13];
  assign t[43] = t[59] ^ x[14];
  assign t[44] = t[60] ^ x[16];
  assign t[45] = t[61] ^ x[17];
  assign t[46] = t[62] ^ x[19];
  assign t[47] = t[63] ^ x[20];
  assign t[48] = t[64] ^ x[25];
  assign t[49] = t[65] ^ x[26];
  assign t[4] = ~(x[6]);
  assign t[50] = t[66] ^ x[33];
  assign t[51] = t[67] ^ x[34];
  assign t[52] = t[68] ^ x[39];
  assign t[53] = t[69] ^ x[40];
  assign t[54] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[55] = (x[2]);
  assign t[56] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[9]);
  assign t[58] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[12]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[15]);
  assign t[62] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[18]);
  assign t[64] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[65] = (x[23]);
  assign t[66] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[67] = (x[31]);
  assign t[68] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[69] = (x[37]);
  assign t[6] = t[11] ^ x[8];
  assign t[7] = ~(t[15] & t[16]);
  assign t[8] = ~(t[17] & t[18]);
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [40:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = t[1] ? t[2] : t[14];
  assign t[10] = ~(t[19] ^ t[13]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[17] ? x[28] : x[27];
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[11];
  assign t[24] = t[32] ^ x[14];
  assign t[25] = t[33] ^ x[17];
  assign t[26] = t[34] ^ x[20];
  assign t[27] = t[35] ^ x[26];
  assign t[28] = t[36] ^ x[34];
  assign t[29] = t[37] ^ x[40];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = (~t[38] & t[39]);
  assign t[31] = (~t[40] & t[41]);
  assign t[32] = (~t[42] & t[43]);
  assign t[33] = (~t[44] & t[45]);
  assign t[34] = (~t[46] & t[47]);
  assign t[35] = (~t[48] & t[49]);
  assign t[36] = (~t[50] & t[51]);
  assign t[37] = (~t[52] & t[53]);
  assign t[38] = t[54] ^ x[4];
  assign t[39] = t[55] ^ x[5];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = t[56] ^ x[10];
  assign t[41] = t[57] ^ x[11];
  assign t[42] = t[58] ^ x[13];
  assign t[43] = t[59] ^ x[14];
  assign t[44] = t[60] ^ x[16];
  assign t[45] = t[61] ^ x[17];
  assign t[46] = t[62] ^ x[19];
  assign t[47] = t[63] ^ x[20];
  assign t[48] = t[64] ^ x[25];
  assign t[49] = t[65] ^ x[26];
  assign t[4] = ~(x[6]);
  assign t[50] = t[66] ^ x[33];
  assign t[51] = t[67] ^ x[34];
  assign t[52] = t[68] ^ x[39];
  assign t[53] = t[69] ^ x[40];
  assign t[54] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[55] = (x[1]);
  assign t[56] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[57] = (x[9]);
  assign t[58] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[59] = (x[12]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[61] = (x[15]);
  assign t[62] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[18]);
  assign t[64] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[65] = (x[22]);
  assign t[66] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[67] = (x[30]);
  assign t[68] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[69] = (x[36]);
  assign t[6] = t[11] ^ x[8];
  assign t[7] = ~(t[15] & t[16]);
  assign t[8] = ~(t[17] & t[18]);
  assign t[9] = t[12] ^ t[10];
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [40:0] x;
 output y;

 wire [104:0] t;
  assign t[0] = t[1] ? t[2] : t[49];
  assign t[100] = (x[21]);
  assign t[101] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[102] = (x[29]);
  assign t[103] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[104] = (x[35]);
  assign t[10] = ~(t[54] ^ t[13]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = ~(t[14] ^ t[15]);
  assign t[13] = ~(t[55] ^ t[56]);
  assign t[14] = t[52] ? x[28] : x[27];
  assign t[15] = t[16] | t[17];
  assign t[16] = ~(t[18] & t[19]);
  assign t[17] = ~(t[20] & t[21]);
  assign t[18] = ~(t[22] & t[23]);
  assign t[19] = ~(t[24] & t[25]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[26] | t[27]);
  assign t[21] = ~(t[28] | t[29]);
  assign t[22] = ~(t[30] | t[50]);
  assign t[23] = ~(t[31] & t[32]);
  assign t[24] = ~(t[51] | t[33]);
  assign t[25] = t[34] & t[50];
  assign t[26] = ~(t[34] | t[35]);
  assign t[27] = ~(t[34] | t[36]);
  assign t[28] = ~(t[34] | t[37]);
  assign t[29] = ~(t[34] | t[38]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = ~(t[52]);
  assign t[31] = ~(t[53] & t[39]);
  assign t[32] = ~(x[7] & t[24]);
  assign t[33] = ~(t[53]);
  assign t[34] = ~(t[30]);
  assign t[35] = t[50] ? t[41] : t[40];
  assign t[36] = t[50] ? t[43] : t[42];
  assign t[37] = t[50] ? t[44] : t[31];
  assign t[38] = t[50] ? t[42] : t[43];
  assign t[39] = ~(x[7] | t[45]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[46] & t[53]);
  assign t[41] = ~(t[47] & t[33]);
  assign t[42] = ~(t[46] & t[33]);
  assign t[43] = ~(t[47] & t[53]);
  assign t[44] = ~(x[7] & t[48]);
  assign t[45] = ~(t[51]);
  assign t[46] = x[7] & t[51];
  assign t[47] = ~(x[7] | t[51]);
  assign t[48] = ~(t[51] | t[53]);
  assign t[49] = (t[57]);
  assign t[4] = ~(x[6]);
  assign t[50] = (t[58]);
  assign t[51] = (t[59]);
  assign t[52] = (t[60]);
  assign t[53] = (t[61]);
  assign t[54] = (t[62]);
  assign t[55] = (t[63]);
  assign t[56] = (t[64]);
  assign t[57] = t[65] ^ x[5];
  assign t[58] = t[66] ^ x[11];
  assign t[59] = t[67] ^ x[14];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[68] ^ x[17];
  assign t[61] = t[69] ^ x[20];
  assign t[62] = t[70] ^ x[26];
  assign t[63] = t[71] ^ x[34];
  assign t[64] = t[72] ^ x[40];
  assign t[65] = (~t[73] & t[74]);
  assign t[66] = (~t[75] & t[76]);
  assign t[67] = (~t[77] & t[78]);
  assign t[68] = (~t[79] & t[80]);
  assign t[69] = (~t[81] & t[82]);
  assign t[6] = t[11] ^ x[8];
  assign t[70] = (~t[83] & t[84]);
  assign t[71] = (~t[85] & t[86]);
  assign t[72] = (~t[87] & t[88]);
  assign t[73] = t[89] ^ x[4];
  assign t[74] = t[90] ^ x[5];
  assign t[75] = t[91] ^ x[10];
  assign t[76] = t[92] ^ x[11];
  assign t[77] = t[93] ^ x[13];
  assign t[78] = t[94] ^ x[14];
  assign t[79] = t[95] ^ x[16];
  assign t[7] = ~(t[50] & t[51]);
  assign t[80] = t[96] ^ x[17];
  assign t[81] = t[97] ^ x[19];
  assign t[82] = t[98] ^ x[20];
  assign t[83] = t[99] ^ x[25];
  assign t[84] = t[100] ^ x[26];
  assign t[85] = t[101] ^ x[33];
  assign t[86] = t[102] ^ x[34];
  assign t[87] = t[103] ^ x[39];
  assign t[88] = t[104] ^ x[40];
  assign t[89] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[8] = ~(t[52] & t[53]);
  assign t[90] = (x[0]);
  assign t[91] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[9]);
  assign t[93] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[12]);
  assign t[95] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[96] = (x[15]);
  assign t[97] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[98] = (x[18]);
  assign t[99] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[9] = ~(t[10] ^ t[12]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [88:0] x;
 output y;

 wire [265:0] t;
  assign t[0] = t[1] ? t[2] : t[84];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[89] ^ t[14]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = t[148] ^ x[5];
  assign t[117] = t[149] ^ x[11];
  assign t[118] = t[150] ^ x[14];
  assign t[119] = t[151] ^ x[17];
  assign t[11] = x[27] ^ x[28];
  assign t[120] = t[152] ^ x[20];
  assign t[121] = t[153] ^ x[26];
  assign t[122] = t[154] ^ x[34];
  assign t[123] = t[155] ^ x[40];
  assign t[124] = t[156] ^ x[46];
  assign t[125] = t[157] ^ x[52];
  assign t[126] = t[158] ^ x[58];
  assign t[127] = t[159] ^ x[59];
  assign t[128] = t[160] ^ x[61];
  assign t[129] = t[161] ^ x[64];
  assign t[12] = ~(t[90] ^ t[15]);
  assign t[130] = t[162] ^ x[65];
  assign t[131] = t[163] ^ x[66];
  assign t[132] = t[164] ^ x[67];
  assign t[133] = t[165] ^ x[68];
  assign t[134] = t[166] ^ x[69];
  assign t[135] = t[167] ^ x[71];
  assign t[136] = t[168] ^ x[74];
  assign t[137] = t[169] ^ x[75];
  assign t[138] = t[170] ^ x[76];
  assign t[139] = t[171] ^ x[77];
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[140] = t[172] ^ x[78];
  assign t[141] = t[173] ^ x[79];
  assign t[142] = t[174] ^ x[81];
  assign t[143] = t[175] ^ x[84];
  assign t[144] = t[176] ^ x[85];
  assign t[145] = t[177] ^ x[86];
  assign t[146] = t[178] ^ x[87];
  assign t[147] = t[179] ^ x[88];
  assign t[148] = (~t[180] & t[181]);
  assign t[149] = (~t[182] & t[183]);
  assign t[14] = ~(t[91] ^ t[92]);
  assign t[150] = (~t[184] & t[185]);
  assign t[151] = (~t[186] & t[187]);
  assign t[152] = (~t[188] & t[189]);
  assign t[153] = (~t[190] & t[191]);
  assign t[154] = (~t[192] & t[193]);
  assign t[155] = (~t[194] & t[195]);
  assign t[156] = (~t[196] & t[197]);
  assign t[157] = (~t[198] & t[199]);
  assign t[158] = (~t[200] & t[201]);
  assign t[159] = (~t[180] & t[202]);
  assign t[15] = ~(t[93] ^ t[94]);
  assign t[160] = (~t[190] & t[203]);
  assign t[161] = (~t[192] & t[204]);
  assign t[162] = (~t[196] & t[205]);
  assign t[163] = (~t[194] & t[206]);
  assign t[164] = (~t[200] & t[207]);
  assign t[165] = (~t[198] & t[208]);
  assign t[166] = (~t[180] & t[209]);
  assign t[167] = (~t[190] & t[210]);
  assign t[168] = (~t[192] & t[211]);
  assign t[169] = (~t[194] & t[212]);
  assign t[16] = t[18] ? x[27] : x[28];
  assign t[170] = (~t[196] & t[213]);
  assign t[171] = (~t[200] & t[214]);
  assign t[172] = (~t[198] & t[215]);
  assign t[173] = (~t[180] & t[216]);
  assign t[174] = (~t[190] & t[217]);
  assign t[175] = (~t[192] & t[218]);
  assign t[176] = (~t[194] & t[219]);
  assign t[177] = (~t[196] & t[220]);
  assign t[178] = (~t[200] & t[221]);
  assign t[179] = (~t[198] & t[222]);
  assign t[17] = ~(t[19] & t[20]);
  assign t[180] = t[223] ^ x[4];
  assign t[181] = t[224] ^ x[5];
  assign t[182] = t[225] ^ x[10];
  assign t[183] = t[226] ^ x[11];
  assign t[184] = t[227] ^ x[13];
  assign t[185] = t[228] ^ x[14];
  assign t[186] = t[229] ^ x[16];
  assign t[187] = t[230] ^ x[17];
  assign t[188] = t[231] ^ x[19];
  assign t[189] = t[232] ^ x[20];
  assign t[18] = ~(t[21]);
  assign t[190] = t[233] ^ x[25];
  assign t[191] = t[234] ^ x[26];
  assign t[192] = t[235] ^ x[33];
  assign t[193] = t[236] ^ x[34];
  assign t[194] = t[237] ^ x[39];
  assign t[195] = t[238] ^ x[40];
  assign t[196] = t[239] ^ x[45];
  assign t[197] = t[240] ^ x[46];
  assign t[198] = t[241] ^ x[51];
  assign t[199] = t[242] ^ x[52];
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[200] = t[243] ^ x[57];
  assign t[201] = t[244] ^ x[58];
  assign t[202] = t[245] ^ x[59];
  assign t[203] = t[246] ^ x[61];
  assign t[204] = t[247] ^ x[64];
  assign t[205] = t[248] ^ x[65];
  assign t[206] = t[249] ^ x[66];
  assign t[207] = t[250] ^ x[67];
  assign t[208] = t[251] ^ x[68];
  assign t[209] = t[252] ^ x[69];
  assign t[20] = ~(t[24]);
  assign t[210] = t[253] ^ x[71];
  assign t[211] = t[254] ^ x[74];
  assign t[212] = t[255] ^ x[75];
  assign t[213] = t[256] ^ x[76];
  assign t[214] = t[257] ^ x[77];
  assign t[215] = t[258] ^ x[78];
  assign t[216] = t[259] ^ x[79];
  assign t[217] = t[260] ^ x[81];
  assign t[218] = t[261] ^ x[84];
  assign t[219] = t[262] ^ x[85];
  assign t[21] = ~(t[87]);
  assign t[220] = t[263] ^ x[86];
  assign t[221] = t[264] ^ x[87];
  assign t[222] = t[265] ^ x[88];
  assign t[223] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[224] = (x[0]);
  assign t[225] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[226] = (x[9]);
  assign t[227] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[228] = (x[12]);
  assign t[229] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[22] = ~(t[25] & t[26]);
  assign t[230] = (x[15]);
  assign t[231] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[232] = (x[18]);
  assign t[233] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[234] = (x[21]);
  assign t[235] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[236] = (x[29]);
  assign t[237] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[238] = (x[35]);
  assign t[239] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[23] = ~(t[27] & t[28]);
  assign t[240] = (x[41]);
  assign t[241] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[242] = (x[47]);
  assign t[243] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[244] = (x[53]);
  assign t[245] = (x[1]);
  assign t[246] = (x[22]);
  assign t[247] = (x[30]);
  assign t[248] = (x[42]);
  assign t[249] = (x[36]);
  assign t[24] = ~(t[29] | t[30]);
  assign t[250] = (x[54]);
  assign t[251] = (x[48]);
  assign t[252] = (x[2]);
  assign t[253] = (x[23]);
  assign t[254] = (x[31]);
  assign t[255] = (x[37]);
  assign t[256] = (x[43]);
  assign t[257] = (x[55]);
  assign t[258] = (x[49]);
  assign t[259] = (x[3]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[260] = (x[24]);
  assign t[261] = (x[32]);
  assign t[262] = (x[38]);
  assign t[263] = (x[44]);
  assign t[264] = (x[56]);
  assign t[265] = (x[50]);
  assign t[26] = ~(t[33] & t[34]);
  assign t[27] = ~(t[35]);
  assign t[28] = t[36] | t[37];
  assign t[29] = ~(t[36]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[85] ? t[39] : t[38];
  assign t[31] = ~(t[36] | t[85]);
  assign t[32] = ~(t[40] & t[41]);
  assign t[33] = ~(t[86] | t[42]);
  assign t[34] = t[29] & t[85];
  assign t[35] = ~(t[36] | t[43]);
  assign t[36] = ~(t[87]);
  assign t[37] = t[85] ? t[45] : t[44];
  assign t[38] = ~(t[46] & t[88]);
  assign t[39] = ~(t[47] & t[42]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[88] & t[48]);
  assign t[41] = ~(x[7] & t[33]);
  assign t[42] = ~(t[88]);
  assign t[43] = t[85] ? t[44] : t[45];
  assign t[44] = ~(t[48] & t[42]);
  assign t[45] = ~(x[7] & t[49]);
  assign t[46] = x[7] & t[86];
  assign t[47] = ~(x[7] | t[86]);
  assign t[48] = ~(x[7] | t[50]);
  assign t[49] = ~(t[86] | t[88]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[86]);
  assign t[51] = t[1] ? t[52] : t[95];
  assign t[52] = x[6] ? t[54] : t[53];
  assign t[53] = x[7] ? t[56] : t[55];
  assign t[54] = t[57] ^ x[60];
  assign t[55] = t[58] ^ t[59];
  assign t[56] = ~(t[96] ^ t[60]);
  assign t[57] = x[62] ^ x[63];
  assign t[58] = t[87] ? x[62] : x[63];
  assign t[59] = ~(t[97] ^ t[61]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = ~(t[98] ^ t[99]);
  assign t[61] = ~(t[100] ^ t[101]);
  assign t[62] = t[1] ? t[63] : t[102];
  assign t[63] = x[6] ? t[65] : t[64];
  assign t[64] = x[7] ? t[67] : t[66];
  assign t[65] = t[68] ^ x[70];
  assign t[66] = t[69] ^ t[70];
  assign t[67] = ~(t[103] ^ t[71]);
  assign t[68] = x[72] ^ x[73];
  assign t[69] = t[87] ? x[72] : x[73];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = ~(t[104] ^ t[72]);
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = ~(t[107] ^ t[108]);
  assign t[73] = t[1] ? t[74] : t[109];
  assign t[74] = x[6] ? t[76] : t[75];
  assign t[75] = x[7] ? t[78] : t[77];
  assign t[76] = t[79] ^ x[80];
  assign t[77] = t[80] ^ t[81];
  assign t[78] = ~(t[110] ^ t[82]);
  assign t[79] = x[82] ^ x[83];
  assign t[7] = ~(t[85] & t[86]);
  assign t[80] = t[87] ? x[82] : x[83];
  assign t[81] = ~(t[111] ^ t[83]);
  assign t[82] = ~(t[112] ^ t[113]);
  assign t[83] = ~(t[114] ^ t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[87] & t[88]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0] & ~t[51] & ~t[62] & ~t[73]) | (~t[0] & t[51] & ~t[62] & ~t[73]) | (~t[0] & ~t[51] & t[62] & ~t[73]) | (~t[0] & ~t[51] & ~t[62] & t[73]) | (t[0] & t[51] & t[62] & ~t[73]) | (t[0] & t[51] & ~t[62] & t[73]) | (t[0] & ~t[51] & t[62] & t[73]) | (~t[0] & t[51] & t[62] & t[73]);
endmodule

module R2ind126(x, y);
 input [58:0] x;
 output y;

 wire [92:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[21] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[19] ? x[27] : x[28];
  assign t[13] = ~(t[22] ^ t[15]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] ^ t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[11];
  assign t[29] = t[40] ^ x[14];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[17];
  assign t[31] = t[42] ^ x[20];
  assign t[32] = t[43] ^ x[26];
  assign t[33] = t[44] ^ x[34];
  assign t[34] = t[45] ^ x[40];
  assign t[35] = t[46] ^ x[46];
  assign t[36] = t[47] ^ x[52];
  assign t[37] = t[48] ^ x[58];
  assign t[38] = (~t[49] & t[50]);
  assign t[39] = (~t[51] & t[52]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[53] & t[54]);
  assign t[41] = (~t[55] & t[56]);
  assign t[42] = (~t[57] & t[58]);
  assign t[43] = (~t[59] & t[60]);
  assign t[44] = (~t[61] & t[62]);
  assign t[45] = (~t[63] & t[64]);
  assign t[46] = (~t[65] & t[66]);
  assign t[47] = (~t[67] & t[68]);
  assign t[48] = (~t[69] & t[70]);
  assign t[49] = t[71] ^ x[4];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[5];
  assign t[51] = t[73] ^ x[10];
  assign t[52] = t[74] ^ x[11];
  assign t[53] = t[75] ^ x[13];
  assign t[54] = t[76] ^ x[14];
  assign t[55] = t[77] ^ x[16];
  assign t[56] = t[78] ^ x[17];
  assign t[57] = t[79] ^ x[19];
  assign t[58] = t[80] ^ x[20];
  assign t[59] = t[81] ^ x[25];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[26];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[39];
  assign t[64] = t[86] ^ x[40];
  assign t[65] = t[87] ^ x[45];
  assign t[66] = t[88] ^ x[46];
  assign t[67] = t[89] ^ x[51];
  assign t[68] = t[90] ^ x[52];
  assign t[69] = t[91] ^ x[57];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[58];
  assign t[71] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[72] = (x[3]);
  assign t[73] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[9]);
  assign t[75] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[12]);
  assign t[77] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[15]);
  assign t[79] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[17] & t[18]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[86] = (x[38]);
  assign t[87] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[88] = (x[44]);
  assign t[89] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[8] = ~(t[19] & t[20]);
  assign t[90] = (x[50]);
  assign t[91] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[92] = (x[56]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [58:0] x;
 output y;

 wire [92:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[21] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[19] ? x[27] : x[28];
  assign t[13] = ~(t[22] ^ t[15]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] ^ t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[11];
  assign t[29] = t[40] ^ x[14];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[17];
  assign t[31] = t[42] ^ x[20];
  assign t[32] = t[43] ^ x[26];
  assign t[33] = t[44] ^ x[34];
  assign t[34] = t[45] ^ x[40];
  assign t[35] = t[46] ^ x[46];
  assign t[36] = t[47] ^ x[52];
  assign t[37] = t[48] ^ x[58];
  assign t[38] = (~t[49] & t[50]);
  assign t[39] = (~t[51] & t[52]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[53] & t[54]);
  assign t[41] = (~t[55] & t[56]);
  assign t[42] = (~t[57] & t[58]);
  assign t[43] = (~t[59] & t[60]);
  assign t[44] = (~t[61] & t[62]);
  assign t[45] = (~t[63] & t[64]);
  assign t[46] = (~t[65] & t[66]);
  assign t[47] = (~t[67] & t[68]);
  assign t[48] = (~t[69] & t[70]);
  assign t[49] = t[71] ^ x[4];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[5];
  assign t[51] = t[73] ^ x[10];
  assign t[52] = t[74] ^ x[11];
  assign t[53] = t[75] ^ x[13];
  assign t[54] = t[76] ^ x[14];
  assign t[55] = t[77] ^ x[16];
  assign t[56] = t[78] ^ x[17];
  assign t[57] = t[79] ^ x[19];
  assign t[58] = t[80] ^ x[20];
  assign t[59] = t[81] ^ x[25];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[26];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[39];
  assign t[64] = t[86] ^ x[40];
  assign t[65] = t[87] ^ x[45];
  assign t[66] = t[88] ^ x[46];
  assign t[67] = t[89] ^ x[51];
  assign t[68] = t[90] ^ x[52];
  assign t[69] = t[91] ^ x[57];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[58];
  assign t[71] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[72] = (x[2]);
  assign t[73] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[9]);
  assign t[75] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[12]);
  assign t[77] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[15]);
  assign t[79] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[17] & t[18]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[82] = (x[23]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[86] = (x[37]);
  assign t[87] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[88] = (x[43]);
  assign t[89] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[8] = ~(t[19] & t[20]);
  assign t[90] = (x[49]);
  assign t[91] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[92] = (x[55]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [58:0] x;
 output y;

 wire [92:0] t;
  assign t[0] = t[1] ? t[2] : t[16];
  assign t[10] = ~(t[21] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[19] ? x[27] : x[28];
  assign t[13] = ~(t[22] ^ t[15]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] ^ t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[11];
  assign t[29] = t[40] ^ x[14];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[17];
  assign t[31] = t[42] ^ x[20];
  assign t[32] = t[43] ^ x[26];
  assign t[33] = t[44] ^ x[34];
  assign t[34] = t[45] ^ x[40];
  assign t[35] = t[46] ^ x[46];
  assign t[36] = t[47] ^ x[52];
  assign t[37] = t[48] ^ x[58];
  assign t[38] = (~t[49] & t[50]);
  assign t[39] = (~t[51] & t[52]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[53] & t[54]);
  assign t[41] = (~t[55] & t[56]);
  assign t[42] = (~t[57] & t[58]);
  assign t[43] = (~t[59] & t[60]);
  assign t[44] = (~t[61] & t[62]);
  assign t[45] = (~t[63] & t[64]);
  assign t[46] = (~t[65] & t[66]);
  assign t[47] = (~t[67] & t[68]);
  assign t[48] = (~t[69] & t[70]);
  assign t[49] = t[71] ^ x[4];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[5];
  assign t[51] = t[73] ^ x[10];
  assign t[52] = t[74] ^ x[11];
  assign t[53] = t[75] ^ x[13];
  assign t[54] = t[76] ^ x[14];
  assign t[55] = t[77] ^ x[16];
  assign t[56] = t[78] ^ x[17];
  assign t[57] = t[79] ^ x[19];
  assign t[58] = t[80] ^ x[20];
  assign t[59] = t[81] ^ x[25];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[26];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[39];
  assign t[64] = t[86] ^ x[40];
  assign t[65] = t[87] ^ x[45];
  assign t[66] = t[88] ^ x[46];
  assign t[67] = t[89] ^ x[51];
  assign t[68] = t[90] ^ x[52];
  assign t[69] = t[91] ^ x[57];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[58];
  assign t[71] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[72] = (x[1]);
  assign t[73] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[9]);
  assign t[75] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[12]);
  assign t[77] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[15]);
  assign t[79] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[17] & t[18]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[82] = (x[22]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[86] = (x[36]);
  assign t[87] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[88] = (x[42]);
  assign t[89] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[8] = ~(t[19] & t[20]);
  assign t[90] = (x[48]);
  assign t[91] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[92] = (x[54]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [58:0] x;
 output y;

 wire [127:0] t;
  assign t[0] = t[1] ? t[2] : t[51];
  assign t[100] = t[122] ^ x[45];
  assign t[101] = t[123] ^ x[46];
  assign t[102] = t[124] ^ x[51];
  assign t[103] = t[125] ^ x[52];
  assign t[104] = t[126] ^ x[57];
  assign t[105] = t[127] ^ x[58];
  assign t[106] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[107] = (x[0]);
  assign t[108] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[109] = (x[9]);
  assign t[10] = ~(t[56] ^ t[14]);
  assign t[110] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[111] = (x[12]);
  assign t[112] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[113] = (x[15]);
  assign t[114] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[115] = (x[18]);
  assign t[116] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[117] = (x[21]);
  assign t[118] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[119] = (x[29]);
  assign t[11] = x[27] ^ x[28];
  assign t[120] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[121] = (x[35]);
  assign t[122] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[123] = (x[41]);
  assign t[124] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[125] = (x[47]);
  assign t[126] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[127] = (x[53]);
  assign t[12] = ~(t[57] ^ t[15]);
  assign t[13] = ~(t[16] ^ t[17]);
  assign t[14] = ~(t[58] ^ t[59]);
  assign t[15] = ~(t[60] ^ t[61]);
  assign t[16] = t[18] ? x[27] : x[28];
  assign t[17] = ~(t[19] & t[20]);
  assign t[18] = ~(t[21]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[54]);
  assign t[22] = ~(t[25] & t[26]);
  assign t[23] = ~(t[27] & t[28]);
  assign t[24] = ~(t[29] | t[30]);
  assign t[25] = ~(t[31] & t[32]);
  assign t[26] = ~(t[33] & t[34]);
  assign t[27] = ~(t[35]);
  assign t[28] = t[36] | t[37];
  assign t[29] = ~(t[36]);
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[52] ? t[39] : t[38];
  assign t[31] = ~(t[36] | t[52]);
  assign t[32] = ~(t[40] & t[41]);
  assign t[33] = ~(t[53] | t[42]);
  assign t[34] = t[29] & t[52];
  assign t[35] = ~(t[36] | t[43]);
  assign t[36] = ~(t[54]);
  assign t[37] = t[52] ? t[45] : t[44];
  assign t[38] = ~(t[46] & t[55]);
  assign t[39] = ~(t[47] & t[42]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = ~(t[55] & t[48]);
  assign t[41] = ~(x[7] & t[33]);
  assign t[42] = ~(t[55]);
  assign t[43] = t[52] ? t[44] : t[45];
  assign t[44] = ~(t[48] & t[42]);
  assign t[45] = ~(x[7] & t[49]);
  assign t[46] = x[7] & t[53];
  assign t[47] = ~(x[7] | t[53]);
  assign t[48] = ~(x[7] | t[50]);
  assign t[49] = ~(t[53] | t[55]);
  assign t[4] = ~(x[6]);
  assign t[50] = ~(t[53]);
  assign t[51] = (t[62]);
  assign t[52] = (t[63]);
  assign t[53] = (t[64]);
  assign t[54] = (t[65]);
  assign t[55] = (t[66]);
  assign t[56] = (t[67]);
  assign t[57] = (t[68]);
  assign t[58] = (t[69]);
  assign t[59] = (t[70]);
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = t[73] ^ x[5];
  assign t[63] = t[74] ^ x[11];
  assign t[64] = t[75] ^ x[14];
  assign t[65] = t[76] ^ x[17];
  assign t[66] = t[77] ^ x[20];
  assign t[67] = t[78] ^ x[26];
  assign t[68] = t[79] ^ x[34];
  assign t[69] = t[80] ^ x[40];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[81] ^ x[46];
  assign t[71] = t[82] ^ x[52];
  assign t[72] = t[83] ^ x[58];
  assign t[73] = (~t[84] & t[85]);
  assign t[74] = (~t[86] & t[87]);
  assign t[75] = (~t[88] & t[89]);
  assign t[76] = (~t[90] & t[91]);
  assign t[77] = (~t[92] & t[93]);
  assign t[78] = (~t[94] & t[95]);
  assign t[79] = (~t[96] & t[97]);
  assign t[7] = ~(t[52] & t[53]);
  assign t[80] = (~t[98] & t[99]);
  assign t[81] = (~t[100] & t[101]);
  assign t[82] = (~t[102] & t[103]);
  assign t[83] = (~t[104] & t[105]);
  assign t[84] = t[106] ^ x[4];
  assign t[85] = t[107] ^ x[5];
  assign t[86] = t[108] ^ x[10];
  assign t[87] = t[109] ^ x[11];
  assign t[88] = t[110] ^ x[13];
  assign t[89] = t[111] ^ x[14];
  assign t[8] = ~(t[54] & t[55]);
  assign t[90] = t[112] ^ x[16];
  assign t[91] = t[113] ^ x[17];
  assign t[92] = t[114] ^ x[19];
  assign t[93] = t[115] ^ x[20];
  assign t[94] = t[116] ^ x[25];
  assign t[95] = t[117] ^ x[26];
  assign t[96] = t[118] ^ x[33];
  assign t[97] = t[119] ^ x[34];
  assign t[98] = t[120] ^ x[39];
  assign t[99] = t[121] ^ x[40];
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [88:0] x;
 output y;

 wire [275:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[5];
  assign t[127] = t[159] ^ x[14];
  assign t[128] = t[160] ^ x[22];
  assign t[129] = t[161] ^ x[28];
  assign t[12] = ~(t[96] ^ t[17]);
  assign t[130] = t[162] ^ x[34];
  assign t[131] = t[163] ^ x[37];
  assign t[132] = t[164] ^ x[40];
  assign t[133] = t[165] ^ x[43];
  assign t[134] = t[166] ^ x[46];
  assign t[135] = t[167] ^ x[52];
  assign t[136] = t[168] ^ x[58];
  assign t[137] = t[169] ^ x[59];
  assign t[138] = t[170] ^ x[61];
  assign t[139] = t[171] ^ x[64];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[65];
  assign t[141] = t[173] ^ x[66];
  assign t[142] = t[174] ^ x[67];
  assign t[143] = t[175] ^ x[68];
  assign t[144] = t[176] ^ x[69];
  assign t[145] = t[177] ^ x[71];
  assign t[146] = t[178] ^ x[74];
  assign t[147] = t[179] ^ x[75];
  assign t[148] = t[180] ^ x[76];
  assign t[149] = t[181] ^ x[77];
  assign t[14] = ~(t[97] ^ t[98]);
  assign t[150] = t[182] ^ x[78];
  assign t[151] = t[183] ^ x[79];
  assign t[152] = t[184] ^ x[81];
  assign t[153] = t[185] ^ x[84];
  assign t[154] = t[186] ^ x[85];
  assign t[155] = t[187] ^ x[86];
  assign t[156] = t[188] ^ x[87];
  assign t[157] = t[189] ^ x[88];
  assign t[158] = (~t[190] & t[191]);
  assign t[159] = (~t[192] & t[193]);
  assign t[15] = ~(t[99] & t[100]);
  assign t[160] = (~t[194] & t[195]);
  assign t[161] = (~t[196] & t[197]);
  assign t[162] = (~t[198] & t[199]);
  assign t[163] = (~t[200] & t[201]);
  assign t[164] = (~t[202] & t[203]);
  assign t[165] = (~t[204] & t[205]);
  assign t[166] = (~t[206] & t[207]);
  assign t[167] = (~t[208] & t[209]);
  assign t[168] = (~t[210] & t[211]);
  assign t[169] = (~t[190] & t[212]);
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (~t[192] & t[213]);
  assign t[171] = (~t[194] & t[214]);
  assign t[172] = (~t[198] & t[215]);
  assign t[173] = (~t[196] & t[216]);
  assign t[174] = (~t[210] & t[217]);
  assign t[175] = (~t[208] & t[218]);
  assign t[176] = (~t[190] & t[219]);
  assign t[177] = (~t[192] & t[220]);
  assign t[178] = (~t[194] & t[221]);
  assign t[179] = (~t[196] & t[222]);
  assign t[17] = ~(t[103] ^ t[104]);
  assign t[180] = (~t[198] & t[223]);
  assign t[181] = (~t[208] & t[224]);
  assign t[182] = (~t[210] & t[225]);
  assign t[183] = (~t[190] & t[226]);
  assign t[184] = (~t[192] & t[227]);
  assign t[185] = (~t[194] & t[228]);
  assign t[186] = (~t[196] & t[229]);
  assign t[187] = (~t[198] & t[230]);
  assign t[188] = (~t[208] & t[231]);
  assign t[189] = (~t[210] & t[232]);
  assign t[18] = t[20] ? x[15] : x[16];
  assign t[190] = t[233] ^ x[4];
  assign t[191] = t[234] ^ x[5];
  assign t[192] = t[235] ^ x[13];
  assign t[193] = t[236] ^ x[14];
  assign t[194] = t[237] ^ x[21];
  assign t[195] = t[238] ^ x[22];
  assign t[196] = t[239] ^ x[27];
  assign t[197] = t[240] ^ x[28];
  assign t[198] = t[241] ^ x[33];
  assign t[199] = t[242] ^ x[34];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[36];
  assign t[201] = t[244] ^ x[37];
  assign t[202] = t[245] ^ x[39];
  assign t[203] = t[246] ^ x[40];
  assign t[204] = t[247] ^ x[42];
  assign t[205] = t[248] ^ x[43];
  assign t[206] = t[249] ^ x[45];
  assign t[207] = t[250] ^ x[46];
  assign t[208] = t[251] ^ x[51];
  assign t[209] = t[252] ^ x[52];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[57];
  assign t[211] = t[254] ^ x[58];
  assign t[212] = t[255] ^ x[59];
  assign t[213] = t[256] ^ x[61];
  assign t[214] = t[257] ^ x[64];
  assign t[215] = t[258] ^ x[65];
  assign t[216] = t[259] ^ x[66];
  assign t[217] = t[260] ^ x[67];
  assign t[218] = t[261] ^ x[68];
  assign t[219] = t[262] ^ x[69];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[71];
  assign t[221] = t[264] ^ x[74];
  assign t[222] = t[265] ^ x[75];
  assign t[223] = t[266] ^ x[76];
  assign t[224] = t[267] ^ x[77];
  assign t[225] = t[268] ^ x[78];
  assign t[226] = t[269] ^ x[79];
  assign t[227] = t[270] ^ x[81];
  assign t[228] = t[271] ^ x[84];
  assign t[229] = t[272] ^ x[85];
  assign t[22] = ~(t[26] | t[27]);
  assign t[230] = t[273] ^ x[86];
  assign t[231] = t[274] ^ x[87];
  assign t[232] = t[275] ^ x[88];
  assign t[233] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[234] = (x[0]);
  assign t[235] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[236] = (x[9]);
  assign t[237] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[238] = (x[17]);
  assign t[239] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[23] = ~(t[101]);
  assign t[240] = (x[23]);
  assign t[241] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[242] = (x[29]);
  assign t[243] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[244] = (x[35]);
  assign t[245] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[246] = (x[38]);
  assign t[247] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[248] = (x[41]);
  assign t[249] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[24] = ~(t[28] & t[29]);
  assign t[250] = (x[44]);
  assign t[251] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[252] = (x[47]);
  assign t[253] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[254] = (x[53]);
  assign t[255] = (x[1]);
  assign t[256] = (x[10]);
  assign t[257] = (x[18]);
  assign t[258] = (x[30]);
  assign t[259] = (x[24]);
  assign t[25] = ~(t[30] & t[31]);
  assign t[260] = (x[54]);
  assign t[261] = (x[48]);
  assign t[262] = (x[2]);
  assign t[263] = (x[11]);
  assign t[264] = (x[19]);
  assign t[265] = (x[25]);
  assign t[266] = (x[31]);
  assign t[267] = (x[49]);
  assign t[268] = (x[55]);
  assign t[269] = (x[3]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[270] = (x[12]);
  assign t[271] = (x[20]);
  assign t[272] = (x[26]);
  assign t[273] = (x[32]);
  assign t[274] = (x[50]);
  assign t[275] = (x[56]);
  assign t[27] = ~(t[32] | t[34]);
  assign t[28] = ~(t[35] | t[36]);
  assign t[29] = ~(t[37] & t[38]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[39] & t[40]);
  assign t[31] = t[37] | t[41];
  assign t[32] = ~(t[37]);
  assign t[33] = t[99] ? t[43] : t[42];
  assign t[34] = t[99] ? t[45] : t[44];
  assign t[35] = ~(t[37] | t[46]);
  assign t[36] = ~(t[32] | t[47]);
  assign t[37] = ~(t[101]);
  assign t[38] = ~(t[48] & t[49]);
  assign t[39] = t[102] & t[50];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] | t[52];
  assign t[41] = t[99] ? t[48] : t[53];
  assign t[42] = ~(t[51] & t[54]);
  assign t[43] = ~(t[52] & t[102]);
  assign t[44] = ~(t[51] & t[102]);
  assign t[45] = ~(t[52] & t[54]);
  assign t[46] = t[99] ? t[42] : t[45];
  assign t[47] = t[99] ? t[53] : t[55];
  assign t[48] = ~(x[7] & t[56]);
  assign t[49] = ~(t[102] & t[57]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[37] | t[99]);
  assign t[51] = ~(x[7] | t[100]);
  assign t[52] = x[7] & t[100];
  assign t[53] = ~(t[57] & t[54]);
  assign t[54] = ~(t[102]);
  assign t[55] = ~(x[7] & t[58]);
  assign t[56] = ~(t[100] | t[102]);
  assign t[57] = ~(x[7] | t[59]);
  assign t[58] = ~(t[100] | t[54]);
  assign t[59] = ~(t[100]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[1] ? t[61] : t[105];
  assign t[61] = x[6] ? t[63] : t[62];
  assign t[62] = x[7] ? t[65] : t[64];
  assign t[63] = t[66] ^ x[60];
  assign t[64] = t[67] ^ t[68];
  assign t[65] = ~(t[106] ^ t[69]);
  assign t[66] = x[62] ^ x[63];
  assign t[67] = t[70] ? x[62] : x[63];
  assign t[68] = ~(t[107] ^ t[71]);
  assign t[69] = ~(t[108] ^ t[109]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[23]);
  assign t[71] = ~(t[110] ^ t[111]);
  assign t[72] = t[1] ? t[73] : t[112];
  assign t[73] = x[6] ? t[75] : t[74];
  assign t[74] = x[7] ? t[77] : t[76];
  assign t[75] = t[78] ^ x[70];
  assign t[76] = t[79] ^ t[80];
  assign t[77] = ~(t[113] ^ t[81]);
  assign t[78] = x[72] ^ x[73];
  assign t[79] = t[20] ? x[72] : x[73];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[114] ^ t[82]);
  assign t[81] = ~(t[115] ^ t[116]);
  assign t[82] = ~(t[117] ^ t[118]);
  assign t[83] = t[1] ? t[84] : t[119];
  assign t[84] = x[6] ? t[86] : t[85];
  assign t[85] = x[7] ? t[88] : t[87];
  assign t[86] = t[89] ^ x[80];
  assign t[87] = t[90] ^ t[91];
  assign t[88] = ~(t[120] ^ t[92]);
  assign t[89] = x[82] ^ x[83];
  assign t[8] = ~(t[95] ^ t[14]);
  assign t[90] = t[20] ? x[82] : x[83];
  assign t[91] = ~(t[121] ^ t[93]);
  assign t[92] = ~(t[122] ^ t[123]);
  assign t[93] = ~(t[124] ^ t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[60] & ~t[72] & ~t[83]) | (~t[0] & t[60] & ~t[72] & ~t[83]) | (~t[0] & ~t[60] & t[72] & ~t[83]) | (~t[0] & ~t[60] & ~t[72] & t[83]) | (t[0] & t[60] & t[72] & ~t[83]) | (t[0] & t[60] & ~t[72] & t[83]) | (t[0] & ~t[60] & t[72] & t[83]) | (~t[0] & t[60] & t[72] & t[83]);
endmodule

module R2ind131(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[2]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[11]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[19]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[25]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[49]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[1]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[10]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[18]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[48]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[54]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [58:0] x;
 output y;

 wire [136:0] t;
  assign t[0] = t[1] ? t[2] : t[60];
  assign t[100] = t[122] ^ x[28];
  assign t[101] = t[123] ^ x[33];
  assign t[102] = t[124] ^ x[34];
  assign t[103] = t[125] ^ x[36];
  assign t[104] = t[126] ^ x[37];
  assign t[105] = t[127] ^ x[39];
  assign t[106] = t[128] ^ x[40];
  assign t[107] = t[129] ^ x[42];
  assign t[108] = t[130] ^ x[43];
  assign t[109] = t[131] ^ x[45];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[132] ^ x[46];
  assign t[111] = t[133] ^ x[51];
  assign t[112] = t[134] ^ x[52];
  assign t[113] = t[135] ^ x[57];
  assign t[114] = t[136] ^ x[58];
  assign t[115] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[116] = (x[0]);
  assign t[117] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[118] = (x[9]);
  assign t[119] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[17]);
  assign t[121] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[122] = (x[23]);
  assign t[123] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[124] = (x[29]);
  assign t[125] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[35]);
  assign t[127] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[38]);
  assign t[129] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[62] ^ t[17]);
  assign t[130] = (x[41]);
  assign t[131] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[132] = (x[44]);
  assign t[133] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[134] = (x[47]);
  assign t[135] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[136] = (x[53]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[63] ^ t[64]);
  assign t[15] = ~(t[65] & t[66]);
  assign t[16] = ~(t[67] & t[68]);
  assign t[17] = ~(t[69] ^ t[70]);
  assign t[18] = t[20] ? x[15] : x[16];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[67]);
  assign t[24] = ~(t[28] & t[29]);
  assign t[25] = ~(t[30] & t[31]);
  assign t[26] = ~(t[32] | t[33]);
  assign t[27] = ~(t[32] | t[34]);
  assign t[28] = ~(t[35] | t[36]);
  assign t[29] = ~(t[37] & t[38]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[39] & t[40]);
  assign t[31] = t[37] | t[41];
  assign t[32] = ~(t[37]);
  assign t[33] = t[65] ? t[43] : t[42];
  assign t[34] = t[65] ? t[45] : t[44];
  assign t[35] = ~(t[37] | t[46]);
  assign t[36] = ~(t[32] | t[47]);
  assign t[37] = ~(t[67]);
  assign t[38] = ~(t[48] & t[49]);
  assign t[39] = t[68] & t[50];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] | t[52];
  assign t[41] = t[65] ? t[48] : t[53];
  assign t[42] = ~(t[51] & t[54]);
  assign t[43] = ~(t[52] & t[68]);
  assign t[44] = ~(t[51] & t[68]);
  assign t[45] = ~(t[52] & t[54]);
  assign t[46] = t[65] ? t[42] : t[45];
  assign t[47] = t[65] ? t[53] : t[55];
  assign t[48] = ~(x[7] & t[56]);
  assign t[49] = ~(t[68] & t[57]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[37] | t[65]);
  assign t[51] = ~(x[7] | t[66]);
  assign t[52] = x[7] & t[66];
  assign t[53] = ~(t[57] & t[54]);
  assign t[54] = ~(t[68]);
  assign t[55] = ~(x[7] & t[58]);
  assign t[56] = ~(t[66] | t[68]);
  assign t[57] = ~(x[7] | t[59]);
  assign t[58] = ~(t[66] | t[54]);
  assign t[59] = ~(t[66]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = (t[73]);
  assign t[63] = (t[74]);
  assign t[64] = (t[75]);
  assign t[65] = (t[76]);
  assign t[66] = (t[77]);
  assign t[67] = (t[78]);
  assign t[68] = (t[79]);
  assign t[69] = (t[80]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[81]);
  assign t[71] = t[82] ^ x[5];
  assign t[72] = t[83] ^ x[14];
  assign t[73] = t[84] ^ x[22];
  assign t[74] = t[85] ^ x[28];
  assign t[75] = t[86] ^ x[34];
  assign t[76] = t[87] ^ x[37];
  assign t[77] = t[88] ^ x[40];
  assign t[78] = t[89] ^ x[43];
  assign t[79] = t[90] ^ x[46];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[91] ^ x[52];
  assign t[81] = t[92] ^ x[58];
  assign t[82] = (~t[93] & t[94]);
  assign t[83] = (~t[95] & t[96]);
  assign t[84] = (~t[97] & t[98]);
  assign t[85] = (~t[99] & t[100]);
  assign t[86] = (~t[101] & t[102]);
  assign t[87] = (~t[103] & t[104]);
  assign t[88] = (~t[105] & t[106]);
  assign t[89] = (~t[107] & t[108]);
  assign t[8] = ~(t[61] ^ t[14]);
  assign t[90] = (~t[109] & t[110]);
  assign t[91] = (~t[111] & t[112]);
  assign t[92] = (~t[113] & t[114]);
  assign t[93] = t[115] ^ x[4];
  assign t[94] = t[116] ^ x[5];
  assign t[95] = t[117] ^ x[13];
  assign t[96] = t[118] ^ x[14];
  assign t[97] = t[119] ^ x[21];
  assign t[98] = t[120] ^ x[22];
  assign t[99] = t[121] ^ x[27];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [88:0] x;
 output y;

 wire [270:0] t;
  assign t[0] = t[1] ? t[2] : t[89];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = t[153] ^ x[5];
  assign t[122] = t[154] ^ x[14];
  assign t[123] = t[155] ^ x[22];
  assign t[124] = t[156] ^ x[28];
  assign t[125] = t[157] ^ x[34];
  assign t[126] = t[158] ^ x[37];
  assign t[127] = t[159] ^ x[40];
  assign t[128] = t[160] ^ x[43];
  assign t[129] = t[161] ^ x[46];
  assign t[12] = ~(t[91] ^ t[17]);
  assign t[130] = t[162] ^ x[52];
  assign t[131] = t[163] ^ x[58];
  assign t[132] = t[164] ^ x[59];
  assign t[133] = t[165] ^ x[61];
  assign t[134] = t[166] ^ x[64];
  assign t[135] = t[167] ^ x[65];
  assign t[136] = t[168] ^ x[66];
  assign t[137] = t[169] ^ x[67];
  assign t[138] = t[170] ^ x[68];
  assign t[139] = t[171] ^ x[69];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[71];
  assign t[141] = t[173] ^ x[74];
  assign t[142] = t[174] ^ x[75];
  assign t[143] = t[175] ^ x[76];
  assign t[144] = t[176] ^ x[77];
  assign t[145] = t[177] ^ x[78];
  assign t[146] = t[178] ^ x[79];
  assign t[147] = t[179] ^ x[81];
  assign t[148] = t[180] ^ x[84];
  assign t[149] = t[181] ^ x[85];
  assign t[14] = ~(t[92] ^ t[93]);
  assign t[150] = t[182] ^ x[86];
  assign t[151] = t[183] ^ x[87];
  assign t[152] = t[184] ^ x[88];
  assign t[153] = (~t[185] & t[186]);
  assign t[154] = (~t[187] & t[188]);
  assign t[155] = (~t[189] & t[190]);
  assign t[156] = (~t[191] & t[192]);
  assign t[157] = (~t[193] & t[194]);
  assign t[158] = (~t[195] & t[196]);
  assign t[159] = (~t[197] & t[198]);
  assign t[15] = ~(t[94] & t[95]);
  assign t[160] = (~t[199] & t[200]);
  assign t[161] = (~t[201] & t[202]);
  assign t[162] = (~t[203] & t[204]);
  assign t[163] = (~t[205] & t[206]);
  assign t[164] = (~t[185] & t[207]);
  assign t[165] = (~t[187] & t[208]);
  assign t[166] = (~t[189] & t[209]);
  assign t[167] = (~t[193] & t[210]);
  assign t[168] = (~t[191] & t[211]);
  assign t[169] = (~t[205] & t[212]);
  assign t[16] = ~(t[96] & t[97]);
  assign t[170] = (~t[203] & t[213]);
  assign t[171] = (~t[185] & t[214]);
  assign t[172] = (~t[187] & t[215]);
  assign t[173] = (~t[189] & t[216]);
  assign t[174] = (~t[193] & t[217]);
  assign t[175] = (~t[191] & t[218]);
  assign t[176] = (~t[203] & t[219]);
  assign t[177] = (~t[205] & t[220]);
  assign t[178] = (~t[185] & t[221]);
  assign t[179] = (~t[187] & t[222]);
  assign t[17] = ~(t[98] ^ t[99]);
  assign t[180] = (~t[189] & t[223]);
  assign t[181] = (~t[193] & t[224]);
  assign t[182] = (~t[191] & t[225]);
  assign t[183] = (~t[203] & t[226]);
  assign t[184] = (~t[205] & t[227]);
  assign t[185] = t[228] ^ x[4];
  assign t[186] = t[229] ^ x[5];
  assign t[187] = t[230] ^ x[13];
  assign t[188] = t[231] ^ x[14];
  assign t[189] = t[232] ^ x[21];
  assign t[18] = t[20] ? x[15] : x[16];
  assign t[190] = t[233] ^ x[22];
  assign t[191] = t[234] ^ x[27];
  assign t[192] = t[235] ^ x[28];
  assign t[193] = t[236] ^ x[33];
  assign t[194] = t[237] ^ x[34];
  assign t[195] = t[238] ^ x[36];
  assign t[196] = t[239] ^ x[37];
  assign t[197] = t[240] ^ x[39];
  assign t[198] = t[241] ^ x[40];
  assign t[199] = t[242] ^ x[42];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[43];
  assign t[201] = t[244] ^ x[45];
  assign t[202] = t[245] ^ x[46];
  assign t[203] = t[246] ^ x[51];
  assign t[204] = t[247] ^ x[52];
  assign t[205] = t[248] ^ x[57];
  assign t[206] = t[249] ^ x[58];
  assign t[207] = t[250] ^ x[59];
  assign t[208] = t[251] ^ x[61];
  assign t[209] = t[252] ^ x[64];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[65];
  assign t[211] = t[254] ^ x[66];
  assign t[212] = t[255] ^ x[67];
  assign t[213] = t[256] ^ x[68];
  assign t[214] = t[257] ^ x[69];
  assign t[215] = t[258] ^ x[71];
  assign t[216] = t[259] ^ x[74];
  assign t[217] = t[260] ^ x[75];
  assign t[218] = t[261] ^ x[76];
  assign t[219] = t[262] ^ x[77];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[78];
  assign t[221] = t[264] ^ x[79];
  assign t[222] = t[265] ^ x[81];
  assign t[223] = t[266] ^ x[84];
  assign t[224] = t[267] ^ x[85];
  assign t[225] = t[268] ^ x[86];
  assign t[226] = t[269] ^ x[87];
  assign t[227] = t[270] ^ x[88];
  assign t[228] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[229] = (x[0]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[230] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[231] = (x[9]);
  assign t[232] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[233] = (x[17]);
  assign t[234] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[235] = (x[23]);
  assign t[236] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[237] = (x[29]);
  assign t[238] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[239] = (x[35]);
  assign t[23] = ~(t[96]);
  assign t[240] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[241] = (x[38]);
  assign t[242] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[243] = (x[41]);
  assign t[244] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[245] = (x[44]);
  assign t[246] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[247] = (x[47]);
  assign t[248] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[249] = (x[53]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[250] = (x[1]);
  assign t[251] = (x[10]);
  assign t[252] = (x[18]);
  assign t[253] = (x[30]);
  assign t[254] = (x[24]);
  assign t[255] = (x[54]);
  assign t[256] = (x[48]);
  assign t[257] = (x[2]);
  assign t[258] = (x[11]);
  assign t[259] = (x[19]);
  assign t[25] = ~(t[30] | t[31]);
  assign t[260] = (x[31]);
  assign t[261] = (x[25]);
  assign t[262] = (x[49]);
  assign t[263] = (x[55]);
  assign t[264] = (x[3]);
  assign t[265] = (x[12]);
  assign t[266] = (x[20]);
  assign t[267] = (x[32]);
  assign t[268] = (x[26]);
  assign t[269] = (x[50]);
  assign t[26] = ~(t[30] | t[32]);
  assign t[270] = (x[56]);
  assign t[27] = ~(t[33] & t[34]);
  assign t[28] = ~(t[96]);
  assign t[29] = t[94] ? t[36] : t[35];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[28]);
  assign t[31] = t[94] ? t[38] : t[37];
  assign t[32] = t[94] ? t[39] : t[35];
  assign t[33] = ~(t[40] | t[41]);
  assign t[34] = t[28] | t[42];
  assign t[35] = ~(t[43] & t[44]);
  assign t[36] = ~(t[45] & t[44]);
  assign t[37] = ~(x[7] & t[46]);
  assign t[38] = ~(t[47] & t[44]);
  assign t[39] = ~(t[45] & t[97]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[30] | t[48]);
  assign t[41] = ~(t[30] | t[49]);
  assign t[42] = t[94] ? t[50] : t[38];
  assign t[43] = x[7] & t[95];
  assign t[44] = ~(t[97]);
  assign t[45] = ~(x[7] | t[95]);
  assign t[46] = ~(t[95] | t[44]);
  assign t[47] = ~(x[7] | t[51]);
  assign t[48] = t[94] ? t[52] : t[36];
  assign t[49] = t[94] ? t[35] : t[39];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(x[7] & t[53]);
  assign t[51] = ~(t[95]);
  assign t[52] = ~(t[43] & t[97]);
  assign t[53] = ~(t[95] | t[97]);
  assign t[54] = t[1] ? t[55] : t[100];
  assign t[55] = x[6] ? t[57] : t[56];
  assign t[56] = x[7] ? t[59] : t[58];
  assign t[57] = t[60] ^ x[60];
  assign t[58] = t[61] ^ t[62];
  assign t[59] = ~(t[101] ^ t[63]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = x[62] ^ x[63];
  assign t[61] = t[20] ? x[62] : x[63];
  assign t[62] = ~(t[102] ^ t[64]);
  assign t[63] = ~(t[103] ^ t[104]);
  assign t[64] = ~(t[105] ^ t[106]);
  assign t[65] = t[1] ? t[66] : t[107];
  assign t[66] = x[6] ? t[68] : t[67];
  assign t[67] = x[7] ? t[70] : t[69];
  assign t[68] = t[71] ^ x[70];
  assign t[69] = t[72] ^ t[73];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] ^ t[74]);
  assign t[71] = x[72] ^ x[73];
  assign t[72] = t[75] ? x[72] : x[73];
  assign t[73] = ~(t[109] ^ t[76]);
  assign t[74] = ~(t[110] ^ t[111]);
  assign t[75] = ~(t[23]);
  assign t[76] = ~(t[112] ^ t[113]);
  assign t[77] = t[1] ? t[78] : t[114];
  assign t[78] = x[6] ? t[80] : t[79];
  assign t[79] = x[7] ? t[82] : t[81];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[83] ^ x[80];
  assign t[81] = t[84] ^ t[85];
  assign t[82] = ~(t[115] ^ t[86]);
  assign t[83] = x[82] ^ x[83];
  assign t[84] = t[87] ? x[82] : x[83];
  assign t[85] = ~(t[116] ^ t[88]);
  assign t[86] = ~(t[117] ^ t[118]);
  assign t[87] = ~(t[23]);
  assign t[88] = ~(t[119] ^ t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[90] ^ t[14]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[54] & ~t[65] & ~t[77]) | (~t[0] & t[54] & ~t[65] & ~t[77]) | (~t[0] & ~t[54] & t[65] & ~t[77]) | (~t[0] & ~t[54] & ~t[65] & t[77]) | (t[0] & t[54] & t[65] & ~t[77]) | (t[0] & t[54] & ~t[65] & t[77]) | (t[0] & ~t[54] & t[65] & t[77]) | (~t[0] & t[54] & t[65] & t[77]);
endmodule

module R2ind136(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[2]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[11]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[19]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[25]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[49]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[1]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[10]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[18]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[48]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[54]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [58:0] x;
 output y;

 wire [130:0] t;
  assign t[0] = t[1] ? t[2] : t[54];
  assign t[100] = t[122] ^ x[40];
  assign t[101] = t[123] ^ x[42];
  assign t[102] = t[124] ^ x[43];
  assign t[103] = t[125] ^ x[45];
  assign t[104] = t[126] ^ x[46];
  assign t[105] = t[127] ^ x[51];
  assign t[106] = t[128] ^ x[52];
  assign t[107] = t[129] ^ x[57];
  assign t[108] = t[130] ^ x[58];
  assign t[109] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (x[0]);
  assign t[111] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[112] = (x[9]);
  assign t[113] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[114] = (x[17]);
  assign t[115] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[116] = (x[23]);
  assign t[117] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[118] = (x[29]);
  assign t[119] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[35]);
  assign t[121] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[38]);
  assign t[123] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[41]);
  assign t[125] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[44]);
  assign t[127] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[128] = (x[47]);
  assign t[129] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[12] = ~(t[56] ^ t[17]);
  assign t[130] = (x[53]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[57] ^ t[58]);
  assign t[15] = ~(t[59] & t[60]);
  assign t[16] = ~(t[61] & t[62]);
  assign t[17] = ~(t[63] ^ t[64]);
  assign t[18] = t[20] ? x[15] : x[16];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[61]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[25] = ~(t[30] | t[31]);
  assign t[26] = ~(t[30] | t[32]);
  assign t[27] = ~(t[33] & t[34]);
  assign t[28] = ~(t[61]);
  assign t[29] = t[59] ? t[36] : t[35];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[28]);
  assign t[31] = t[59] ? t[38] : t[37];
  assign t[32] = t[59] ? t[39] : t[35];
  assign t[33] = ~(t[40] | t[41]);
  assign t[34] = t[28] | t[42];
  assign t[35] = ~(t[43] & t[44]);
  assign t[36] = ~(t[45] & t[44]);
  assign t[37] = ~(x[7] & t[46]);
  assign t[38] = ~(t[47] & t[44]);
  assign t[39] = ~(t[45] & t[62]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[30] | t[48]);
  assign t[41] = ~(t[30] | t[49]);
  assign t[42] = t[59] ? t[50] : t[38];
  assign t[43] = x[7] & t[60];
  assign t[44] = ~(t[62]);
  assign t[45] = ~(x[7] | t[60]);
  assign t[46] = ~(t[60] | t[44]);
  assign t[47] = ~(x[7] | t[51]);
  assign t[48] = t[59] ? t[52] : t[36];
  assign t[49] = t[59] ? t[35] : t[39];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(x[7] & t[53]);
  assign t[51] = ~(t[60]);
  assign t[52] = ~(t[43] & t[62]);
  assign t[53] = ~(t[60] | t[62]);
  assign t[54] = (t[65]);
  assign t[55] = (t[66]);
  assign t[56] = (t[67]);
  assign t[57] = (t[68]);
  assign t[58] = (t[69]);
  assign t[59] = (t[70]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = (t[73]);
  assign t[63] = (t[74]);
  assign t[64] = (t[75]);
  assign t[65] = t[76] ^ x[5];
  assign t[66] = t[77] ^ x[14];
  assign t[67] = t[78] ^ x[22];
  assign t[68] = t[79] ^ x[28];
  assign t[69] = t[80] ^ x[34];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[81] ^ x[37];
  assign t[71] = t[82] ^ x[40];
  assign t[72] = t[83] ^ x[43];
  assign t[73] = t[84] ^ x[46];
  assign t[74] = t[85] ^ x[52];
  assign t[75] = t[86] ^ x[58];
  assign t[76] = (~t[87] & t[88]);
  assign t[77] = (~t[89] & t[90]);
  assign t[78] = (~t[91] & t[92]);
  assign t[79] = (~t[93] & t[94]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[95] & t[96]);
  assign t[81] = (~t[97] & t[98]);
  assign t[82] = (~t[99] & t[100]);
  assign t[83] = (~t[101] & t[102]);
  assign t[84] = (~t[103] & t[104]);
  assign t[85] = (~t[105] & t[106]);
  assign t[86] = (~t[107] & t[108]);
  assign t[87] = t[109] ^ x[4];
  assign t[88] = t[110] ^ x[5];
  assign t[89] = t[111] ^ x[13];
  assign t[8] = ~(t[55] ^ t[14]);
  assign t[90] = t[112] ^ x[14];
  assign t[91] = t[113] ^ x[21];
  assign t[92] = t[114] ^ x[22];
  assign t[93] = t[115] ^ x[27];
  assign t[94] = t[116] ^ x[28];
  assign t[95] = t[117] ^ x[33];
  assign t[96] = t[118] ^ x[34];
  assign t[97] = t[119] ^ x[36];
  assign t[98] = t[120] ^ x[37];
  assign t[99] = t[121] ^ x[39];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [70:0] x;
 output y;

 wire [220:0] t;
  assign t[0] = t[1] ? t[2] : t[83];
  assign t[100] = (t[124]);
  assign t[101] = (t[125]);
  assign t[102] = (t[126]);
  assign t[103] = (t[127]);
  assign t[104] = (t[128]);
  assign t[105] = (t[129]);
  assign t[106] = (t[130]);
  assign t[107] = t[131] ^ x[5];
  assign t[108] = t[132] ^ x[14];
  assign t[109] = t[133] ^ x[22];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[134] ^ x[28];
  assign t[111] = t[135] ^ x[34];
  assign t[112] = t[136] ^ x[37];
  assign t[113] = t[137] ^ x[40];
  assign t[114] = t[138] ^ x[43];
  assign t[115] = t[139] ^ x[46];
  assign t[116] = t[140] ^ x[47];
  assign t[117] = t[141] ^ x[49];
  assign t[118] = t[142] ^ x[52];
  assign t[119] = t[143] ^ x[53];
  assign t[11] = ~(x[6]);
  assign t[120] = t[144] ^ x[54];
  assign t[121] = t[145] ^ x[55];
  assign t[122] = t[146] ^ x[57];
  assign t[123] = t[147] ^ x[60];
  assign t[124] = t[148] ^ x[61];
  assign t[125] = t[149] ^ x[62];
  assign t[126] = t[150] ^ x[63];
  assign t[127] = t[151] ^ x[65];
  assign t[128] = t[152] ^ x[68];
  assign t[129] = t[153] ^ x[69];
  assign t[12] = ~(t[85] ^ t[14]);
  assign t[130] = t[154] ^ x[70];
  assign t[131] = (~t[155] & t[156]);
  assign t[132] = (~t[157] & t[158]);
  assign t[133] = (~t[159] & t[160]);
  assign t[134] = (~t[161] & t[162]);
  assign t[135] = (~t[163] & t[164]);
  assign t[136] = (~t[165] & t[166]);
  assign t[137] = (~t[167] & t[168]);
  assign t[138] = (~t[169] & t[170]);
  assign t[139] = (~t[171] & t[172]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (~t[155] & t[173]);
  assign t[141] = (~t[157] & t[174]);
  assign t[142] = (~t[159] & t[175]);
  assign t[143] = (~t[163] & t[176]);
  assign t[144] = (~t[161] & t[177]);
  assign t[145] = (~t[155] & t[178]);
  assign t[146] = (~t[157] & t[179]);
  assign t[147] = (~t[159] & t[180]);
  assign t[148] = (~t[163] & t[181]);
  assign t[149] = (~t[161] & t[182]);
  assign t[14] = ~(t[86] ^ t[87]);
  assign t[150] = (~t[155] & t[183]);
  assign t[151] = (~t[157] & t[184]);
  assign t[152] = (~t[159] & t[185]);
  assign t[153] = (~t[163] & t[186]);
  assign t[154] = (~t[161] & t[187]);
  assign t[155] = t[188] ^ x[4];
  assign t[156] = t[189] ^ x[5];
  assign t[157] = t[190] ^ x[13];
  assign t[158] = t[191] ^ x[14];
  assign t[159] = t[192] ^ x[21];
  assign t[15] = ~(t[88] & t[89]);
  assign t[160] = t[193] ^ x[22];
  assign t[161] = t[194] ^ x[27];
  assign t[162] = t[195] ^ x[28];
  assign t[163] = t[196] ^ x[33];
  assign t[164] = t[197] ^ x[34];
  assign t[165] = t[198] ^ x[36];
  assign t[166] = t[199] ^ x[37];
  assign t[167] = t[200] ^ x[39];
  assign t[168] = t[201] ^ x[40];
  assign t[169] = t[202] ^ x[42];
  assign t[16] = ~(t[90] & t[91]);
  assign t[170] = t[203] ^ x[43];
  assign t[171] = t[204] ^ x[45];
  assign t[172] = t[205] ^ x[46];
  assign t[173] = t[206] ^ x[47];
  assign t[174] = t[207] ^ x[49];
  assign t[175] = t[208] ^ x[52];
  assign t[176] = t[209] ^ x[53];
  assign t[177] = t[210] ^ x[54];
  assign t[178] = t[211] ^ x[55];
  assign t[179] = t[212] ^ x[57];
  assign t[17] = t[19] ? x[15] : x[16];
  assign t[180] = t[213] ^ x[60];
  assign t[181] = t[214] ^ x[61];
  assign t[182] = t[215] ^ x[62];
  assign t[183] = t[216] ^ x[63];
  assign t[184] = t[217] ^ x[65];
  assign t[185] = t[218] ^ x[68];
  assign t[186] = t[219] ^ x[69];
  assign t[187] = t[220] ^ x[70];
  assign t[188] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[189] = (x[0]);
  assign t[18] = ~(t[20] & t[21]);
  assign t[190] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[191] = (x[9]);
  assign t[192] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[193] = (x[17]);
  assign t[194] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[195] = (x[23]);
  assign t[196] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[197] = (x[29]);
  assign t[198] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[199] = (x[35]);
  assign t[19] = ~(t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[201] = (x[38]);
  assign t[202] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[203] = (x[41]);
  assign t[204] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[205] = (x[44]);
  assign t[206] = (x[1]);
  assign t[207] = (x[10]);
  assign t[208] = (x[18]);
  assign t[209] = (x[30]);
  assign t[20] = ~(t[23] | t[24]);
  assign t[210] = (x[24]);
  assign t[211] = (x[2]);
  assign t[212] = (x[11]);
  assign t[213] = (x[19]);
  assign t[214] = (x[31]);
  assign t[215] = (x[25]);
  assign t[216] = (x[3]);
  assign t[217] = (x[12]);
  assign t[218] = (x[20]);
  assign t[219] = (x[32]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[220] = (x[26]);
  assign t[22] = ~(t[90]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[27] | t[29]);
  assign t[25] = ~(t[30] | t[31]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[30]);
  assign t[28] = t[88] ? t[35] : t[34];
  assign t[29] = t[88] ? t[37] : t[36];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[90]);
  assign t[31] = t[88] ? t[35] : t[36];
  assign t[32] = ~(t[38] | t[39]);
  assign t[33] = ~(t[40] & t[41]);
  assign t[34] = ~(t[42] & t[91]);
  assign t[35] = ~(t[43] & t[44]);
  assign t[36] = ~(t[42] & t[44]);
  assign t[37] = ~(t[43] & t[91]);
  assign t[38] = ~(t[30] | t[45]);
  assign t[39] = ~(t[30] | t[46]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[89] | t[44]);
  assign t[41] = t[27] & t[88];
  assign t[42] = x[7] & t[89];
  assign t[43] = ~(x[7] | t[89]);
  assign t[44] = ~(t[91]);
  assign t[45] = t[88] ? t[36] : t[35];
  assign t[46] = t[88] ? t[48] : t[47];
  assign t[47] = ~(x[7] & t[49]);
  assign t[48] = ~(t[50] & t[44]);
  assign t[49] = ~(t[89] | t[91]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(x[7] | t[51]);
  assign t[51] = ~(t[89]);
  assign t[52] = t[1] ? t[53] : t[92];
  assign t[53] = x[6] ? t[55] : t[54];
  assign t[54] = x[7] ? t[57] : t[56];
  assign t[55] = t[58] ^ x[48];
  assign t[56] = t[59] ^ t[60];
  assign t[57] = ~(t[93] ^ t[61]);
  assign t[58] = x[50] ^ x[51];
  assign t[59] = t[62] ? x[50] : x[51];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[94] ^ t[61]);
  assign t[61] = ~(t[95] ^ t[96]);
  assign t[62] = ~(t[22]);
  assign t[63] = t[1] ? t[64] : t[97];
  assign t[64] = x[6] ? t[66] : t[65];
  assign t[65] = x[7] ? t[68] : t[67];
  assign t[66] = t[69] ^ x[56];
  assign t[67] = t[70] ^ t[71];
  assign t[68] = ~(t[98] ^ t[72]);
  assign t[69] = x[58] ^ x[59];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[90] ? x[58] : x[59];
  assign t[71] = ~(t[99] ^ t[72]);
  assign t[72] = ~(t[100] ^ t[101]);
  assign t[73] = t[1] ? t[74] : t[102];
  assign t[74] = x[6] ? t[76] : t[75];
  assign t[75] = x[7] ? t[78] : t[77];
  assign t[76] = t[79] ^ x[64];
  assign t[77] = t[80] ^ t[81];
  assign t[78] = ~(t[103] ^ t[82]);
  assign t[79] = x[66] ^ x[67];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[19] ? x[66] : x[67];
  assign t[81] = ~(t[104] ^ t[82]);
  assign t[82] = ~(t[105] ^ t[106]);
  assign t[83] = (t[107]);
  assign t[84] = (t[108]);
  assign t[85] = (t[109]);
  assign t[86] = (t[110]);
  assign t[87] = (t[111]);
  assign t[88] = (t[112]);
  assign t[89] = (t[113]);
  assign t[8] = ~(t[84] ^ t[14]);
  assign t[90] = (t[114]);
  assign t[91] = (t[115]);
  assign t[92] = (t[116]);
  assign t[93] = (t[117]);
  assign t[94] = (t[118]);
  assign t[95] = (t[119]);
  assign t[96] = (t[120]);
  assign t[97] = (t[121]);
  assign t[98] = (t[122]);
  assign t[99] = (t[123]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[52] & ~t[63] & ~t[73]) | (~t[0] & t[52] & ~t[63] & ~t[73]) | (~t[0] & ~t[52] & t[63] & ~t[73]) | (~t[0] & ~t[52] & ~t[63] & t[73]) | (t[0] & t[52] & t[63] & ~t[73]) | (t[0] & t[52] & ~t[63] & t[73]) | (t[0] & ~t[52] & t[63] & t[73]) | (~t[0] & t[52] & t[63] & t[73]);
endmodule

module R2ind141(x, y);
 input [46:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = t[1] ? t[2] : t[19];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[21] ^ t[14]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[26] & t[27]);
  assign t[17] = ~(t[18]);
  assign t[18] = ~(t[26]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = t[37] ^ x[5];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[39] ^ x[22];
  assign t[31] = t[40] ^ x[28];
  assign t[32] = t[41] ^ x[34];
  assign t[33] = t[42] ^ x[37];
  assign t[34] = t[43] ^ x[40];
  assign t[35] = t[44] ^ x[43];
  assign t[36] = t[45] ^ x[46];
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[48] & t[49]);
  assign t[39] = (~t[50] & t[51]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[52] & t[53]);
  assign t[41] = (~t[54] & t[55]);
  assign t[42] = (~t[56] & t[57]);
  assign t[43] = (~t[58] & t[59]);
  assign t[44] = (~t[60] & t[61]);
  assign t[45] = (~t[62] & t[63]);
  assign t[46] = t[64] ^ x[4];
  assign t[47] = t[65] ^ x[5];
  assign t[48] = t[66] ^ x[13];
  assign t[49] = t[67] ^ x[14];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[68] ^ x[21];
  assign t[51] = t[69] ^ x[22];
  assign t[52] = t[70] ^ x[27];
  assign t[53] = t[71] ^ x[28];
  assign t[54] = t[72] ^ x[33];
  assign t[55] = t[73] ^ x[34];
  assign t[56] = t[74] ^ x[36];
  assign t[57] = t[75] ^ x[37];
  assign t[58] = t[76] ^ x[39];
  assign t[59] = t[77] ^ x[40];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[78] ^ x[42];
  assign t[61] = t[79] ^ x[43];
  assign t[62] = t[80] ^ x[45];
  assign t[63] = t[81] ^ x[46];
  assign t[64] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[65] = (x[3]);
  assign t[66] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[67] = (x[12]);
  assign t[68] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[69] = (x[20]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[71] = (x[26]);
  assign t[72] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[73] = (x[32]);
  assign t[74] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[35]);
  assign t[76] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[38]);
  assign t[78] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[41]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[44]);
  assign t[8] = ~(t[20] ^ t[14]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [46:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = t[1] ? t[2] : t[17];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[19] ? x[15] : x[16];
  assign t[13] = ~(t[20] ^ t[14]);
  assign t[14] = ~(t[21] ^ t[22]);
  assign t[15] = ~(t[23] & t[24]);
  assign t[16] = ~(t[19] & t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = t[35] ^ x[5];
  assign t[27] = t[36] ^ x[14];
  assign t[28] = t[37] ^ x[19];
  assign t[29] = t[38] ^ x[25];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[39] ^ x[31];
  assign t[31] = t[40] ^ x[37];
  assign t[32] = t[41] ^ x[40];
  assign t[33] = t[42] ^ x[43];
  assign t[34] = t[43] ^ x[46];
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[46] & t[47]);
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = (~t[58] & t[59]);
  assign t[43] = (~t[60] & t[61]);
  assign t[44] = t[62] ^ x[4];
  assign t[45] = t[63] ^ x[5];
  assign t[46] = t[64] ^ x[13];
  assign t[47] = t[65] ^ x[14];
  assign t[48] = t[66] ^ x[18];
  assign t[49] = t[67] ^ x[19];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[68] ^ x[24];
  assign t[51] = t[69] ^ x[25];
  assign t[52] = t[70] ^ x[30];
  assign t[53] = t[71] ^ x[31];
  assign t[54] = t[72] ^ x[36];
  assign t[55] = t[73] ^ x[37];
  assign t[56] = t[74] ^ x[39];
  assign t[57] = t[75] ^ x[40];
  assign t[58] = t[76] ^ x[42];
  assign t[59] = t[77] ^ x[43];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[78] ^ x[45];
  assign t[61] = t[79] ^ x[46];
  assign t[62] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[63] = (x[2]);
  assign t[64] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[65] = (x[11]);
  assign t[66] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[17]);
  assign t[68] = (x[20] & ~x[21] & ~x[22] & ~x[23]) | (~x[20] & x[21] & ~x[22] & ~x[23]) | (~x[20] & ~x[21] & x[22] & ~x[23]) | (~x[20] & ~x[21] & ~x[22] & x[23]) | (x[20] & x[21] & x[22] & ~x[23]) | (x[20] & x[21] & ~x[22] & x[23]) | (x[20] & ~x[21] & x[22] & x[23]) | (~x[20] & x[21] & x[22] & x[23]);
  assign t[69] = (x[22]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[26] & ~x[27] & ~x[28] & ~x[29]) | (~x[26] & x[27] & ~x[28] & ~x[29]) | (~x[26] & ~x[27] & x[28] & ~x[29]) | (~x[26] & ~x[27] & ~x[28] & x[29]) | (x[26] & x[27] & x[28] & ~x[29]) | (x[26] & x[27] & ~x[28] & x[29]) | (x[26] & ~x[27] & x[28] & x[29]) | (~x[26] & x[27] & x[28] & x[29]);
  assign t[71] = (x[28]);
  assign t[72] = (x[32] & ~x[33] & ~x[34] & ~x[35]) | (~x[32] & x[33] & ~x[34] & ~x[35]) | (~x[32] & ~x[33] & x[34] & ~x[35]) | (~x[32] & ~x[33] & ~x[34] & x[35]) | (x[32] & x[33] & x[34] & ~x[35]) | (x[32] & x[33] & ~x[34] & x[35]) | (x[32] & ~x[33] & x[34] & x[35]) | (~x[32] & x[33] & x[34] & x[35]);
  assign t[73] = (x[34]);
  assign t[74] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[38]);
  assign t[76] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[41]);
  assign t[78] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[44]);
  assign t[7] = t[12] ^ t[13];
  assign t[8] = ~(t[18] ^ t[14]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [46:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = t[1] ? t[2] : t[19];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[21] ^ t[14]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[26] & t[27]);
  assign t[17] = ~(t[18]);
  assign t[18] = ~(t[26]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = t[37] ^ x[5];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[39] ^ x[22];
  assign t[31] = t[40] ^ x[28];
  assign t[32] = t[41] ^ x[34];
  assign t[33] = t[42] ^ x[37];
  assign t[34] = t[43] ^ x[40];
  assign t[35] = t[44] ^ x[43];
  assign t[36] = t[45] ^ x[46];
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[48] & t[49]);
  assign t[39] = (~t[50] & t[51]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[52] & t[53]);
  assign t[41] = (~t[54] & t[55]);
  assign t[42] = (~t[56] & t[57]);
  assign t[43] = (~t[58] & t[59]);
  assign t[44] = (~t[60] & t[61]);
  assign t[45] = (~t[62] & t[63]);
  assign t[46] = t[64] ^ x[4];
  assign t[47] = t[65] ^ x[5];
  assign t[48] = t[66] ^ x[13];
  assign t[49] = t[67] ^ x[14];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[68] ^ x[21];
  assign t[51] = t[69] ^ x[22];
  assign t[52] = t[70] ^ x[27];
  assign t[53] = t[71] ^ x[28];
  assign t[54] = t[72] ^ x[33];
  assign t[55] = t[73] ^ x[34];
  assign t[56] = t[74] ^ x[36];
  assign t[57] = t[75] ^ x[37];
  assign t[58] = t[76] ^ x[39];
  assign t[59] = t[77] ^ x[40];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[78] ^ x[42];
  assign t[61] = t[79] ^ x[43];
  assign t[62] = t[80] ^ x[45];
  assign t[63] = t[81] ^ x[46];
  assign t[64] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[65] = (x[1]);
  assign t[66] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[67] = (x[10]);
  assign t[68] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[69] = (x[18]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[71] = (x[24]);
  assign t[72] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[73] = (x[30]);
  assign t[74] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[35]);
  assign t[76] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[38]);
  assign t[78] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[41]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[44]);
  assign t[8] = ~(t[20] ^ t[14]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [46:0] x;
 output y;

 wire [114:0] t;
  assign t[0] = t[1] ? t[2] : t[52];
  assign t[100] = (x[9]);
  assign t[101] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[102] = (x[17]);
  assign t[103] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[104] = (x[23]);
  assign t[105] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[106] = (x[29]);
  assign t[107] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[108] = (x[35]);
  assign t[109] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (x[38]);
  assign t[111] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[112] = (x[41]);
  assign t[113] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[114] = (x[44]);
  assign t[11] = ~(x[6]);
  assign t[12] = ~(t[54] ^ t[14]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[14] = ~(t[55] ^ t[56]);
  assign t[15] = ~(t[57] & t[58]);
  assign t[16] = ~(t[59] & t[60]);
  assign t[17] = t[19] ? x[15] : x[16];
  assign t[18] = ~(t[20] & t[21]);
  assign t[19] = ~(t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23] | t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[59]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[27] | t[29]);
  assign t[25] = ~(t[30] | t[31]);
  assign t[26] = ~(t[32] & t[33]);
  assign t[27] = ~(t[30]);
  assign t[28] = t[57] ? t[35] : t[34];
  assign t[29] = t[57] ? t[37] : t[36];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[59]);
  assign t[31] = t[57] ? t[35] : t[36];
  assign t[32] = ~(t[38] | t[39]);
  assign t[33] = ~(t[40] & t[41]);
  assign t[34] = ~(t[42] & t[60]);
  assign t[35] = ~(t[43] & t[44]);
  assign t[36] = ~(t[42] & t[44]);
  assign t[37] = ~(t[43] & t[60]);
  assign t[38] = ~(t[30] | t[45]);
  assign t[39] = ~(t[30] | t[46]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[58] | t[44]);
  assign t[41] = t[27] & t[57];
  assign t[42] = x[7] & t[58];
  assign t[43] = ~(x[7] | t[58]);
  assign t[44] = ~(t[60]);
  assign t[45] = t[57] ? t[36] : t[35];
  assign t[46] = t[57] ? t[48] : t[47];
  assign t[47] = ~(x[7] & t[49]);
  assign t[48] = ~(t[50] & t[44]);
  assign t[49] = ~(t[58] | t[60]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(x[7] | t[51]);
  assign t[51] = ~(t[58]);
  assign t[52] = (t[61]);
  assign t[53] = (t[62]);
  assign t[54] = (t[63]);
  assign t[55] = (t[64]);
  assign t[56] = (t[65]);
  assign t[57] = (t[66]);
  assign t[58] = (t[67]);
  assign t[59] = (t[68]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[69]);
  assign t[61] = t[70] ^ x[5];
  assign t[62] = t[71] ^ x[14];
  assign t[63] = t[72] ^ x[22];
  assign t[64] = t[73] ^ x[28];
  assign t[65] = t[74] ^ x[34];
  assign t[66] = t[75] ^ x[37];
  assign t[67] = t[76] ^ x[40];
  assign t[68] = t[77] ^ x[43];
  assign t[69] = t[78] ^ x[46];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (~t[79] & t[80]);
  assign t[71] = (~t[81] & t[82]);
  assign t[72] = (~t[83] & t[84]);
  assign t[73] = (~t[85] & t[86]);
  assign t[74] = (~t[87] & t[88]);
  assign t[75] = (~t[89] & t[90]);
  assign t[76] = (~t[91] & t[92]);
  assign t[77] = (~t[93] & t[94]);
  assign t[78] = (~t[95] & t[96]);
  assign t[79] = t[97] ^ x[4];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[98] ^ x[5];
  assign t[81] = t[99] ^ x[13];
  assign t[82] = t[100] ^ x[14];
  assign t[83] = t[101] ^ x[21];
  assign t[84] = t[102] ^ x[22];
  assign t[85] = t[103] ^ x[27];
  assign t[86] = t[104] ^ x[28];
  assign t[87] = t[105] ^ x[33];
  assign t[88] = t[106] ^ x[34];
  assign t[89] = t[107] ^ x[36];
  assign t[8] = ~(t[53] ^ t[14]);
  assign t[90] = t[108] ^ x[37];
  assign t[91] = t[109] ^ x[39];
  assign t[92] = t[110] ^ x[40];
  assign t[93] = t[111] ^ x[42];
  assign t[94] = t[112] ^ x[43];
  assign t[95] = t[113] ^ x[45];
  assign t[96] = t[114] ^ x[46];
  assign t[97] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[98] = (x[0]);
  assign t[99] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [88:0] x;
 output y;

 wire [279:0] t;
  assign t[0] = t[1] ? t[2] : t[98];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = (t[158]);
  assign t[127] = (t[159]);
  assign t[128] = (t[160]);
  assign t[129] = (t[161]);
  assign t[12] = ~(t[100] ^ t[17]);
  assign t[130] = t[162] ^ x[5];
  assign t[131] = t[163] ^ x[14];
  assign t[132] = t[164] ^ x[22];
  assign t[133] = t[165] ^ x[28];
  assign t[134] = t[166] ^ x[34];
  assign t[135] = t[167] ^ x[37];
  assign t[136] = t[168] ^ x[40];
  assign t[137] = t[169] ^ x[43];
  assign t[138] = t[170] ^ x[46];
  assign t[139] = t[171] ^ x[52];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[58];
  assign t[141] = t[173] ^ x[59];
  assign t[142] = t[174] ^ x[61];
  assign t[143] = t[175] ^ x[64];
  assign t[144] = t[176] ^ x[65];
  assign t[145] = t[177] ^ x[66];
  assign t[146] = t[178] ^ x[67];
  assign t[147] = t[179] ^ x[68];
  assign t[148] = t[180] ^ x[69];
  assign t[149] = t[181] ^ x[71];
  assign t[14] = ~(t[101] ^ t[102]);
  assign t[150] = t[182] ^ x[74];
  assign t[151] = t[183] ^ x[75];
  assign t[152] = t[184] ^ x[76];
  assign t[153] = t[185] ^ x[77];
  assign t[154] = t[186] ^ x[78];
  assign t[155] = t[187] ^ x[79];
  assign t[156] = t[188] ^ x[81];
  assign t[157] = t[189] ^ x[84];
  assign t[158] = t[190] ^ x[85];
  assign t[159] = t[191] ^ x[86];
  assign t[15] = ~(t[103] & t[104]);
  assign t[160] = t[192] ^ x[87];
  assign t[161] = t[193] ^ x[88];
  assign t[162] = (~t[194] & t[195]);
  assign t[163] = (~t[196] & t[197]);
  assign t[164] = (~t[198] & t[199]);
  assign t[165] = (~t[200] & t[201]);
  assign t[166] = (~t[202] & t[203]);
  assign t[167] = (~t[204] & t[205]);
  assign t[168] = (~t[206] & t[207]);
  assign t[169] = (~t[208] & t[209]);
  assign t[16] = ~(t[105] & t[106]);
  assign t[170] = (~t[210] & t[211]);
  assign t[171] = (~t[212] & t[213]);
  assign t[172] = (~t[214] & t[215]);
  assign t[173] = (~t[194] & t[216]);
  assign t[174] = (~t[196] & t[217]);
  assign t[175] = (~t[198] & t[218]);
  assign t[176] = (~t[202] & t[219]);
  assign t[177] = (~t[200] & t[220]);
  assign t[178] = (~t[214] & t[221]);
  assign t[179] = (~t[212] & t[222]);
  assign t[17] = ~(t[107] ^ t[108]);
  assign t[180] = (~t[194] & t[223]);
  assign t[181] = (~t[196] & t[224]);
  assign t[182] = (~t[198] & t[225]);
  assign t[183] = (~t[200] & t[226]);
  assign t[184] = (~t[202] & t[227]);
  assign t[185] = (~t[214] & t[228]);
  assign t[186] = (~t[212] & t[229]);
  assign t[187] = (~t[194] & t[230]);
  assign t[188] = (~t[196] & t[231]);
  assign t[189] = (~t[198] & t[232]);
  assign t[18] = t[20] ? x[15] : x[16];
  assign t[190] = (~t[200] & t[233]);
  assign t[191] = (~t[202] & t[234]);
  assign t[192] = (~t[214] & t[235]);
  assign t[193] = (~t[212] & t[236]);
  assign t[194] = t[237] ^ x[4];
  assign t[195] = t[238] ^ x[5];
  assign t[196] = t[239] ^ x[13];
  assign t[197] = t[240] ^ x[14];
  assign t[198] = t[241] ^ x[21];
  assign t[199] = t[242] ^ x[22];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[27];
  assign t[201] = t[244] ^ x[28];
  assign t[202] = t[245] ^ x[33];
  assign t[203] = t[246] ^ x[34];
  assign t[204] = t[247] ^ x[36];
  assign t[205] = t[248] ^ x[37];
  assign t[206] = t[249] ^ x[39];
  assign t[207] = t[250] ^ x[40];
  assign t[208] = t[251] ^ x[42];
  assign t[209] = t[252] ^ x[43];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[45];
  assign t[211] = t[254] ^ x[46];
  assign t[212] = t[255] ^ x[51];
  assign t[213] = t[256] ^ x[52];
  assign t[214] = t[257] ^ x[57];
  assign t[215] = t[258] ^ x[58];
  assign t[216] = t[259] ^ x[59];
  assign t[217] = t[260] ^ x[61];
  assign t[218] = t[261] ^ x[64];
  assign t[219] = t[262] ^ x[65];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[66];
  assign t[221] = t[264] ^ x[67];
  assign t[222] = t[265] ^ x[68];
  assign t[223] = t[266] ^ x[69];
  assign t[224] = t[267] ^ x[71];
  assign t[225] = t[268] ^ x[74];
  assign t[226] = t[269] ^ x[75];
  assign t[227] = t[270] ^ x[76];
  assign t[228] = t[271] ^ x[77];
  assign t[229] = t[272] ^ x[78];
  assign t[22] = ~(t[26] | t[27]);
  assign t[230] = t[273] ^ x[79];
  assign t[231] = t[274] ^ x[81];
  assign t[232] = t[275] ^ x[84];
  assign t[233] = t[276] ^ x[85];
  assign t[234] = t[277] ^ x[86];
  assign t[235] = t[278] ^ x[87];
  assign t[236] = t[279] ^ x[88];
  assign t[237] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[238] = (x[0]);
  assign t[239] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[23] = ~(t[105]);
  assign t[240] = (x[9]);
  assign t[241] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[242] = (x[17]);
  assign t[243] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[244] = (x[23]);
  assign t[245] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[246] = (x[29]);
  assign t[247] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[248] = (x[35]);
  assign t[249] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[24] = ~(t[28] | t[29]);
  assign t[250] = (x[38]);
  assign t[251] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[252] = (x[41]);
  assign t[253] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[254] = (x[44]);
  assign t[255] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[256] = (x[47]);
  assign t[257] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[258] = (x[53]);
  assign t[259] = (x[1]);
  assign t[25] = ~(t[28] | t[30]);
  assign t[260] = (x[10]);
  assign t[261] = (x[18]);
  assign t[262] = (x[30]);
  assign t[263] = (x[24]);
  assign t[264] = (x[54]);
  assign t[265] = (x[48]);
  assign t[266] = (x[2]);
  assign t[267] = (x[11]);
  assign t[268] = (x[19]);
  assign t[269] = (x[25]);
  assign t[26] = t[31] | t[32];
  assign t[270] = (x[31]);
  assign t[271] = (x[55]);
  assign t[272] = (x[49]);
  assign t[273] = (x[3]);
  assign t[274] = (x[12]);
  assign t[275] = (x[20]);
  assign t[276] = (x[26]);
  assign t[277] = (x[32]);
  assign t[278] = (x[56]);
  assign t[279] = (x[50]);
  assign t[27] = ~(t[33] & t[34]);
  assign t[28] = ~(t[35]);
  assign t[29] = t[103] ? t[37] : t[36];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[103] ? t[39] : t[38];
  assign t[31] = ~(t[40] & t[41]);
  assign t[32] = ~(t[28] | t[42]);
  assign t[33] = ~(t[43] | t[44]);
  assign t[34] = t[35] | t[45];
  assign t[35] = ~(t[105]);
  assign t[36] = ~(t[46] & t[47]);
  assign t[37] = ~(t[48] & t[106]);
  assign t[38] = ~(t[106] & t[49]);
  assign t[39] = ~(x[7] & t[50]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[51] | t[52]);
  assign t[41] = ~(t[53] & t[54]);
  assign t[42] = t[103] ? t[38] : t[39];
  assign t[43] = ~(t[55]);
  assign t[44] = ~(t[28] | t[56]);
  assign t[45] = t[103] ? t[39] : t[57];
  assign t[46] = ~(x[7] | t[104]);
  assign t[47] = ~(t[106]);
  assign t[48] = x[7] & t[104];
  assign t[49] = ~(x[7] | t[58]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[104] | t[106]);
  assign t[51] = ~(t[35] | t[59]);
  assign t[52] = ~(t[35] | t[60]);
  assign t[53] = ~(t[104] | t[47]);
  assign t[54] = t[28] & t[103];
  assign t[55] = ~(t[61] & t[62]);
  assign t[56] = t[103] ? t[63] : t[57];
  assign t[57] = ~(t[49] & t[47]);
  assign t[58] = ~(t[104]);
  assign t[59] = t[103] ? t[64] : t[36];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[103] ? t[57] : t[39];
  assign t[61] = ~(t[35] | t[103]);
  assign t[62] = ~(t[38] & t[63]);
  assign t[63] = ~(x[7] & t[53]);
  assign t[64] = ~(t[48] & t[47]);
  assign t[65] = t[1] ? t[66] : t[109];
  assign t[66] = x[6] ? t[68] : t[67];
  assign t[67] = x[7] ? t[70] : t[69];
  assign t[68] = t[71] ^ x[60];
  assign t[69] = t[72] ^ t[73];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[110] ^ t[74]);
  assign t[71] = x[62] ^ x[63];
  assign t[72] = t[20] ? x[62] : x[63];
  assign t[73] = ~(t[111] ^ t[75]);
  assign t[74] = ~(t[112] ^ t[113]);
  assign t[75] = ~(t[114] ^ t[115]);
  assign t[76] = t[1] ? t[77] : t[116];
  assign t[77] = x[6] ? t[79] : t[78];
  assign t[78] = x[7] ? t[81] : t[80];
  assign t[79] = t[82] ^ x[70];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[83] ^ t[84];
  assign t[81] = ~(t[117] ^ t[85]);
  assign t[82] = x[72] ^ x[73];
  assign t[83] = t[20] ? x[72] : x[73];
  assign t[84] = ~(t[118] ^ t[86]);
  assign t[85] = ~(t[119] ^ t[120]);
  assign t[86] = ~(t[121] ^ t[122]);
  assign t[87] = t[1] ? t[88] : t[123];
  assign t[88] = x[6] ? t[90] : t[89];
  assign t[89] = x[7] ? t[92] : t[91];
  assign t[8] = ~(t[99] ^ t[14]);
  assign t[90] = t[93] ^ x[80];
  assign t[91] = t[94] ^ t[95];
  assign t[92] = ~(t[124] ^ t[96]);
  assign t[93] = x[82] ^ x[83];
  assign t[94] = t[20] ? x[82] : x[83];
  assign t[95] = ~(t[125] ^ t[97]);
  assign t[96] = ~(t[126] ^ t[127]);
  assign t[97] = ~(t[128] ^ t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[65] & ~t[76] & ~t[87]) | (~t[0] & t[65] & ~t[76] & ~t[87]) | (~t[0] & ~t[65] & t[76] & ~t[87]) | (~t[0] & ~t[65] & ~t[76] & t[87]) | (t[0] & t[65] & t[76] & ~t[87]) | (t[0] & t[65] & ~t[76] & t[87]) | (t[0] & ~t[65] & t[76] & t[87]) | (~t[0] & t[65] & t[76] & t[87]);
endmodule

module R2ind146(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[2]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[11]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[19]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[25]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[49]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[1]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[10]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[18]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[48]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[54]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [58:0] x;
 output y;

 wire [141:0] t;
  assign t[0] = t[1] ? t[2] : t[65];
  assign t[100] = t[122] ^ x[13];
  assign t[101] = t[123] ^ x[14];
  assign t[102] = t[124] ^ x[21];
  assign t[103] = t[125] ^ x[22];
  assign t[104] = t[126] ^ x[27];
  assign t[105] = t[127] ^ x[28];
  assign t[106] = t[128] ^ x[33];
  assign t[107] = t[129] ^ x[34];
  assign t[108] = t[130] ^ x[36];
  assign t[109] = t[131] ^ x[37];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[132] ^ x[39];
  assign t[111] = t[133] ^ x[40];
  assign t[112] = t[134] ^ x[42];
  assign t[113] = t[135] ^ x[43];
  assign t[114] = t[136] ^ x[45];
  assign t[115] = t[137] ^ x[46];
  assign t[116] = t[138] ^ x[51];
  assign t[117] = t[139] ^ x[52];
  assign t[118] = t[140] ^ x[57];
  assign t[119] = t[141] ^ x[58];
  assign t[11] = ~(x[6]);
  assign t[120] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[121] = (x[0]);
  assign t[122] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[123] = (x[9]);
  assign t[124] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[125] = (x[17]);
  assign t[126] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[127] = (x[23]);
  assign t[128] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[129] = (x[29]);
  assign t[12] = ~(t[67] ^ t[17]);
  assign t[130] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[35]);
  assign t[132] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[133] = (x[38]);
  assign t[134] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[135] = (x[41]);
  assign t[136] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[137] = (x[44]);
  assign t[138] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[139] = (x[47]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[141] = (x[53]);
  assign t[14] = ~(t[68] ^ t[69]);
  assign t[15] = ~(t[70] & t[71]);
  assign t[16] = ~(t[72] & t[73]);
  assign t[17] = ~(t[74] ^ t[75]);
  assign t[18] = t[20] ? x[15] : x[16];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[72]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[25] = ~(t[28] | t[30]);
  assign t[26] = t[31] | t[32];
  assign t[27] = ~(t[33] & t[34]);
  assign t[28] = ~(t[35]);
  assign t[29] = t[70] ? t[37] : t[36];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[70] ? t[39] : t[38];
  assign t[31] = ~(t[40] & t[41]);
  assign t[32] = ~(t[28] | t[42]);
  assign t[33] = ~(t[43] | t[44]);
  assign t[34] = t[35] | t[45];
  assign t[35] = ~(t[72]);
  assign t[36] = ~(t[46] & t[47]);
  assign t[37] = ~(t[48] & t[73]);
  assign t[38] = ~(t[73] & t[49]);
  assign t[39] = ~(x[7] & t[50]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[51] | t[52]);
  assign t[41] = ~(t[53] & t[54]);
  assign t[42] = t[70] ? t[38] : t[39];
  assign t[43] = ~(t[55]);
  assign t[44] = ~(t[28] | t[56]);
  assign t[45] = t[70] ? t[39] : t[57];
  assign t[46] = ~(x[7] | t[71]);
  assign t[47] = ~(t[73]);
  assign t[48] = x[7] & t[71];
  assign t[49] = ~(x[7] | t[58]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[71] | t[73]);
  assign t[51] = ~(t[35] | t[59]);
  assign t[52] = ~(t[35] | t[60]);
  assign t[53] = ~(t[71] | t[47]);
  assign t[54] = t[28] & t[70];
  assign t[55] = ~(t[61] & t[62]);
  assign t[56] = t[70] ? t[63] : t[57];
  assign t[57] = ~(t[49] & t[47]);
  assign t[58] = ~(t[71]);
  assign t[59] = t[70] ? t[64] : t[36];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[70] ? t[57] : t[39];
  assign t[61] = ~(t[35] | t[70]);
  assign t[62] = ~(t[38] & t[63]);
  assign t[63] = ~(x[7] & t[53]);
  assign t[64] = ~(t[48] & t[47]);
  assign t[65] = (t[76]);
  assign t[66] = (t[77]);
  assign t[67] = (t[78]);
  assign t[68] = (t[79]);
  assign t[69] = (t[80]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[81]);
  assign t[71] = (t[82]);
  assign t[72] = (t[83]);
  assign t[73] = (t[84]);
  assign t[74] = (t[85]);
  assign t[75] = (t[86]);
  assign t[76] = t[87] ^ x[5];
  assign t[77] = t[88] ^ x[14];
  assign t[78] = t[89] ^ x[22];
  assign t[79] = t[90] ^ x[28];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[91] ^ x[34];
  assign t[81] = t[92] ^ x[37];
  assign t[82] = t[93] ^ x[40];
  assign t[83] = t[94] ^ x[43];
  assign t[84] = t[95] ^ x[46];
  assign t[85] = t[96] ^ x[52];
  assign t[86] = t[97] ^ x[58];
  assign t[87] = (~t[98] & t[99]);
  assign t[88] = (~t[100] & t[101]);
  assign t[89] = (~t[102] & t[103]);
  assign t[8] = ~(t[66] ^ t[14]);
  assign t[90] = (~t[104] & t[105]);
  assign t[91] = (~t[106] & t[107]);
  assign t[92] = (~t[108] & t[109]);
  assign t[93] = (~t[110] & t[111]);
  assign t[94] = (~t[112] & t[113]);
  assign t[95] = (~t[114] & t[115]);
  assign t[96] = (~t[116] & t[117]);
  assign t[97] = (~t[118] & t[119]);
  assign t[98] = t[120] ^ x[4];
  assign t[99] = t[121] ^ x[5];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [88:0] x;
 output y;

 wire [265:0] t;
  assign t[0] = t[1] ? t[2] : t[84];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = t[148] ^ x[5];
  assign t[117] = t[149] ^ x[14];
  assign t[118] = t[150] ^ x[22];
  assign t[119] = t[151] ^ x[28];
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[34];
  assign t[121] = t[153] ^ x[37];
  assign t[122] = t[154] ^ x[40];
  assign t[123] = t[155] ^ x[43];
  assign t[124] = t[156] ^ x[46];
  assign t[125] = t[157] ^ x[52];
  assign t[126] = t[158] ^ x[58];
  assign t[127] = t[159] ^ x[59];
  assign t[128] = t[160] ^ x[61];
  assign t[129] = t[161] ^ x[64];
  assign t[12] = ~(t[86] ^ t[17]);
  assign t[130] = t[162] ^ x[65];
  assign t[131] = t[163] ^ x[66];
  assign t[132] = t[164] ^ x[67];
  assign t[133] = t[165] ^ x[68];
  assign t[134] = t[166] ^ x[69];
  assign t[135] = t[167] ^ x[71];
  assign t[136] = t[168] ^ x[74];
  assign t[137] = t[169] ^ x[75];
  assign t[138] = t[170] ^ x[76];
  assign t[139] = t[171] ^ x[77];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[78];
  assign t[141] = t[173] ^ x[79];
  assign t[142] = t[174] ^ x[81];
  assign t[143] = t[175] ^ x[84];
  assign t[144] = t[176] ^ x[85];
  assign t[145] = t[177] ^ x[86];
  assign t[146] = t[178] ^ x[87];
  assign t[147] = t[179] ^ x[88];
  assign t[148] = (~t[180] & t[181]);
  assign t[149] = (~t[182] & t[183]);
  assign t[14] = ~(t[87] ^ t[88]);
  assign t[150] = (~t[184] & t[185]);
  assign t[151] = (~t[186] & t[187]);
  assign t[152] = (~t[188] & t[189]);
  assign t[153] = (~t[190] & t[191]);
  assign t[154] = (~t[192] & t[193]);
  assign t[155] = (~t[194] & t[195]);
  assign t[156] = (~t[196] & t[197]);
  assign t[157] = (~t[198] & t[199]);
  assign t[158] = (~t[200] & t[201]);
  assign t[159] = (~t[180] & t[202]);
  assign t[15] = ~(t[89] & t[90]);
  assign t[160] = (~t[182] & t[203]);
  assign t[161] = (~t[184] & t[204]);
  assign t[162] = (~t[188] & t[205]);
  assign t[163] = (~t[186] & t[206]);
  assign t[164] = (~t[200] & t[207]);
  assign t[165] = (~t[198] & t[208]);
  assign t[166] = (~t[180] & t[209]);
  assign t[167] = (~t[182] & t[210]);
  assign t[168] = (~t[184] & t[211]);
  assign t[169] = (~t[188] & t[212]);
  assign t[16] = ~(t[91] & t[92]);
  assign t[170] = (~t[186] & t[213]);
  assign t[171] = (~t[198] & t[214]);
  assign t[172] = (~t[200] & t[215]);
  assign t[173] = (~t[180] & t[216]);
  assign t[174] = (~t[182] & t[217]);
  assign t[175] = (~t[184] & t[218]);
  assign t[176] = (~t[188] & t[219]);
  assign t[177] = (~t[186] & t[220]);
  assign t[178] = (~t[198] & t[221]);
  assign t[179] = (~t[200] & t[222]);
  assign t[17] = ~(t[93] ^ t[94]);
  assign t[180] = t[223] ^ x[4];
  assign t[181] = t[224] ^ x[5];
  assign t[182] = t[225] ^ x[13];
  assign t[183] = t[226] ^ x[14];
  assign t[184] = t[227] ^ x[21];
  assign t[185] = t[228] ^ x[22];
  assign t[186] = t[229] ^ x[27];
  assign t[187] = t[230] ^ x[28];
  assign t[188] = t[231] ^ x[33];
  assign t[189] = t[232] ^ x[34];
  assign t[18] = t[20] ? x[15] : x[16];
  assign t[190] = t[233] ^ x[36];
  assign t[191] = t[234] ^ x[37];
  assign t[192] = t[235] ^ x[39];
  assign t[193] = t[236] ^ x[40];
  assign t[194] = t[237] ^ x[42];
  assign t[195] = t[238] ^ x[43];
  assign t[196] = t[239] ^ x[45];
  assign t[197] = t[240] ^ x[46];
  assign t[198] = t[241] ^ x[51];
  assign t[199] = t[242] ^ x[52];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[57];
  assign t[201] = t[244] ^ x[58];
  assign t[202] = t[245] ^ x[59];
  assign t[203] = t[246] ^ x[61];
  assign t[204] = t[247] ^ x[64];
  assign t[205] = t[248] ^ x[65];
  assign t[206] = t[249] ^ x[66];
  assign t[207] = t[250] ^ x[67];
  assign t[208] = t[251] ^ x[68];
  assign t[209] = t[252] ^ x[69];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[71];
  assign t[211] = t[254] ^ x[74];
  assign t[212] = t[255] ^ x[75];
  assign t[213] = t[256] ^ x[76];
  assign t[214] = t[257] ^ x[77];
  assign t[215] = t[258] ^ x[78];
  assign t[216] = t[259] ^ x[79];
  assign t[217] = t[260] ^ x[81];
  assign t[218] = t[261] ^ x[84];
  assign t[219] = t[262] ^ x[85];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[86];
  assign t[221] = t[264] ^ x[87];
  assign t[222] = t[265] ^ x[88];
  assign t[223] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[224] = (x[0]);
  assign t[225] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[226] = (x[9]);
  assign t[227] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[228] = (x[17]);
  assign t[229] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[230] = (x[23]);
  assign t[231] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[232] = (x[29]);
  assign t[233] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[234] = (x[35]);
  assign t[235] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[236] = (x[38]);
  assign t[237] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[238] = (x[41]);
  assign t[239] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[23] = ~(t[91]);
  assign t[240] = (x[44]);
  assign t[241] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[242] = (x[47]);
  assign t[243] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[244] = (x[53]);
  assign t[245] = (x[1]);
  assign t[246] = (x[10]);
  assign t[247] = (x[18]);
  assign t[248] = (x[30]);
  assign t[249] = (x[24]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[250] = (x[54]);
  assign t[251] = (x[48]);
  assign t[252] = (x[2]);
  assign t[253] = (x[11]);
  assign t[254] = (x[19]);
  assign t[255] = (x[31]);
  assign t[256] = (x[25]);
  assign t[257] = (x[49]);
  assign t[258] = (x[55]);
  assign t[259] = (x[3]);
  assign t[25] = ~(t[30] & t[31]);
  assign t[260] = (x[12]);
  assign t[261] = (x[20]);
  assign t[262] = (x[32]);
  assign t[263] = (x[26]);
  assign t[264] = (x[50]);
  assign t[265] = (x[56]);
  assign t[26] = ~(t[90] | t[32]);
  assign t[27] = t[28] & t[89];
  assign t[28] = ~(t[33]);
  assign t[29] = t[89] ? t[35] : t[34];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[33] & t[38]);
  assign t[32] = ~(t[92]);
  assign t[33] = ~(t[91]);
  assign t[34] = ~(t[39] & t[32]);
  assign t[35] = ~(t[40] & t[92]);
  assign t[36] = ~(t[33] | t[41]);
  assign t[37] = ~(t[28] | t[42]);
  assign t[38] = ~(t[43] & t[44]);
  assign t[39] = ~(x[7] | t[90]);
  assign t[3] = ~(t[6]);
  assign t[40] = x[7] & t[90];
  assign t[41] = t[89] ? t[34] : t[45];
  assign t[42] = t[89] ? t[47] : t[46];
  assign t[43] = ~(x[7] & t[48]);
  assign t[44] = ~(t[92] & t[49]);
  assign t[45] = ~(t[40] & t[32]);
  assign t[46] = ~(x[7] & t[26]);
  assign t[47] = ~(t[49] & t[32]);
  assign t[48] = ~(t[90] | t[92]);
  assign t[49] = ~(x[7] | t[50]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[90]);
  assign t[51] = t[1] ? t[52] : t[95];
  assign t[52] = x[6] ? t[54] : t[53];
  assign t[53] = x[7] ? t[56] : t[55];
  assign t[54] = t[57] ^ x[60];
  assign t[55] = t[58] ^ t[59];
  assign t[56] = ~(t[96] ^ t[60]);
  assign t[57] = x[62] ^ x[63];
  assign t[58] = t[20] ? x[62] : x[63];
  assign t[59] = ~(t[97] ^ t[61]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[98] ^ t[99]);
  assign t[61] = ~(t[100] ^ t[101]);
  assign t[62] = t[1] ? t[63] : t[102];
  assign t[63] = x[6] ? t[65] : t[64];
  assign t[64] = x[7] ? t[67] : t[66];
  assign t[65] = t[68] ^ x[70];
  assign t[66] = t[69] ^ t[70];
  assign t[67] = ~(t[103] ^ t[71]);
  assign t[68] = x[72] ^ x[73];
  assign t[69] = t[20] ? x[72] : x[73];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104] ^ t[72]);
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = ~(t[107] ^ t[108]);
  assign t[73] = t[1] ? t[74] : t[109];
  assign t[74] = x[6] ? t[76] : t[75];
  assign t[75] = x[7] ? t[78] : t[77];
  assign t[76] = t[79] ^ x[80];
  assign t[77] = t[80] ^ t[81];
  assign t[78] = ~(t[110] ^ t[82]);
  assign t[79] = x[82] ^ x[83];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[20] ? x[82] : x[83];
  assign t[81] = ~(t[111] ^ t[83]);
  assign t[82] = ~(t[112] ^ t[113]);
  assign t[83] = ~(t[114] ^ t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[85] ^ t[14]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[51] & ~t[62] & ~t[73]) | (~t[0] & t[51] & ~t[62] & ~t[73]) | (~t[0] & ~t[51] & t[62] & ~t[73]) | (~t[0] & ~t[51] & ~t[62] & t[73]) | (t[0] & t[51] & t[62] & ~t[73]) | (t[0] & t[51] & ~t[62] & t[73]) | (t[0] & ~t[51] & t[62] & t[73]) | (~t[0] & t[51] & t[62] & t[73]);
endmodule

module R2ind151(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[2]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[11]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[19]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[25]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[49]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[15] : x[16];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[1]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[10]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[18]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[48]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[54]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [58:0] x;
 output y;

 wire [127:0] t;
  assign t[0] = t[1] ? t[2] : t[51];
  assign t[100] = t[122] ^ x[45];
  assign t[101] = t[123] ^ x[46];
  assign t[102] = t[124] ^ x[51];
  assign t[103] = t[125] ^ x[52];
  assign t[104] = t[126] ^ x[57];
  assign t[105] = t[127] ^ x[58];
  assign t[106] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[107] = (x[0]);
  assign t[108] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[109] = (x[9]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[111] = (x[17]);
  assign t[112] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[113] = (x[23]);
  assign t[114] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[115] = (x[29]);
  assign t[116] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[117] = (x[35]);
  assign t[118] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[119] = (x[38]);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[121] = (x[41]);
  assign t[122] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[44]);
  assign t[124] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[125] = (x[47]);
  assign t[126] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[127] = (x[53]);
  assign t[12] = ~(t[53] ^ t[17]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[54] ^ t[55]);
  assign t[15] = ~(t[56] & t[57]);
  assign t[16] = ~(t[58] & t[59]);
  assign t[17] = ~(t[60] ^ t[61]);
  assign t[18] = t[20] ? x[15] : x[16];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[58]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[25] = ~(t[30] & t[31]);
  assign t[26] = ~(t[57] | t[32]);
  assign t[27] = t[28] & t[56];
  assign t[28] = ~(t[33]);
  assign t[29] = t[56] ? t[35] : t[34];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[36] | t[37]);
  assign t[31] = ~(t[33] & t[38]);
  assign t[32] = ~(t[59]);
  assign t[33] = ~(t[58]);
  assign t[34] = ~(t[39] & t[32]);
  assign t[35] = ~(t[40] & t[59]);
  assign t[36] = ~(t[33] | t[41]);
  assign t[37] = ~(t[28] | t[42]);
  assign t[38] = ~(t[43] & t[44]);
  assign t[39] = ~(x[7] | t[57]);
  assign t[3] = ~(t[6]);
  assign t[40] = x[7] & t[57];
  assign t[41] = t[56] ? t[34] : t[45];
  assign t[42] = t[56] ? t[47] : t[46];
  assign t[43] = ~(x[7] & t[48]);
  assign t[44] = ~(t[59] & t[49]);
  assign t[45] = ~(t[40] & t[32]);
  assign t[46] = ~(x[7] & t[26]);
  assign t[47] = ~(t[49] & t[32]);
  assign t[48] = ~(t[57] | t[59]);
  assign t[49] = ~(x[7] | t[50]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[57]);
  assign t[51] = (t[62]);
  assign t[52] = (t[63]);
  assign t[53] = (t[64]);
  assign t[54] = (t[65]);
  assign t[55] = (t[66]);
  assign t[56] = (t[67]);
  assign t[57] = (t[68]);
  assign t[58] = (t[69]);
  assign t[59] = (t[70]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = t[73] ^ x[5];
  assign t[63] = t[74] ^ x[14];
  assign t[64] = t[75] ^ x[22];
  assign t[65] = t[76] ^ x[28];
  assign t[66] = t[77] ^ x[34];
  assign t[67] = t[78] ^ x[37];
  assign t[68] = t[79] ^ x[40];
  assign t[69] = t[80] ^ x[43];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[81] ^ x[46];
  assign t[71] = t[82] ^ x[52];
  assign t[72] = t[83] ^ x[58];
  assign t[73] = (~t[84] & t[85]);
  assign t[74] = (~t[86] & t[87]);
  assign t[75] = (~t[88] & t[89]);
  assign t[76] = (~t[90] & t[91]);
  assign t[77] = (~t[92] & t[93]);
  assign t[78] = (~t[94] & t[95]);
  assign t[79] = (~t[96] & t[97]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[98] & t[99]);
  assign t[81] = (~t[100] & t[101]);
  assign t[82] = (~t[102] & t[103]);
  assign t[83] = (~t[104] & t[105]);
  assign t[84] = t[106] ^ x[4];
  assign t[85] = t[107] ^ x[5];
  assign t[86] = t[108] ^ x[13];
  assign t[87] = t[109] ^ x[14];
  assign t[88] = t[110] ^ x[21];
  assign t[89] = t[111] ^ x[22];
  assign t[8] = ~(t[52] ^ t[14]);
  assign t[90] = t[112] ^ x[27];
  assign t[91] = t[113] ^ x[28];
  assign t[92] = t[114] ^ x[33];
  assign t[93] = t[115] ^ x[34];
  assign t[94] = t[116] ^ x[36];
  assign t[95] = t[117] ^ x[37];
  assign t[96] = t[118] ^ x[39];
  assign t[97] = t[119] ^ x[40];
  assign t[98] = t[120] ^ x[42];
  assign t[99] = t[121] ^ x[43];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [88:0] x;
 output y;

 wire [265:0] t;
  assign t[0] = t[1] ? t[2] : t[84];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = t[148] ^ x[5];
  assign t[117] = t[149] ^ x[14];
  assign t[118] = t[150] ^ x[22];
  assign t[119] = t[151] ^ x[28];
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[34];
  assign t[121] = t[153] ^ x[37];
  assign t[122] = t[154] ^ x[40];
  assign t[123] = t[155] ^ x[43];
  assign t[124] = t[156] ^ x[46];
  assign t[125] = t[157] ^ x[52];
  assign t[126] = t[158] ^ x[58];
  assign t[127] = t[159] ^ x[59];
  assign t[128] = t[160] ^ x[61];
  assign t[129] = t[161] ^ x[64];
  assign t[12] = ~(t[86] ^ t[17]);
  assign t[130] = t[162] ^ x[65];
  assign t[131] = t[163] ^ x[66];
  assign t[132] = t[164] ^ x[67];
  assign t[133] = t[165] ^ x[68];
  assign t[134] = t[166] ^ x[69];
  assign t[135] = t[167] ^ x[71];
  assign t[136] = t[168] ^ x[74];
  assign t[137] = t[169] ^ x[75];
  assign t[138] = t[170] ^ x[76];
  assign t[139] = t[171] ^ x[77];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[78];
  assign t[141] = t[173] ^ x[79];
  assign t[142] = t[174] ^ x[81];
  assign t[143] = t[175] ^ x[84];
  assign t[144] = t[176] ^ x[85];
  assign t[145] = t[177] ^ x[86];
  assign t[146] = t[178] ^ x[87];
  assign t[147] = t[179] ^ x[88];
  assign t[148] = (~t[180] & t[181]);
  assign t[149] = (~t[182] & t[183]);
  assign t[14] = ~(t[87] ^ t[88]);
  assign t[150] = (~t[184] & t[185]);
  assign t[151] = (~t[186] & t[187]);
  assign t[152] = (~t[188] & t[189]);
  assign t[153] = (~t[190] & t[191]);
  assign t[154] = (~t[192] & t[193]);
  assign t[155] = (~t[194] & t[195]);
  assign t[156] = (~t[196] & t[197]);
  assign t[157] = (~t[198] & t[199]);
  assign t[158] = (~t[200] & t[201]);
  assign t[159] = (~t[180] & t[202]);
  assign t[15] = ~(t[89] & t[90]);
  assign t[160] = (~t[182] & t[203]);
  assign t[161] = (~t[184] & t[204]);
  assign t[162] = (~t[188] & t[205]);
  assign t[163] = (~t[186] & t[206]);
  assign t[164] = (~t[200] & t[207]);
  assign t[165] = (~t[198] & t[208]);
  assign t[166] = (~t[180] & t[209]);
  assign t[167] = (~t[182] & t[210]);
  assign t[168] = (~t[184] & t[211]);
  assign t[169] = (~t[186] & t[212]);
  assign t[16] = ~(t[91] & t[92]);
  assign t[170] = (~t[188] & t[213]);
  assign t[171] = (~t[198] & t[214]);
  assign t[172] = (~t[200] & t[215]);
  assign t[173] = (~t[180] & t[216]);
  assign t[174] = (~t[182] & t[217]);
  assign t[175] = (~t[184] & t[218]);
  assign t[176] = (~t[186] & t[219]);
  assign t[177] = (~t[188] & t[220]);
  assign t[178] = (~t[198] & t[221]);
  assign t[179] = (~t[200] & t[222]);
  assign t[17] = ~(t[93] ^ t[94]);
  assign t[180] = t[223] ^ x[4];
  assign t[181] = t[224] ^ x[5];
  assign t[182] = t[225] ^ x[13];
  assign t[183] = t[226] ^ x[14];
  assign t[184] = t[227] ^ x[21];
  assign t[185] = t[228] ^ x[22];
  assign t[186] = t[229] ^ x[27];
  assign t[187] = t[230] ^ x[28];
  assign t[188] = t[231] ^ x[33];
  assign t[189] = t[232] ^ x[34];
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[190] = t[233] ^ x[36];
  assign t[191] = t[234] ^ x[37];
  assign t[192] = t[235] ^ x[39];
  assign t[193] = t[236] ^ x[40];
  assign t[194] = t[237] ^ x[42];
  assign t[195] = t[238] ^ x[43];
  assign t[196] = t[239] ^ x[45];
  assign t[197] = t[240] ^ x[46];
  assign t[198] = t[241] ^ x[51];
  assign t[199] = t[242] ^ x[52];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[57];
  assign t[201] = t[244] ^ x[58];
  assign t[202] = t[245] ^ x[59];
  assign t[203] = t[246] ^ x[61];
  assign t[204] = t[247] ^ x[64];
  assign t[205] = t[248] ^ x[65];
  assign t[206] = t[249] ^ x[66];
  assign t[207] = t[250] ^ x[67];
  assign t[208] = t[251] ^ x[68];
  assign t[209] = t[252] ^ x[69];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[71];
  assign t[211] = t[254] ^ x[74];
  assign t[212] = t[255] ^ x[75];
  assign t[213] = t[256] ^ x[76];
  assign t[214] = t[257] ^ x[77];
  assign t[215] = t[258] ^ x[78];
  assign t[216] = t[259] ^ x[79];
  assign t[217] = t[260] ^ x[81];
  assign t[218] = t[261] ^ x[84];
  assign t[219] = t[262] ^ x[85];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[86];
  assign t[221] = t[264] ^ x[87];
  assign t[222] = t[265] ^ x[88];
  assign t[223] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[224] = (x[0]);
  assign t[225] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[226] = (x[9]);
  assign t[227] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[228] = (x[17]);
  assign t[229] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[230] = (x[23]);
  assign t[231] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[232] = (x[29]);
  assign t[233] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[234] = (x[35]);
  assign t[235] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[236] = (x[38]);
  assign t[237] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[238] = (x[41]);
  assign t[239] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[23] = ~(t[91]);
  assign t[240] = (x[44]);
  assign t[241] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[242] = (x[47]);
  assign t[243] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[244] = (x[53]);
  assign t[245] = (x[1]);
  assign t[246] = (x[10]);
  assign t[247] = (x[18]);
  assign t[248] = (x[30]);
  assign t[249] = (x[24]);
  assign t[24] = ~(t[28] & t[29]);
  assign t[250] = (x[54]);
  assign t[251] = (x[48]);
  assign t[252] = (x[2]);
  assign t[253] = (x[11]);
  assign t[254] = (x[19]);
  assign t[255] = (x[25]);
  assign t[256] = (x[31]);
  assign t[257] = (x[49]);
  assign t[258] = (x[55]);
  assign t[259] = (x[3]);
  assign t[25] = t[30] | t[31];
  assign t[260] = (x[12]);
  assign t[261] = (x[20]);
  assign t[262] = (x[26]);
  assign t[263] = (x[32]);
  assign t[264] = (x[50]);
  assign t[265] = (x[56]);
  assign t[26] = t[92] & t[32];
  assign t[27] = t[33] | t[34];
  assign t[28] = ~(t[32] & t[35]);
  assign t[29] = ~(t[36] & t[37]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[38] | t[39]);
  assign t[31] = ~(t[38] | t[40]);
  assign t[32] = ~(t[41] | t[89]);
  assign t[33] = ~(x[7] | t[90]);
  assign t[34] = x[7] & t[90];
  assign t[35] = ~(t[42] & t[43]);
  assign t[36] = ~(t[90] | t[44]);
  assign t[37] = t[38] & t[89];
  assign t[38] = ~(t[41]);
  assign t[39] = t[89] ? t[42] : t[45];
  assign t[3] = ~(t[6]);
  assign t[40] = t[89] ? t[47] : t[46];
  assign t[41] = ~(t[91]);
  assign t[42] = ~(t[92] & t[48]);
  assign t[43] = ~(x[7] & t[36]);
  assign t[44] = ~(t[92]);
  assign t[45] = ~(x[7] & t[49]);
  assign t[46] = ~(t[34] & t[44]);
  assign t[47] = ~(t[33] & t[92]);
  assign t[48] = ~(x[7] | t[50]);
  assign t[49] = ~(t[90] | t[92]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[90]);
  assign t[51] = t[1] ? t[52] : t[95];
  assign t[52] = x[6] ? t[54] : t[53];
  assign t[53] = x[7] ? t[56] : t[55];
  assign t[54] = t[57] ^ x[60];
  assign t[55] = t[58] ^ t[59];
  assign t[56] = ~(t[96] ^ t[60]);
  assign t[57] = x[62] ^ x[63];
  assign t[58] = t[20] ? x[63] : x[62];
  assign t[59] = ~(t[97] ^ t[61]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[98] ^ t[99]);
  assign t[61] = ~(t[100] ^ t[101]);
  assign t[62] = t[1] ? t[63] : t[102];
  assign t[63] = x[6] ? t[65] : t[64];
  assign t[64] = x[7] ? t[67] : t[66];
  assign t[65] = t[68] ^ x[70];
  assign t[66] = t[69] ^ t[70];
  assign t[67] = ~(t[103] ^ t[71]);
  assign t[68] = x[72] ^ x[73];
  assign t[69] = t[20] ? x[73] : x[72];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104] ^ t[72]);
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = ~(t[107] ^ t[108]);
  assign t[73] = t[1] ? t[74] : t[109];
  assign t[74] = x[6] ? t[76] : t[75];
  assign t[75] = x[7] ? t[78] : t[77];
  assign t[76] = t[79] ^ x[80];
  assign t[77] = t[80] ^ t[81];
  assign t[78] = ~(t[110] ^ t[82]);
  assign t[79] = x[82] ^ x[83];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[20] ? x[83] : x[82];
  assign t[81] = ~(t[111] ^ t[83]);
  assign t[82] = ~(t[112] ^ t[113]);
  assign t[83] = ~(t[114] ^ t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[85] ^ t[14]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[51] & ~t[62] & ~t[73]) | (~t[0] & t[51] & ~t[62] & ~t[73]) | (~t[0] & ~t[51] & t[62] & ~t[73]) | (~t[0] & ~t[51] & ~t[62] & t[73]) | (t[0] & t[51] & t[62] & ~t[73]) | (t[0] & t[51] & ~t[62] & t[73]) | (t[0] & ~t[51] & t[62] & t[73]) | (~t[0] & t[51] & t[62] & t[73]);
endmodule

module R2ind156(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[2]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[11]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[19]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[25]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[49]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[1]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[10]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[18]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[48]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[54]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [58:0] x;
 output y;

 wire [127:0] t;
  assign t[0] = t[1] ? t[2] : t[51];
  assign t[100] = t[122] ^ x[45];
  assign t[101] = t[123] ^ x[46];
  assign t[102] = t[124] ^ x[51];
  assign t[103] = t[125] ^ x[52];
  assign t[104] = t[126] ^ x[57];
  assign t[105] = t[127] ^ x[58];
  assign t[106] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[107] = (x[0]);
  assign t[108] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[109] = (x[9]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[111] = (x[17]);
  assign t[112] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[113] = (x[23]);
  assign t[114] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[115] = (x[29]);
  assign t[116] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[117] = (x[35]);
  assign t[118] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[119] = (x[38]);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[121] = (x[41]);
  assign t[122] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[44]);
  assign t[124] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[125] = (x[47]);
  assign t[126] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[127] = (x[53]);
  assign t[12] = ~(t[53] ^ t[17]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[54] ^ t[55]);
  assign t[15] = ~(t[56] & t[57]);
  assign t[16] = ~(t[58] & t[59]);
  assign t[17] = ~(t[60] ^ t[61]);
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] & t[27]);
  assign t[23] = ~(t[58]);
  assign t[24] = ~(t[28] & t[29]);
  assign t[25] = t[30] | t[31];
  assign t[26] = t[59] & t[32];
  assign t[27] = t[33] | t[34];
  assign t[28] = ~(t[32] & t[35]);
  assign t[29] = ~(t[36] & t[37]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[38] | t[39]);
  assign t[31] = ~(t[38] | t[40]);
  assign t[32] = ~(t[41] | t[56]);
  assign t[33] = ~(x[7] | t[57]);
  assign t[34] = x[7] & t[57];
  assign t[35] = ~(t[42] & t[43]);
  assign t[36] = ~(t[57] | t[44]);
  assign t[37] = t[38] & t[56];
  assign t[38] = ~(t[41]);
  assign t[39] = t[56] ? t[42] : t[45];
  assign t[3] = ~(t[6]);
  assign t[40] = t[56] ? t[47] : t[46];
  assign t[41] = ~(t[58]);
  assign t[42] = ~(t[59] & t[48]);
  assign t[43] = ~(x[7] & t[36]);
  assign t[44] = ~(t[59]);
  assign t[45] = ~(x[7] & t[49]);
  assign t[46] = ~(t[34] & t[44]);
  assign t[47] = ~(t[33] & t[59]);
  assign t[48] = ~(x[7] | t[50]);
  assign t[49] = ~(t[57] | t[59]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[57]);
  assign t[51] = (t[62]);
  assign t[52] = (t[63]);
  assign t[53] = (t[64]);
  assign t[54] = (t[65]);
  assign t[55] = (t[66]);
  assign t[56] = (t[67]);
  assign t[57] = (t[68]);
  assign t[58] = (t[69]);
  assign t[59] = (t[70]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = t[73] ^ x[5];
  assign t[63] = t[74] ^ x[14];
  assign t[64] = t[75] ^ x[22];
  assign t[65] = t[76] ^ x[28];
  assign t[66] = t[77] ^ x[34];
  assign t[67] = t[78] ^ x[37];
  assign t[68] = t[79] ^ x[40];
  assign t[69] = t[80] ^ x[43];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[81] ^ x[46];
  assign t[71] = t[82] ^ x[52];
  assign t[72] = t[83] ^ x[58];
  assign t[73] = (~t[84] & t[85]);
  assign t[74] = (~t[86] & t[87]);
  assign t[75] = (~t[88] & t[89]);
  assign t[76] = (~t[90] & t[91]);
  assign t[77] = (~t[92] & t[93]);
  assign t[78] = (~t[94] & t[95]);
  assign t[79] = (~t[96] & t[97]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[98] & t[99]);
  assign t[81] = (~t[100] & t[101]);
  assign t[82] = (~t[102] & t[103]);
  assign t[83] = (~t[104] & t[105]);
  assign t[84] = t[106] ^ x[4];
  assign t[85] = t[107] ^ x[5];
  assign t[86] = t[108] ^ x[13];
  assign t[87] = t[109] ^ x[14];
  assign t[88] = t[110] ^ x[21];
  assign t[89] = t[111] ^ x[22];
  assign t[8] = ~(t[52] ^ t[14]);
  assign t[90] = t[112] ^ x[27];
  assign t[91] = t[113] ^ x[28];
  assign t[92] = t[114] ^ x[33];
  assign t[93] = t[115] ^ x[34];
  assign t[94] = t[116] ^ x[36];
  assign t[95] = t[117] ^ x[37];
  assign t[96] = t[118] ^ x[39];
  assign t[97] = t[119] ^ x[40];
  assign t[98] = t[120] ^ x[42];
  assign t[99] = t[121] ^ x[43];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [88:0] x;
 output y;

 wire [265:0] t;
  assign t[0] = t[1] ? t[2] : t[84];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = t[148] ^ x[5];
  assign t[117] = t[149] ^ x[14];
  assign t[118] = t[150] ^ x[22];
  assign t[119] = t[151] ^ x[28];
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[34];
  assign t[121] = t[153] ^ x[37];
  assign t[122] = t[154] ^ x[40];
  assign t[123] = t[155] ^ x[43];
  assign t[124] = t[156] ^ x[46];
  assign t[125] = t[157] ^ x[52];
  assign t[126] = t[158] ^ x[58];
  assign t[127] = t[159] ^ x[59];
  assign t[128] = t[160] ^ x[61];
  assign t[129] = t[161] ^ x[64];
  assign t[12] = ~(t[86] ^ t[17]);
  assign t[130] = t[162] ^ x[65];
  assign t[131] = t[163] ^ x[66];
  assign t[132] = t[164] ^ x[67];
  assign t[133] = t[165] ^ x[68];
  assign t[134] = t[166] ^ x[69];
  assign t[135] = t[167] ^ x[71];
  assign t[136] = t[168] ^ x[74];
  assign t[137] = t[169] ^ x[75];
  assign t[138] = t[170] ^ x[76];
  assign t[139] = t[171] ^ x[77];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[78];
  assign t[141] = t[173] ^ x[79];
  assign t[142] = t[174] ^ x[81];
  assign t[143] = t[175] ^ x[84];
  assign t[144] = t[176] ^ x[85];
  assign t[145] = t[177] ^ x[86];
  assign t[146] = t[178] ^ x[87];
  assign t[147] = t[179] ^ x[88];
  assign t[148] = (~t[180] & t[181]);
  assign t[149] = (~t[182] & t[183]);
  assign t[14] = ~(t[87] ^ t[88]);
  assign t[150] = (~t[184] & t[185]);
  assign t[151] = (~t[186] & t[187]);
  assign t[152] = (~t[188] & t[189]);
  assign t[153] = (~t[190] & t[191]);
  assign t[154] = (~t[192] & t[193]);
  assign t[155] = (~t[194] & t[195]);
  assign t[156] = (~t[196] & t[197]);
  assign t[157] = (~t[198] & t[199]);
  assign t[158] = (~t[200] & t[201]);
  assign t[159] = (~t[180] & t[202]);
  assign t[15] = ~(t[89] & t[90]);
  assign t[160] = (~t[182] & t[203]);
  assign t[161] = (~t[184] & t[204]);
  assign t[162] = (~t[188] & t[205]);
  assign t[163] = (~t[186] & t[206]);
  assign t[164] = (~t[200] & t[207]);
  assign t[165] = (~t[198] & t[208]);
  assign t[166] = (~t[180] & t[209]);
  assign t[167] = (~t[182] & t[210]);
  assign t[168] = (~t[184] & t[211]);
  assign t[169] = (~t[186] & t[212]);
  assign t[16] = ~(t[91] & t[92]);
  assign t[170] = (~t[188] & t[213]);
  assign t[171] = (~t[200] & t[214]);
  assign t[172] = (~t[198] & t[215]);
  assign t[173] = (~t[180] & t[216]);
  assign t[174] = (~t[182] & t[217]);
  assign t[175] = (~t[184] & t[218]);
  assign t[176] = (~t[186] & t[219]);
  assign t[177] = (~t[188] & t[220]);
  assign t[178] = (~t[200] & t[221]);
  assign t[179] = (~t[198] & t[222]);
  assign t[17] = ~(t[93] ^ t[94]);
  assign t[180] = t[223] ^ x[4];
  assign t[181] = t[224] ^ x[5];
  assign t[182] = t[225] ^ x[13];
  assign t[183] = t[226] ^ x[14];
  assign t[184] = t[227] ^ x[21];
  assign t[185] = t[228] ^ x[22];
  assign t[186] = t[229] ^ x[27];
  assign t[187] = t[230] ^ x[28];
  assign t[188] = t[231] ^ x[33];
  assign t[189] = t[232] ^ x[34];
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[190] = t[233] ^ x[36];
  assign t[191] = t[234] ^ x[37];
  assign t[192] = t[235] ^ x[39];
  assign t[193] = t[236] ^ x[40];
  assign t[194] = t[237] ^ x[42];
  assign t[195] = t[238] ^ x[43];
  assign t[196] = t[239] ^ x[45];
  assign t[197] = t[240] ^ x[46];
  assign t[198] = t[241] ^ x[51];
  assign t[199] = t[242] ^ x[52];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[57];
  assign t[201] = t[244] ^ x[58];
  assign t[202] = t[245] ^ x[59];
  assign t[203] = t[246] ^ x[61];
  assign t[204] = t[247] ^ x[64];
  assign t[205] = t[248] ^ x[65];
  assign t[206] = t[249] ^ x[66];
  assign t[207] = t[250] ^ x[67];
  assign t[208] = t[251] ^ x[68];
  assign t[209] = t[252] ^ x[69];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[71];
  assign t[211] = t[254] ^ x[74];
  assign t[212] = t[255] ^ x[75];
  assign t[213] = t[256] ^ x[76];
  assign t[214] = t[257] ^ x[77];
  assign t[215] = t[258] ^ x[78];
  assign t[216] = t[259] ^ x[79];
  assign t[217] = t[260] ^ x[81];
  assign t[218] = t[261] ^ x[84];
  assign t[219] = t[262] ^ x[85];
  assign t[21] = ~(t[24]);
  assign t[220] = t[263] ^ x[86];
  assign t[221] = t[264] ^ x[87];
  assign t[222] = t[265] ^ x[88];
  assign t[223] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[224] = (x[0]);
  assign t[225] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[226] = (x[9]);
  assign t[227] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[228] = (x[17]);
  assign t[229] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[22] = ~(t[25] | t[26]);
  assign t[230] = (x[23]);
  assign t[231] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[232] = (x[29]);
  assign t[233] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[234] = (x[35]);
  assign t[235] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[236] = (x[38]);
  assign t[237] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[238] = (x[41]);
  assign t[239] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[23] = ~(t[91]);
  assign t[240] = (x[44]);
  assign t[241] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[242] = (x[47]);
  assign t[243] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[244] = (x[53]);
  assign t[245] = (x[1]);
  assign t[246] = (x[10]);
  assign t[247] = (x[18]);
  assign t[248] = (x[30]);
  assign t[249] = (x[24]);
  assign t[24] = ~(t[27] | t[28]);
  assign t[250] = (x[54]);
  assign t[251] = (x[48]);
  assign t[252] = (x[2]);
  assign t[253] = (x[11]);
  assign t[254] = (x[19]);
  assign t[255] = (x[25]);
  assign t[256] = (x[31]);
  assign t[257] = (x[55]);
  assign t[258] = (x[49]);
  assign t[259] = (x[3]);
  assign t[25] = ~(t[29]);
  assign t[260] = (x[12]);
  assign t[261] = (x[20]);
  assign t[262] = (x[26]);
  assign t[263] = (x[32]);
  assign t[264] = (x[56]);
  assign t[265] = (x[50]);
  assign t[26] = ~(t[27] | t[30]);
  assign t[27] = ~(t[31]);
  assign t[28] = t[89] ? t[33] : t[32];
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[89] ? t[37] : t[36];
  assign t[31] = ~(t[91]);
  assign t[32] = ~(t[38] & t[39]);
  assign t[33] = ~(t[40] & t[92]);
  assign t[34] = ~(t[27] | t[41]);
  assign t[35] = ~(t[27] | t[42]);
  assign t[36] = ~(x[7] & t[43]);
  assign t[37] = ~(t[92] & t[44]);
  assign t[38] = ~(x[7] | t[90]);
  assign t[39] = ~(t[92]);
  assign t[3] = ~(t[6]);
  assign t[40] = x[7] & t[90];
  assign t[41] = t[89] ? t[46] : t[45];
  assign t[42] = t[89] ? t[48] : t[47];
  assign t[43] = ~(t[90] | t[92]);
  assign t[44] = ~(x[7] | t[49]);
  assign t[45] = ~(t[44] & t[39]);
  assign t[46] = ~(x[7] & t[50]);
  assign t[47] = ~(t[38] & t[92]);
  assign t[48] = ~(t[40] & t[39]);
  assign t[49] = ~(t[90]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[90] | t[39]);
  assign t[51] = t[6] ? t[52] : t[95];
  assign t[52] = x[6] ? t[54] : t[53];
  assign t[53] = x[7] ? t[56] : t[55];
  assign t[54] = t[57] ^ x[60];
  assign t[55] = t[58] ^ t[59];
  assign t[56] = ~(t[96] ^ t[60]);
  assign t[57] = x[62] ^ x[63];
  assign t[58] = t[20] ? x[63] : x[62];
  assign t[59] = ~(t[97] ^ t[61]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[98] ^ t[99]);
  assign t[61] = ~(t[100] ^ t[101]);
  assign t[62] = t[6] ? t[63] : t[102];
  assign t[63] = x[6] ? t[65] : t[64];
  assign t[64] = x[7] ? t[67] : t[66];
  assign t[65] = t[68] ^ x[70];
  assign t[66] = t[69] ^ t[70];
  assign t[67] = ~(t[103] ^ t[71]);
  assign t[68] = x[72] ^ x[73];
  assign t[69] = t[20] ? x[73] : x[72];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104] ^ t[72]);
  assign t[71] = ~(t[105] ^ t[106]);
  assign t[72] = ~(t[107] ^ t[108]);
  assign t[73] = t[1] ? t[74] : t[109];
  assign t[74] = x[6] ? t[76] : t[75];
  assign t[75] = x[7] ? t[78] : t[77];
  assign t[76] = t[79] ^ x[80];
  assign t[77] = t[80] ^ t[81];
  assign t[78] = ~(t[110] ^ t[82]);
  assign t[79] = x[82] ^ x[83];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[20] ? x[83] : x[82];
  assign t[81] = ~(t[111] ^ t[83]);
  assign t[82] = ~(t[112] ^ t[113]);
  assign t[83] = ~(t[114] ^ t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[85] ^ t[14]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[51] & ~t[62] & ~t[73]) | (~t[0] & t[51] & ~t[62] & ~t[73]) | (~t[0] & ~t[51] & t[62] & ~t[73]) | (~t[0] & ~t[51] & ~t[62] & t[73]) | (t[0] & t[51] & t[62] & ~t[73]) | (t[0] & t[51] & ~t[62] & t[73]) | (t[0] & ~t[51] & t[62] & t[73]) | (~t[0] & t[51] & t[62] & t[73]);
endmodule

module R2ind161(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [58:0] x;
 output y;

 wire [94:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[23] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[15] ? x[28] : x[27];
  assign t[13] = ~(t[24] ^ t[16]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[15] = ~(t[17]);
  assign t[16] = ~(t[27] ^ t[28]);
  assign t[17] = ~(t[21]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = t[40] ^ x[5];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[11];
  assign t[31] = t[42] ^ x[14];
  assign t[32] = t[43] ^ x[17];
  assign t[33] = t[44] ^ x[20];
  assign t[34] = t[45] ^ x[26];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[40];
  assign t[37] = t[48] ^ x[46];
  assign t[38] = t[49] ^ x[52];
  assign t[39] = t[50] ^ x[58];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[51] & t[52]);
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[6]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = t[73] ^ x[4];
  assign t[52] = t[74] ^ x[5];
  assign t[53] = t[75] ^ x[10];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[16];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[19];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[25];
  assign t[62] = t[84] ^ x[26];
  assign t[63] = t[85] ^ x[33];
  assign t[64] = t[86] ^ x[34];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[45];
  assign t[68] = t[90] ^ x[46];
  assign t[69] = t[91] ^ x[51];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[52];
  assign t[71] = t[93] ^ x[57];
  assign t[72] = t[94] ^ x[58];
  assign t[73] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[74] = (x[2]);
  assign t[75] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[9]);
  assign t[77] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[12]);
  assign t[79] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[15]);
  assign t[81] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[18]);
  assign t[83] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[84] = (x[23]);
  assign t[85] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[86] = (x[31]);
  assign t[87] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[88] = (x[37]);
  assign t[89] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[43]);
  assign t[91] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[92] = (x[49]);
  assign t[93] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[94] = (x[55]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [58:0] x;
 output y;

 wire [94:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[23] ^ t[14]);
  assign t[11] = x[27] ^ x[28];
  assign t[12] = t[15] ? x[28] : x[27];
  assign t[13] = ~(t[24] ^ t[16]);
  assign t[14] = ~(t[25] ^ t[26]);
  assign t[15] = ~(t[17]);
  assign t[16] = ~(t[27] ^ t[28]);
  assign t[17] = ~(t[21]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = t[40] ^ x[5];
  assign t[2] = x[6] ? t[6] : t[5];
  assign t[30] = t[41] ^ x[11];
  assign t[31] = t[42] ^ x[14];
  assign t[32] = t[43] ^ x[17];
  assign t[33] = t[44] ^ x[20];
  assign t[34] = t[45] ^ x[26];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[40];
  assign t[37] = t[48] ^ x[46];
  assign t[38] = t[49] ^ x[52];
  assign t[39] = t[50] ^ x[58];
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (~t[51] & t[52]);
  assign t[41] = (~t[53] & t[54]);
  assign t[42] = (~t[55] & t[56]);
  assign t[43] = (~t[57] & t[58]);
  assign t[44] = (~t[59] & t[60]);
  assign t[45] = (~t[61] & t[62]);
  assign t[46] = (~t[63] & t[64]);
  assign t[47] = (~t[65] & t[66]);
  assign t[48] = (~t[67] & t[68]);
  assign t[49] = (~t[69] & t[70]);
  assign t[4] = ~(x[6]);
  assign t[50] = (~t[71] & t[72]);
  assign t[51] = t[73] ^ x[4];
  assign t[52] = t[74] ^ x[5];
  assign t[53] = t[75] ^ x[10];
  assign t[54] = t[76] ^ x[11];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[16];
  assign t[58] = t[80] ^ x[17];
  assign t[59] = t[81] ^ x[19];
  assign t[5] = x[7] ? t[10] : t[9];
  assign t[60] = t[82] ^ x[20];
  assign t[61] = t[83] ^ x[25];
  assign t[62] = t[84] ^ x[26];
  assign t[63] = t[85] ^ x[33];
  assign t[64] = t[86] ^ x[34];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[45];
  assign t[68] = t[90] ^ x[46];
  assign t[69] = t[91] ^ x[51];
  assign t[6] = t[11] ^ x[8];
  assign t[70] = t[92] ^ x[52];
  assign t[71] = t[93] ^ x[57];
  assign t[72] = t[94] ^ x[58];
  assign t[73] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[74] = (x[1]);
  assign t[75] = (x[9] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[9] & 1'b0 & ~1'b0 & ~1'b0) | (~x[9] & ~1'b0 & 1'b0 & ~1'b0) | (~x[9] & ~1'b0 & ~1'b0 & 1'b0) | (x[9] & 1'b0 & 1'b0 & ~1'b0) | (x[9] & 1'b0 & ~1'b0 & 1'b0) | (x[9] & ~1'b0 & 1'b0 & 1'b0) | (~x[9] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[9]);
  assign t[77] = (x[12] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[12] & 1'b0 & ~1'b0 & ~1'b0) | (~x[12] & ~1'b0 & 1'b0 & ~1'b0) | (~x[12] & ~1'b0 & ~1'b0 & 1'b0) | (x[12] & 1'b0 & 1'b0 & ~1'b0) | (x[12] & 1'b0 & ~1'b0 & 1'b0) | (x[12] & ~1'b0 & 1'b0 & 1'b0) | (~x[12] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[12]);
  assign t[79] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[19] & t[20]);
  assign t[80] = (x[15]);
  assign t[81] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[18]);
  assign t[83] = (x[21] & ~x[22] & ~x[23] & ~x[24]) | (~x[21] & x[22] & ~x[23] & ~x[24]) | (~x[21] & ~x[22] & x[23] & ~x[24]) | (~x[21] & ~x[22] & ~x[23] & x[24]) | (x[21] & x[22] & x[23] & ~x[24]) | (x[21] & x[22] & ~x[23] & x[24]) | (x[21] & ~x[22] & x[23] & x[24]) | (~x[21] & x[22] & x[23] & x[24]);
  assign t[84] = (x[22]);
  assign t[85] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[86] = (x[30]);
  assign t[87] = (x[35] & ~x[36] & ~x[37] & ~x[38]) | (~x[35] & x[36] & ~x[37] & ~x[38]) | (~x[35] & ~x[36] & x[37] & ~x[38]) | (~x[35] & ~x[36] & ~x[37] & x[38]) | (x[35] & x[36] & x[37] & ~x[38]) | (x[35] & x[36] & ~x[37] & x[38]) | (x[35] & ~x[36] & x[37] & x[38]) | (~x[35] & x[36] & x[37] & x[38]);
  assign t[88] = (x[36]);
  assign t[89] = (x[41] & ~x[42] & ~x[43] & ~x[44]) | (~x[41] & x[42] & ~x[43] & ~x[44]) | (~x[41] & ~x[42] & x[43] & ~x[44]) | (~x[41] & ~x[42] & ~x[43] & x[44]) | (x[41] & x[42] & x[43] & ~x[44]) | (x[41] & x[42] & ~x[43] & x[44]) | (x[41] & ~x[42] & x[43] & x[44]) | (~x[41] & x[42] & x[43] & x[44]);
  assign t[8] = ~(t[21] & t[22]);
  assign t[90] = (x[42]);
  assign t[91] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[92] = (x[48]);
  assign t[93] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[94] = (x[54]);
  assign t[9] = t[12] ^ t[13];
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [58:0] x;
 output y;

 wire [127:0] t;
  assign t[0] = t[1] ? t[2] : t[51];
  assign t[100] = t[122] ^ x[45];
  assign t[101] = t[123] ^ x[46];
  assign t[102] = t[124] ^ x[51];
  assign t[103] = t[125] ^ x[52];
  assign t[104] = t[126] ^ x[57];
  assign t[105] = t[127] ^ x[58];
  assign t[106] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[107] = (x[0]);
  assign t[108] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[109] = (x[9]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[111] = (x[17]);
  assign t[112] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[113] = (x[23]);
  assign t[114] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[115] = (x[29]);
  assign t[116] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[117] = (x[35]);
  assign t[118] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[119] = (x[38]);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[121] = (x[41]);
  assign t[122] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[123] = (x[44]);
  assign t[124] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[125] = (x[47]);
  assign t[126] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[127] = (x[53]);
  assign t[12] = ~(t[53] ^ t[17]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[54] ^ t[55]);
  assign t[15] = ~(t[56] & t[57]);
  assign t[16] = ~(t[58] & t[59]);
  assign t[17] = ~(t[60] ^ t[61]);
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[25] | t[26]);
  assign t[23] = ~(t[58]);
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29]);
  assign t[26] = ~(t[27] | t[30]);
  assign t[27] = ~(t[31]);
  assign t[28] = t[56] ? t[33] : t[32];
  assign t[29] = ~(t[34] | t[35]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[56] ? t[37] : t[36];
  assign t[31] = ~(t[58]);
  assign t[32] = ~(t[38] & t[39]);
  assign t[33] = ~(t[40] & t[59]);
  assign t[34] = ~(t[27] | t[41]);
  assign t[35] = ~(t[27] | t[42]);
  assign t[36] = ~(x[7] & t[43]);
  assign t[37] = ~(t[59] & t[44]);
  assign t[38] = ~(x[7] | t[57]);
  assign t[39] = ~(t[59]);
  assign t[3] = ~(t[6]);
  assign t[40] = x[7] & t[57];
  assign t[41] = t[56] ? t[46] : t[45];
  assign t[42] = t[56] ? t[48] : t[47];
  assign t[43] = ~(t[57] | t[59]);
  assign t[44] = ~(x[7] | t[49]);
  assign t[45] = ~(t[44] & t[39]);
  assign t[46] = ~(x[7] & t[50]);
  assign t[47] = ~(t[38] & t[59]);
  assign t[48] = ~(t[40] & t[39]);
  assign t[49] = ~(t[57]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[57] | t[39]);
  assign t[51] = (t[62]);
  assign t[52] = (t[63]);
  assign t[53] = (t[64]);
  assign t[54] = (t[65]);
  assign t[55] = (t[66]);
  assign t[56] = (t[67]);
  assign t[57] = (t[68]);
  assign t[58] = (t[69]);
  assign t[59] = (t[70]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = t[73] ^ x[5];
  assign t[63] = t[74] ^ x[14];
  assign t[64] = t[75] ^ x[22];
  assign t[65] = t[76] ^ x[28];
  assign t[66] = t[77] ^ x[34];
  assign t[67] = t[78] ^ x[37];
  assign t[68] = t[79] ^ x[40];
  assign t[69] = t[80] ^ x[43];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[81] ^ x[46];
  assign t[71] = t[82] ^ x[52];
  assign t[72] = t[83] ^ x[58];
  assign t[73] = (~t[84] & t[85]);
  assign t[74] = (~t[86] & t[87]);
  assign t[75] = (~t[88] & t[89]);
  assign t[76] = (~t[90] & t[91]);
  assign t[77] = (~t[92] & t[93]);
  assign t[78] = (~t[94] & t[95]);
  assign t[79] = (~t[96] & t[97]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[98] & t[99]);
  assign t[81] = (~t[100] & t[101]);
  assign t[82] = (~t[102] & t[103]);
  assign t[83] = (~t[104] & t[105]);
  assign t[84] = t[106] ^ x[4];
  assign t[85] = t[107] ^ x[5];
  assign t[86] = t[108] ^ x[13];
  assign t[87] = t[109] ^ x[14];
  assign t[88] = t[110] ^ x[21];
  assign t[89] = t[111] ^ x[22];
  assign t[8] = ~(t[52] ^ t[14]);
  assign t[90] = t[112] ^ x[27];
  assign t[91] = t[113] ^ x[28];
  assign t[92] = t[114] ^ x[33];
  assign t[93] = t[115] ^ x[34];
  assign t[94] = t[116] ^ x[36];
  assign t[95] = t[117] ^ x[37];
  assign t[96] = t[118] ^ x[39];
  assign t[97] = t[119] ^ x[40];
  assign t[98] = t[120] ^ x[42];
  assign t[99] = t[121] ^ x[43];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [70:0] x;
 output y;

 wire [212:0] t;
  assign t[0] = t[1] ? t[2] : t[75];
  assign t[100] = t[124] ^ x[14];
  assign t[101] = t[125] ^ x[22];
  assign t[102] = t[126] ^ x[28];
  assign t[103] = t[127] ^ x[34];
  assign t[104] = t[128] ^ x[37];
  assign t[105] = t[129] ^ x[40];
  assign t[106] = t[130] ^ x[43];
  assign t[107] = t[131] ^ x[46];
  assign t[108] = t[132] ^ x[47];
  assign t[109] = t[133] ^ x[49];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[134] ^ x[52];
  assign t[111] = t[135] ^ x[53];
  assign t[112] = t[136] ^ x[54];
  assign t[113] = t[137] ^ x[55];
  assign t[114] = t[138] ^ x[57];
  assign t[115] = t[139] ^ x[60];
  assign t[116] = t[140] ^ x[61];
  assign t[117] = t[141] ^ x[62];
  assign t[118] = t[142] ^ x[63];
  assign t[119] = t[143] ^ x[65];
  assign t[11] = ~(x[6]);
  assign t[120] = t[144] ^ x[68];
  assign t[121] = t[145] ^ x[69];
  assign t[122] = t[146] ^ x[70];
  assign t[123] = (~t[147] & t[148]);
  assign t[124] = (~t[149] & t[150]);
  assign t[125] = (~t[151] & t[152]);
  assign t[126] = (~t[153] & t[154]);
  assign t[127] = (~t[155] & t[156]);
  assign t[128] = (~t[157] & t[158]);
  assign t[129] = (~t[159] & t[160]);
  assign t[12] = ~(t[77] ^ t[14]);
  assign t[130] = (~t[161] & t[162]);
  assign t[131] = (~t[163] & t[164]);
  assign t[132] = (~t[147] & t[165]);
  assign t[133] = (~t[149] & t[166]);
  assign t[134] = (~t[151] & t[167]);
  assign t[135] = (~t[155] & t[168]);
  assign t[136] = (~t[153] & t[169]);
  assign t[137] = (~t[147] & t[170]);
  assign t[138] = (~t[149] & t[171]);
  assign t[139] = (~t[151] & t[172]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[140] = (~t[155] & t[173]);
  assign t[141] = (~t[153] & t[174]);
  assign t[142] = (~t[147] & t[175]);
  assign t[143] = (~t[149] & t[176]);
  assign t[144] = (~t[151] & t[177]);
  assign t[145] = (~t[155] & t[178]);
  assign t[146] = (~t[153] & t[179]);
  assign t[147] = t[180] ^ x[4];
  assign t[148] = t[181] ^ x[5];
  assign t[149] = t[182] ^ x[13];
  assign t[14] = ~(t[78] ^ t[79]);
  assign t[150] = t[183] ^ x[14];
  assign t[151] = t[184] ^ x[21];
  assign t[152] = t[185] ^ x[22];
  assign t[153] = t[186] ^ x[27];
  assign t[154] = t[187] ^ x[28];
  assign t[155] = t[188] ^ x[33];
  assign t[156] = t[189] ^ x[34];
  assign t[157] = t[190] ^ x[36];
  assign t[158] = t[191] ^ x[37];
  assign t[159] = t[192] ^ x[39];
  assign t[15] = ~(t[80] & t[81]);
  assign t[160] = t[193] ^ x[40];
  assign t[161] = t[194] ^ x[42];
  assign t[162] = t[195] ^ x[43];
  assign t[163] = t[196] ^ x[45];
  assign t[164] = t[197] ^ x[46];
  assign t[165] = t[198] ^ x[47];
  assign t[166] = t[199] ^ x[49];
  assign t[167] = t[200] ^ x[52];
  assign t[168] = t[201] ^ x[53];
  assign t[169] = t[202] ^ x[54];
  assign t[16] = ~(t[82] & t[83]);
  assign t[170] = t[203] ^ x[55];
  assign t[171] = t[204] ^ x[57];
  assign t[172] = t[205] ^ x[60];
  assign t[173] = t[206] ^ x[61];
  assign t[174] = t[207] ^ x[62];
  assign t[175] = t[208] ^ x[63];
  assign t[176] = t[209] ^ x[65];
  assign t[177] = t[210] ^ x[68];
  assign t[178] = t[211] ^ x[69];
  assign t[179] = t[212] ^ x[70];
  assign t[17] = t[19] ? x[16] : x[15];
  assign t[180] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[181] = (x[0]);
  assign t[182] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[183] = (x[9]);
  assign t[184] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[185] = (x[17]);
  assign t[186] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[187] = (x[23]);
  assign t[188] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[189] = (x[29]);
  assign t[18] = t[20] | t[21];
  assign t[190] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[191] = (x[35]);
  assign t[192] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[193] = (x[38]);
  assign t[194] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[195] = (x[41]);
  assign t[196] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[197] = (x[44]);
  assign t[198] = (x[1]);
  assign t[199] = (x[10]);
  assign t[19] = ~(t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = (x[18]);
  assign t[201] = (x[30]);
  assign t[202] = (x[24]);
  assign t[203] = (x[2]);
  assign t[204] = (x[11]);
  assign t[205] = (x[19]);
  assign t[206] = (x[31]);
  assign t[207] = (x[25]);
  assign t[208] = (x[3]);
  assign t[209] = (x[12]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[210] = (x[20]);
  assign t[211] = (x[32]);
  assign t[212] = (x[26]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[82]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[29] & t[30]);
  assign t[25] = ~(t[31]);
  assign t[26] = t[80] ? t[33] : t[32];
  assign t[27] = ~(t[31] | t[34]);
  assign t[28] = ~(t[31] | t[35]);
  assign t[29] = ~(t[81] | t[36]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[25] & t[80];
  assign t[31] = ~(t[82]);
  assign t[32] = ~(x[7] & t[37]);
  assign t[33] = ~(t[83] & t[38]);
  assign t[34] = t[80] ? t[40] : t[39];
  assign t[35] = t[80] ? t[41] : t[32];
  assign t[36] = ~(t[83]);
  assign t[37] = ~(t[81] | t[83]);
  assign t[38] = ~(x[7] | t[42]);
  assign t[39] = ~(t[43] & t[36]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[44] & t[36]);
  assign t[41] = ~(t[38] & t[36]);
  assign t[42] = ~(t[81]);
  assign t[43] = ~(x[7] | t[81]);
  assign t[44] = x[7] & t[81];
  assign t[45] = t[1] ? t[46] : t[84];
  assign t[46] = x[6] ? t[48] : t[47];
  assign t[47] = x[7] ? t[50] : t[49];
  assign t[48] = t[51] ^ x[48];
  assign t[49] = t[52] ^ t[53];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(t[85] ^ t[54]);
  assign t[51] = x[50] ^ x[51];
  assign t[52] = t[19] ? x[51] : x[50];
  assign t[53] = ~(t[86] ^ t[54]);
  assign t[54] = ~(t[87] ^ t[88]);
  assign t[55] = t[1] ? t[56] : t[89];
  assign t[56] = x[6] ? t[58] : t[57];
  assign t[57] = x[7] ? t[60] : t[59];
  assign t[58] = t[61] ^ x[56];
  assign t[59] = t[62] ^ t[63];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[90] ^ t[64]);
  assign t[61] = x[58] ^ x[59];
  assign t[62] = t[19] ? x[59] : x[58];
  assign t[63] = ~(t[91] ^ t[64]);
  assign t[64] = ~(t[92] ^ t[93]);
  assign t[65] = t[1] ? t[66] : t[94];
  assign t[66] = x[6] ? t[68] : t[67];
  assign t[67] = x[7] ? t[70] : t[69];
  assign t[68] = t[71] ^ x[64];
  assign t[69] = t[72] ^ t[73];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[95] ^ t[74]);
  assign t[71] = x[66] ^ x[67];
  assign t[72] = t[19] ? x[67] : x[66];
  assign t[73] = ~(t[96] ^ t[74]);
  assign t[74] = ~(t[97] ^ t[98]);
  assign t[75] = (t[99]);
  assign t[76] = (t[100]);
  assign t[77] = (t[101]);
  assign t[78] = (t[102]);
  assign t[79] = (t[103]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (t[104]);
  assign t[81] = (t[105]);
  assign t[82] = (t[106]);
  assign t[83] = (t[107]);
  assign t[84] = (t[108]);
  assign t[85] = (t[109]);
  assign t[86] = (t[110]);
  assign t[87] = (t[111]);
  assign t[88] = (t[112]);
  assign t[89] = (t[113]);
  assign t[8] = ~(t[76] ^ t[14]);
  assign t[90] = (t[114]);
  assign t[91] = (t[115]);
  assign t[92] = (t[116]);
  assign t[93] = (t[117]);
  assign t[94] = (t[118]);
  assign t[95] = (t[119]);
  assign t[96] = (t[120]);
  assign t[97] = (t[121]);
  assign t[98] = (t[122]);
  assign t[99] = t[123] ^ x[5];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[45] & ~t[55] & ~t[65]) | (~t[0] & t[45] & ~t[55] & ~t[65]) | (~t[0] & ~t[45] & t[55] & ~t[65]) | (~t[0] & ~t[45] & ~t[55] & t[65]) | (t[0] & t[45] & t[55] & ~t[65]) | (t[0] & t[45] & ~t[55] & t[65]) | (t[0] & ~t[45] & t[55] & t[65]) | (~t[0] & t[45] & t[55] & t[65]);
endmodule

module R2ind166(x, y);
 input [46:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = t[1] ? t[2] : t[19];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[21] ^ t[14]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[26] & t[27]);
  assign t[17] = ~(t[18]);
  assign t[18] = ~(t[26]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = t[37] ^ x[5];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[39] ^ x[22];
  assign t[31] = t[40] ^ x[28];
  assign t[32] = t[41] ^ x[34];
  assign t[33] = t[42] ^ x[37];
  assign t[34] = t[43] ^ x[40];
  assign t[35] = t[44] ^ x[43];
  assign t[36] = t[45] ^ x[46];
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[48] & t[49]);
  assign t[39] = (~t[50] & t[51]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[52] & t[53]);
  assign t[41] = (~t[54] & t[55]);
  assign t[42] = (~t[56] & t[57]);
  assign t[43] = (~t[58] & t[59]);
  assign t[44] = (~t[60] & t[61]);
  assign t[45] = (~t[62] & t[63]);
  assign t[46] = t[64] ^ x[4];
  assign t[47] = t[65] ^ x[5];
  assign t[48] = t[66] ^ x[13];
  assign t[49] = t[67] ^ x[14];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[68] ^ x[21];
  assign t[51] = t[69] ^ x[22];
  assign t[52] = t[70] ^ x[27];
  assign t[53] = t[71] ^ x[28];
  assign t[54] = t[72] ^ x[33];
  assign t[55] = t[73] ^ x[34];
  assign t[56] = t[74] ^ x[36];
  assign t[57] = t[75] ^ x[37];
  assign t[58] = t[76] ^ x[39];
  assign t[59] = t[77] ^ x[40];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[78] ^ x[42];
  assign t[61] = t[79] ^ x[43];
  assign t[62] = t[80] ^ x[45];
  assign t[63] = t[81] ^ x[46];
  assign t[64] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[65] = (x[3]);
  assign t[66] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[67] = (x[12]);
  assign t[68] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[69] = (x[20]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[71] = (x[26]);
  assign t[72] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[73] = (x[32]);
  assign t[74] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[35]);
  assign t[76] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[38]);
  assign t[78] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[41]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[44]);
  assign t[8] = ~(t[20] ^ t[14]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [46:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = t[1] ? t[2] : t[19];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[21] ^ t[14]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[26] & t[27]);
  assign t[17] = ~(t[18]);
  assign t[18] = ~(t[26]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = t[37] ^ x[5];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[39] ^ x[22];
  assign t[31] = t[40] ^ x[28];
  assign t[32] = t[41] ^ x[34];
  assign t[33] = t[42] ^ x[37];
  assign t[34] = t[43] ^ x[40];
  assign t[35] = t[44] ^ x[43];
  assign t[36] = t[45] ^ x[46];
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[48] & t[49]);
  assign t[39] = (~t[50] & t[51]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[52] & t[53]);
  assign t[41] = (~t[54] & t[55]);
  assign t[42] = (~t[56] & t[57]);
  assign t[43] = (~t[58] & t[59]);
  assign t[44] = (~t[60] & t[61]);
  assign t[45] = (~t[62] & t[63]);
  assign t[46] = t[64] ^ x[4];
  assign t[47] = t[65] ^ x[5];
  assign t[48] = t[66] ^ x[13];
  assign t[49] = t[67] ^ x[14];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[68] ^ x[21];
  assign t[51] = t[69] ^ x[22];
  assign t[52] = t[70] ^ x[27];
  assign t[53] = t[71] ^ x[28];
  assign t[54] = t[72] ^ x[33];
  assign t[55] = t[73] ^ x[34];
  assign t[56] = t[74] ^ x[36];
  assign t[57] = t[75] ^ x[37];
  assign t[58] = t[76] ^ x[39];
  assign t[59] = t[77] ^ x[40];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[78] ^ x[42];
  assign t[61] = t[79] ^ x[43];
  assign t[62] = t[80] ^ x[45];
  assign t[63] = t[81] ^ x[46];
  assign t[64] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[65] = (x[2]);
  assign t[66] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[67] = (x[11]);
  assign t[68] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[69] = (x[19]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[71] = (x[25]);
  assign t[72] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[73] = (x[31]);
  assign t[74] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[35]);
  assign t[76] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[38]);
  assign t[78] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[41]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[44]);
  assign t[8] = ~(t[20] ^ t[14]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [46:0] x;
 output y;

 wire [81:0] t;
  assign t[0] = t[1] ? t[2] : t[19];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[21] ^ t[14]);
  assign t[14] = ~(t[22] ^ t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[26] & t[27]);
  assign t[17] = ~(t[18]);
  assign t[18] = ~(t[26]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = (t[33]);
  assign t[25] = (t[34]);
  assign t[26] = (t[35]);
  assign t[27] = (t[36]);
  assign t[28] = t[37] ^ x[5];
  assign t[29] = t[38] ^ x[14];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[39] ^ x[22];
  assign t[31] = t[40] ^ x[28];
  assign t[32] = t[41] ^ x[34];
  assign t[33] = t[42] ^ x[37];
  assign t[34] = t[43] ^ x[40];
  assign t[35] = t[44] ^ x[43];
  assign t[36] = t[45] ^ x[46];
  assign t[37] = (~t[46] & t[47]);
  assign t[38] = (~t[48] & t[49]);
  assign t[39] = (~t[50] & t[51]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[52] & t[53]);
  assign t[41] = (~t[54] & t[55]);
  assign t[42] = (~t[56] & t[57]);
  assign t[43] = (~t[58] & t[59]);
  assign t[44] = (~t[60] & t[61]);
  assign t[45] = (~t[62] & t[63]);
  assign t[46] = t[64] ^ x[4];
  assign t[47] = t[65] ^ x[5];
  assign t[48] = t[66] ^ x[13];
  assign t[49] = t[67] ^ x[14];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[68] ^ x[21];
  assign t[51] = t[69] ^ x[22];
  assign t[52] = t[70] ^ x[27];
  assign t[53] = t[71] ^ x[28];
  assign t[54] = t[72] ^ x[33];
  assign t[55] = t[73] ^ x[34];
  assign t[56] = t[74] ^ x[36];
  assign t[57] = t[75] ^ x[37];
  assign t[58] = t[76] ^ x[39];
  assign t[59] = t[77] ^ x[40];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[78] ^ x[42];
  assign t[61] = t[79] ^ x[43];
  assign t[62] = t[80] ^ x[45];
  assign t[63] = t[81] ^ x[46];
  assign t[64] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[65] = (x[1]);
  assign t[66] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[67] = (x[10]);
  assign t[68] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[69] = (x[18]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[71] = (x[24]);
  assign t[72] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[73] = (x[30]);
  assign t[74] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[35]);
  assign t[76] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[38]);
  assign t[78] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[41]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[44]);
  assign t[8] = ~(t[20] ^ t[14]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [46:0] x;
 output y;

 wire [107:0] t;
  assign t[0] = t[1] ? t[2] : t[45];
  assign t[100] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[101] = (x[35]);
  assign t[102] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[103] = (x[38]);
  assign t[104] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[105] = (x[41]);
  assign t[106] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[107] = (x[44]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = ~(t[47] ^ t[14]);
  assign t[13] = ~(t[17] ^ t[18]);
  assign t[14] = ~(t[48] ^ t[49]);
  assign t[15] = ~(t[50] & t[51]);
  assign t[16] = ~(t[52] & t[53]);
  assign t[17] = t[19] ? x[16] : x[15];
  assign t[18] = t[20] | t[21];
  assign t[19] = ~(t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23] & t[24]);
  assign t[21] = ~(t[25] | t[26]);
  assign t[22] = ~(t[52]);
  assign t[23] = ~(t[27] | t[28]);
  assign t[24] = ~(t[29] & t[30]);
  assign t[25] = ~(t[31]);
  assign t[26] = t[50] ? t[33] : t[32];
  assign t[27] = ~(t[31] | t[34]);
  assign t[28] = ~(t[31] | t[35]);
  assign t[29] = ~(t[51] | t[36]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[25] & t[50];
  assign t[31] = ~(t[52]);
  assign t[32] = ~(x[7] & t[37]);
  assign t[33] = ~(t[53] & t[38]);
  assign t[34] = t[50] ? t[40] : t[39];
  assign t[35] = t[50] ? t[41] : t[32];
  assign t[36] = ~(t[53]);
  assign t[37] = ~(t[51] | t[53]);
  assign t[38] = ~(x[7] | t[42]);
  assign t[39] = ~(t[43] & t[36]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[44] & t[36]);
  assign t[41] = ~(t[38] & t[36]);
  assign t[42] = ~(t[51]);
  assign t[43] = ~(x[7] | t[51]);
  assign t[44] = x[7] & t[51];
  assign t[45] = (t[54]);
  assign t[46] = (t[55]);
  assign t[47] = (t[56]);
  assign t[48] = (t[57]);
  assign t[49] = (t[58]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (t[59]);
  assign t[51] = (t[60]);
  assign t[52] = (t[61]);
  assign t[53] = (t[62]);
  assign t[54] = t[63] ^ x[5];
  assign t[55] = t[64] ^ x[14];
  assign t[56] = t[65] ^ x[22];
  assign t[57] = t[66] ^ x[28];
  assign t[58] = t[67] ^ x[34];
  assign t[59] = t[68] ^ x[37];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[69] ^ x[40];
  assign t[61] = t[70] ^ x[43];
  assign t[62] = t[71] ^ x[46];
  assign t[63] = (~t[72] & t[73]);
  assign t[64] = (~t[74] & t[75]);
  assign t[65] = (~t[76] & t[77]);
  assign t[66] = (~t[78] & t[79]);
  assign t[67] = (~t[80] & t[81]);
  assign t[68] = (~t[82] & t[83]);
  assign t[69] = (~t[84] & t[85]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (~t[86] & t[87]);
  assign t[71] = (~t[88] & t[89]);
  assign t[72] = t[90] ^ x[4];
  assign t[73] = t[91] ^ x[5];
  assign t[74] = t[92] ^ x[13];
  assign t[75] = t[93] ^ x[14];
  assign t[76] = t[94] ^ x[21];
  assign t[77] = t[95] ^ x[22];
  assign t[78] = t[96] ^ x[27];
  assign t[79] = t[97] ^ x[28];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[98] ^ x[33];
  assign t[81] = t[99] ^ x[34];
  assign t[82] = t[100] ^ x[36];
  assign t[83] = t[101] ^ x[37];
  assign t[84] = t[102] ^ x[39];
  assign t[85] = t[103] ^ x[40];
  assign t[86] = t[104] ^ x[42];
  assign t[87] = t[105] ^ x[43];
  assign t[88] = t[106] ^ x[45];
  assign t[89] = t[107] ^ x[46];
  assign t[8] = ~(t[46] ^ t[14]);
  assign t[90] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[91] = (x[0]);
  assign t[92] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[93] = (x[9]);
  assign t[94] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[95] = (x[17]);
  assign t[96] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[97] = (x[23]);
  assign t[98] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[99] = (x[29]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [88:0] x;
 output y;

 wire [275:0] t;
  assign t[0] = t[1] ? t[2] : t[94];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = (t[155]);
  assign t[124] = (t[156]);
  assign t[125] = (t[157]);
  assign t[126] = t[158] ^ x[5];
  assign t[127] = t[159] ^ x[14];
  assign t[128] = t[160] ^ x[22];
  assign t[129] = t[161] ^ x[28];
  assign t[12] = ~(t[96] ^ t[17]);
  assign t[130] = t[162] ^ x[34];
  assign t[131] = t[163] ^ x[37];
  assign t[132] = t[164] ^ x[40];
  assign t[133] = t[165] ^ x[43];
  assign t[134] = t[166] ^ x[46];
  assign t[135] = t[167] ^ x[52];
  assign t[136] = t[168] ^ x[58];
  assign t[137] = t[169] ^ x[59];
  assign t[138] = t[170] ^ x[61];
  assign t[139] = t[171] ^ x[64];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[65];
  assign t[141] = t[173] ^ x[66];
  assign t[142] = t[174] ^ x[67];
  assign t[143] = t[175] ^ x[68];
  assign t[144] = t[176] ^ x[69];
  assign t[145] = t[177] ^ x[71];
  assign t[146] = t[178] ^ x[74];
  assign t[147] = t[179] ^ x[75];
  assign t[148] = t[180] ^ x[76];
  assign t[149] = t[181] ^ x[77];
  assign t[14] = ~(t[97] ^ t[98]);
  assign t[150] = t[182] ^ x[78];
  assign t[151] = t[183] ^ x[79];
  assign t[152] = t[184] ^ x[81];
  assign t[153] = t[185] ^ x[84];
  assign t[154] = t[186] ^ x[85];
  assign t[155] = t[187] ^ x[86];
  assign t[156] = t[188] ^ x[87];
  assign t[157] = t[189] ^ x[88];
  assign t[158] = (~t[190] & t[191]);
  assign t[159] = (~t[192] & t[193]);
  assign t[15] = ~(t[99] & t[100]);
  assign t[160] = (~t[194] & t[195]);
  assign t[161] = (~t[196] & t[197]);
  assign t[162] = (~t[198] & t[199]);
  assign t[163] = (~t[200] & t[201]);
  assign t[164] = (~t[202] & t[203]);
  assign t[165] = (~t[204] & t[205]);
  assign t[166] = (~t[206] & t[207]);
  assign t[167] = (~t[208] & t[209]);
  assign t[168] = (~t[210] & t[211]);
  assign t[169] = (~t[190] & t[212]);
  assign t[16] = ~(t[101] & t[102]);
  assign t[170] = (~t[192] & t[213]);
  assign t[171] = (~t[194] & t[214]);
  assign t[172] = (~t[198] & t[215]);
  assign t[173] = (~t[196] & t[216]);
  assign t[174] = (~t[210] & t[217]);
  assign t[175] = (~t[208] & t[218]);
  assign t[176] = (~t[190] & t[219]);
  assign t[177] = (~t[192] & t[220]);
  assign t[178] = (~t[194] & t[221]);
  assign t[179] = (~t[198] & t[222]);
  assign t[17] = ~(t[103] ^ t[104]);
  assign t[180] = (~t[196] & t[223]);
  assign t[181] = (~t[208] & t[224]);
  assign t[182] = (~t[210] & t[225]);
  assign t[183] = (~t[190] & t[226]);
  assign t[184] = (~t[192] & t[227]);
  assign t[185] = (~t[194] & t[228]);
  assign t[186] = (~t[198] & t[229]);
  assign t[187] = (~t[196] & t[230]);
  assign t[188] = (~t[208] & t[231]);
  assign t[189] = (~t[210] & t[232]);
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[190] = t[233] ^ x[4];
  assign t[191] = t[234] ^ x[5];
  assign t[192] = t[235] ^ x[13];
  assign t[193] = t[236] ^ x[14];
  assign t[194] = t[237] ^ x[21];
  assign t[195] = t[238] ^ x[22];
  assign t[196] = t[239] ^ x[27];
  assign t[197] = t[240] ^ x[28];
  assign t[198] = t[241] ^ x[33];
  assign t[199] = t[242] ^ x[34];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[36];
  assign t[201] = t[244] ^ x[37];
  assign t[202] = t[245] ^ x[39];
  assign t[203] = t[246] ^ x[40];
  assign t[204] = t[247] ^ x[42];
  assign t[205] = t[248] ^ x[43];
  assign t[206] = t[249] ^ x[45];
  assign t[207] = t[250] ^ x[46];
  assign t[208] = t[251] ^ x[51];
  assign t[209] = t[252] ^ x[52];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[57];
  assign t[211] = t[254] ^ x[58];
  assign t[212] = t[255] ^ x[59];
  assign t[213] = t[256] ^ x[61];
  assign t[214] = t[257] ^ x[64];
  assign t[215] = t[258] ^ x[65];
  assign t[216] = t[259] ^ x[66];
  assign t[217] = t[260] ^ x[67];
  assign t[218] = t[261] ^ x[68];
  assign t[219] = t[262] ^ x[69];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[71];
  assign t[221] = t[264] ^ x[74];
  assign t[222] = t[265] ^ x[75];
  assign t[223] = t[266] ^ x[76];
  assign t[224] = t[267] ^ x[77];
  assign t[225] = t[268] ^ x[78];
  assign t[226] = t[269] ^ x[79];
  assign t[227] = t[270] ^ x[81];
  assign t[228] = t[271] ^ x[84];
  assign t[229] = t[272] ^ x[85];
  assign t[22] = ~(t[26]);
  assign t[230] = t[273] ^ x[86];
  assign t[231] = t[274] ^ x[87];
  assign t[232] = t[275] ^ x[88];
  assign t[233] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[234] = (x[0]);
  assign t[235] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[236] = (x[9]);
  assign t[237] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[238] = (x[17]);
  assign t[239] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[23] = ~(t[101]);
  assign t[240] = (x[23]);
  assign t[241] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[242] = (x[29]);
  assign t[243] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[244] = (x[35]);
  assign t[245] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[246] = (x[38]);
  assign t[247] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[248] = (x[41]);
  assign t[249] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[24] = ~(t[27] | t[28]);
  assign t[250] = (x[44]);
  assign t[251] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[252] = (x[47]);
  assign t[253] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[254] = (x[53]);
  assign t[255] = (x[1]);
  assign t[256] = (x[10]);
  assign t[257] = (x[18]);
  assign t[258] = (x[30]);
  assign t[259] = (x[24]);
  assign t[25] = ~(t[29] & t[30]);
  assign t[260] = (x[54]);
  assign t[261] = (x[48]);
  assign t[262] = (x[2]);
  assign t[263] = (x[11]);
  assign t[264] = (x[19]);
  assign t[265] = (x[31]);
  assign t[266] = (x[25]);
  assign t[267] = (x[49]);
  assign t[268] = (x[55]);
  assign t[269] = (x[3]);
  assign t[26] = ~(t[27] | t[31]);
  assign t[270] = (x[12]);
  assign t[271] = (x[20]);
  assign t[272] = (x[32]);
  assign t[273] = (x[26]);
  assign t[274] = (x[50]);
  assign t[275] = (x[56]);
  assign t[27] = ~(t[32]);
  assign t[28] = t[99] ? t[34] : t[33];
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[37] | t[38]);
  assign t[31] = t[99] ? t[40] : t[39];
  assign t[32] = ~(t[101]);
  assign t[33] = ~(t[41] & t[42]);
  assign t[34] = ~(x[7] & t[43]);
  assign t[35] = ~(t[27] | t[44]);
  assign t[36] = ~(t[45] & t[46]);
  assign t[37] = ~(t[32] | t[47]);
  assign t[38] = ~(t[32] | t[48]);
  assign t[39] = ~(t[49] & t[102]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[50] & t[42]);
  assign t[41] = ~(x[7] | t[51]);
  assign t[42] = ~(t[102]);
  assign t[43] = ~(t[100] | t[42]);
  assign t[44] = t[99] ? t[39] : t[40];
  assign t[45] = ~(t[52] | t[53]);
  assign t[46] = ~(t[32] & t[54]);
  assign t[47] = t[99] ? t[55] : t[40];
  assign t[48] = t[99] ? t[33] : t[56];
  assign t[49] = x[7] & t[100];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(x[7] | t[100]);
  assign t[51] = ~(t[100]);
  assign t[52] = ~(t[32] | t[57]);
  assign t[53] = ~(t[27] | t[58]);
  assign t[54] = ~(t[56] & t[59]);
  assign t[55] = ~(t[49] & t[42]);
  assign t[56] = ~(x[7] & t[60]);
  assign t[57] = t[99] ? t[40] : t[55];
  assign t[58] = t[99] ? t[33] : t[34];
  assign t[59] = ~(t[102] & t[41]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[100] | t[102]);
  assign t[61] = t[1] ? t[62] : t[105];
  assign t[62] = x[6] ? t[64] : t[63];
  assign t[63] = x[7] ? t[66] : t[65];
  assign t[64] = t[67] ^ x[60];
  assign t[65] = t[68] ^ t[69];
  assign t[66] = ~(t[106] ^ t[70]);
  assign t[67] = x[62] ^ x[63];
  assign t[68] = t[20] ? x[63] : x[62];
  assign t[69] = ~(t[107] ^ t[71]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[108] ^ t[109]);
  assign t[71] = ~(t[110] ^ t[111]);
  assign t[72] = t[1] ? t[73] : t[112];
  assign t[73] = x[6] ? t[75] : t[74];
  assign t[74] = x[7] ? t[77] : t[76];
  assign t[75] = t[78] ^ x[70];
  assign t[76] = t[79] ^ t[80];
  assign t[77] = ~(t[113] ^ t[81]);
  assign t[78] = x[72] ^ x[73];
  assign t[79] = t[20] ? x[73] : x[72];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[114] ^ t[82]);
  assign t[81] = ~(t[115] ^ t[116]);
  assign t[82] = ~(t[117] ^ t[118]);
  assign t[83] = t[1] ? t[84] : t[119];
  assign t[84] = x[6] ? t[86] : t[85];
  assign t[85] = x[7] ? t[88] : t[87];
  assign t[86] = t[89] ^ x[80];
  assign t[87] = t[90] ^ t[91];
  assign t[88] = ~(t[120] ^ t[92]);
  assign t[89] = x[82] ^ x[83];
  assign t[8] = ~(t[95] ^ t[14]);
  assign t[90] = t[20] ? x[83] : x[82];
  assign t[91] = ~(t[121] ^ t[93]);
  assign t[92] = ~(t[122] ^ t[123]);
  assign t[93] = ~(t[124] ^ t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[61] & ~t[72] & ~t[83]) | (~t[0] & t[61] & ~t[72] & ~t[83]) | (~t[0] & ~t[61] & t[72] & ~t[83]) | (~t[0] & ~t[61] & ~t[72] & t[83]) | (t[0] & t[61] & t[72] & ~t[83]) | (t[0] & t[61] & ~t[72] & t[83]) | (t[0] & ~t[61] & t[72] & t[83]) | (~t[0] & t[61] & t[72] & t[83]);
endmodule

module R2ind171(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[2]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[11]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[19]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[25]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[49]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[1]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[10]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[18]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[48]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[54]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [58:0] x;
 output y;

 wire [137:0] t;
  assign t[0] = t[1] ? t[2] : t[61];
  assign t[100] = t[122] ^ x[27];
  assign t[101] = t[123] ^ x[28];
  assign t[102] = t[124] ^ x[33];
  assign t[103] = t[125] ^ x[34];
  assign t[104] = t[126] ^ x[36];
  assign t[105] = t[127] ^ x[37];
  assign t[106] = t[128] ^ x[39];
  assign t[107] = t[129] ^ x[40];
  assign t[108] = t[130] ^ x[42];
  assign t[109] = t[131] ^ x[43];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[132] ^ x[45];
  assign t[111] = t[133] ^ x[46];
  assign t[112] = t[134] ^ x[51];
  assign t[113] = t[135] ^ x[52];
  assign t[114] = t[136] ^ x[57];
  assign t[115] = t[137] ^ x[58];
  assign t[116] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[117] = (x[0]);
  assign t[118] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[119] = (x[9]);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[121] = (x[17]);
  assign t[122] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[123] = (x[23]);
  assign t[124] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[125] = (x[29]);
  assign t[126] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[127] = (x[35]);
  assign t[128] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[129] = (x[38]);
  assign t[12] = ~(t[63] ^ t[17]);
  assign t[130] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[131] = (x[41]);
  assign t[132] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[133] = (x[44]);
  assign t[134] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[135] = (x[47]);
  assign t[136] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[137] = (x[53]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[64] ^ t[65]);
  assign t[15] = ~(t[66] & t[67]);
  assign t[16] = ~(t[68] & t[69]);
  assign t[17] = ~(t[70] ^ t[71]);
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26]);
  assign t[23] = ~(t[68]);
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[29] & t[30]);
  assign t[26] = ~(t[27] | t[31]);
  assign t[27] = ~(t[32]);
  assign t[28] = t[66] ? t[34] : t[33];
  assign t[29] = ~(t[35] | t[36]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[37] | t[38]);
  assign t[31] = t[66] ? t[40] : t[39];
  assign t[32] = ~(t[68]);
  assign t[33] = ~(t[41] & t[42]);
  assign t[34] = ~(x[7] & t[43]);
  assign t[35] = ~(t[27] | t[44]);
  assign t[36] = ~(t[45] & t[46]);
  assign t[37] = ~(t[32] | t[47]);
  assign t[38] = ~(t[32] | t[48]);
  assign t[39] = ~(t[49] & t[69]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[50] & t[42]);
  assign t[41] = ~(x[7] | t[51]);
  assign t[42] = ~(t[69]);
  assign t[43] = ~(t[67] | t[42]);
  assign t[44] = t[66] ? t[39] : t[40];
  assign t[45] = ~(t[52] | t[53]);
  assign t[46] = ~(t[32] & t[54]);
  assign t[47] = t[66] ? t[55] : t[40];
  assign t[48] = t[66] ? t[33] : t[56];
  assign t[49] = x[7] & t[67];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = ~(x[7] | t[67]);
  assign t[51] = ~(t[67]);
  assign t[52] = ~(t[32] | t[57]);
  assign t[53] = ~(t[27] | t[58]);
  assign t[54] = ~(t[56] & t[59]);
  assign t[55] = ~(t[49] & t[42]);
  assign t[56] = ~(x[7] & t[60]);
  assign t[57] = t[66] ? t[40] : t[55];
  assign t[58] = t[66] ? t[33] : t[34];
  assign t[59] = ~(t[69] & t[41]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[67] | t[69]);
  assign t[61] = (t[72]);
  assign t[62] = (t[73]);
  assign t[63] = (t[74]);
  assign t[64] = (t[75]);
  assign t[65] = (t[76]);
  assign t[66] = (t[77]);
  assign t[67] = (t[78]);
  assign t[68] = (t[79]);
  assign t[69] = (t[80]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (t[81]);
  assign t[71] = (t[82]);
  assign t[72] = t[83] ^ x[5];
  assign t[73] = t[84] ^ x[14];
  assign t[74] = t[85] ^ x[22];
  assign t[75] = t[86] ^ x[28];
  assign t[76] = t[87] ^ x[34];
  assign t[77] = t[88] ^ x[37];
  assign t[78] = t[89] ^ x[40];
  assign t[79] = t[90] ^ x[43];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[91] ^ x[46];
  assign t[81] = t[92] ^ x[52];
  assign t[82] = t[93] ^ x[58];
  assign t[83] = (~t[94] & t[95]);
  assign t[84] = (~t[96] & t[97]);
  assign t[85] = (~t[98] & t[99]);
  assign t[86] = (~t[100] & t[101]);
  assign t[87] = (~t[102] & t[103]);
  assign t[88] = (~t[104] & t[105]);
  assign t[89] = (~t[106] & t[107]);
  assign t[8] = ~(t[62] ^ t[14]);
  assign t[90] = (~t[108] & t[109]);
  assign t[91] = (~t[110] & t[111]);
  assign t[92] = (~t[112] & t[113]);
  assign t[93] = (~t[114] & t[115]);
  assign t[94] = t[116] ^ x[4];
  assign t[95] = t[117] ^ x[5];
  assign t[96] = t[118] ^ x[13];
  assign t[97] = t[119] ^ x[14];
  assign t[98] = t[120] ^ x[21];
  assign t[99] = t[121] ^ x[22];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [88:0] x;
 output y;

 wire [264:0] t;
  assign t[0] = t[1] ? t[2] : t[83];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = t[147] ^ x[5];
  assign t[116] = t[148] ^ x[14];
  assign t[117] = t[149] ^ x[22];
  assign t[118] = t[150] ^ x[28];
  assign t[119] = t[151] ^ x[34];
  assign t[11] = ~(x[6]);
  assign t[120] = t[152] ^ x[37];
  assign t[121] = t[153] ^ x[40];
  assign t[122] = t[154] ^ x[43];
  assign t[123] = t[155] ^ x[46];
  assign t[124] = t[156] ^ x[52];
  assign t[125] = t[157] ^ x[58];
  assign t[126] = t[158] ^ x[59];
  assign t[127] = t[159] ^ x[61];
  assign t[128] = t[160] ^ x[64];
  assign t[129] = t[161] ^ x[65];
  assign t[12] = ~(t[85] ^ t[17]);
  assign t[130] = t[162] ^ x[66];
  assign t[131] = t[163] ^ x[67];
  assign t[132] = t[164] ^ x[68];
  assign t[133] = t[165] ^ x[69];
  assign t[134] = t[166] ^ x[71];
  assign t[135] = t[167] ^ x[74];
  assign t[136] = t[168] ^ x[75];
  assign t[137] = t[169] ^ x[76];
  assign t[138] = t[170] ^ x[77];
  assign t[139] = t[171] ^ x[78];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[79];
  assign t[141] = t[173] ^ x[81];
  assign t[142] = t[174] ^ x[84];
  assign t[143] = t[175] ^ x[85];
  assign t[144] = t[176] ^ x[86];
  assign t[145] = t[177] ^ x[87];
  assign t[146] = t[178] ^ x[88];
  assign t[147] = (~t[179] & t[180]);
  assign t[148] = (~t[181] & t[182]);
  assign t[149] = (~t[183] & t[184]);
  assign t[14] = ~(t[86] ^ t[87]);
  assign t[150] = (~t[185] & t[186]);
  assign t[151] = (~t[187] & t[188]);
  assign t[152] = (~t[189] & t[190]);
  assign t[153] = (~t[191] & t[192]);
  assign t[154] = (~t[193] & t[194]);
  assign t[155] = (~t[195] & t[196]);
  assign t[156] = (~t[197] & t[198]);
  assign t[157] = (~t[199] & t[200]);
  assign t[158] = (~t[179] & t[201]);
  assign t[159] = (~t[181] & t[202]);
  assign t[15] = ~(t[88] & t[89]);
  assign t[160] = (~t[183] & t[203]);
  assign t[161] = (~t[187] & t[204]);
  assign t[162] = (~t[185] & t[205]);
  assign t[163] = (~t[199] & t[206]);
  assign t[164] = (~t[197] & t[207]);
  assign t[165] = (~t[179] & t[208]);
  assign t[166] = (~t[181] & t[209]);
  assign t[167] = (~t[183] & t[210]);
  assign t[168] = (~t[185] & t[211]);
  assign t[169] = (~t[187] & t[212]);
  assign t[16] = ~(t[90] & t[91]);
  assign t[170] = (~t[197] & t[213]);
  assign t[171] = (~t[199] & t[214]);
  assign t[172] = (~t[179] & t[215]);
  assign t[173] = (~t[181] & t[216]);
  assign t[174] = (~t[183] & t[217]);
  assign t[175] = (~t[185] & t[218]);
  assign t[176] = (~t[187] & t[219]);
  assign t[177] = (~t[197] & t[220]);
  assign t[178] = (~t[199] & t[221]);
  assign t[179] = t[222] ^ x[4];
  assign t[17] = ~(t[92] ^ t[93]);
  assign t[180] = t[223] ^ x[5];
  assign t[181] = t[224] ^ x[13];
  assign t[182] = t[225] ^ x[14];
  assign t[183] = t[226] ^ x[21];
  assign t[184] = t[227] ^ x[22];
  assign t[185] = t[228] ^ x[27];
  assign t[186] = t[229] ^ x[28];
  assign t[187] = t[230] ^ x[33];
  assign t[188] = t[231] ^ x[34];
  assign t[189] = t[232] ^ x[36];
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[190] = t[233] ^ x[37];
  assign t[191] = t[234] ^ x[39];
  assign t[192] = t[235] ^ x[40];
  assign t[193] = t[236] ^ x[42];
  assign t[194] = t[237] ^ x[43];
  assign t[195] = t[238] ^ x[45];
  assign t[196] = t[239] ^ x[46];
  assign t[197] = t[240] ^ x[51];
  assign t[198] = t[241] ^ x[52];
  assign t[199] = t[242] ^ x[57];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[58];
  assign t[201] = t[244] ^ x[59];
  assign t[202] = t[245] ^ x[61];
  assign t[203] = t[246] ^ x[64];
  assign t[204] = t[247] ^ x[65];
  assign t[205] = t[248] ^ x[66];
  assign t[206] = t[249] ^ x[67];
  assign t[207] = t[250] ^ x[68];
  assign t[208] = t[251] ^ x[69];
  assign t[209] = t[252] ^ x[71];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[74];
  assign t[211] = t[254] ^ x[75];
  assign t[212] = t[255] ^ x[76];
  assign t[213] = t[256] ^ x[77];
  assign t[214] = t[257] ^ x[78];
  assign t[215] = t[258] ^ x[79];
  assign t[216] = t[259] ^ x[81];
  assign t[217] = t[260] ^ x[84];
  assign t[218] = t[261] ^ x[85];
  assign t[219] = t[262] ^ x[86];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[87];
  assign t[221] = t[264] ^ x[88];
  assign t[222] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[223] = (x[0]);
  assign t[224] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[225] = (x[9]);
  assign t[226] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[227] = (x[17]);
  assign t[228] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[229] = (x[23]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[230] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[231] = (x[29]);
  assign t[232] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[233] = (x[35]);
  assign t[234] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[235] = (x[38]);
  assign t[236] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[237] = (x[41]);
  assign t[238] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[239] = (x[44]);
  assign t[23] = ~(t[90]);
  assign t[240] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[241] = (x[47]);
  assign t[242] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[243] = (x[53]);
  assign t[244] = (x[1]);
  assign t[245] = (x[10]);
  assign t[246] = (x[18]);
  assign t[247] = (x[30]);
  assign t[248] = (x[24]);
  assign t[249] = (x[54]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[250] = (x[48]);
  assign t[251] = (x[2]);
  assign t[252] = (x[11]);
  assign t[253] = (x[19]);
  assign t[254] = (x[25]);
  assign t[255] = (x[31]);
  assign t[256] = (x[49]);
  assign t[257] = (x[55]);
  assign t[258] = (x[3]);
  assign t[259] = (x[12]);
  assign t[25] = ~(t[28] | t[30]);
  assign t[260] = (x[20]);
  assign t[261] = (x[26]);
  assign t[262] = (x[32]);
  assign t[263] = (x[50]);
  assign t[264] = (x[56]);
  assign t[26] = t[91] & t[31];
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[33]);
  assign t[29] = t[88] ? t[35] : t[34];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[88] ? t[37] : t[36];
  assign t[31] = ~(t[33] | t[88]);
  assign t[32] = ~(t[38] | t[39]);
  assign t[33] = ~(t[90]);
  assign t[34] = ~(t[91] & t[40]);
  assign t[35] = ~(x[7] & t[41]);
  assign t[36] = ~(t[42] & t[91]);
  assign t[37] = ~(t[43] & t[44]);
  assign t[38] = ~(t[33] | t[45]);
  assign t[39] = ~(t[33] | t[46]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(x[7] | t[47]);
  assign t[41] = ~(t[89] | t[91]);
  assign t[42] = ~(x[7] | t[89]);
  assign t[43] = x[7] & t[89];
  assign t[44] = ~(t[91]);
  assign t[45] = t[88] ? t[37] : t[48];
  assign t[46] = t[88] ? t[49] : t[35];
  assign t[47] = ~(t[89]);
  assign t[48] = ~(t[42] & t[44]);
  assign t[49] = ~(t[40] & t[44]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[1] ? t[51] : t[94];
  assign t[51] = x[6] ? t[53] : t[52];
  assign t[52] = x[7] ? t[55] : t[54];
  assign t[53] = t[56] ^ x[60];
  assign t[54] = t[57] ^ t[58];
  assign t[55] = ~(t[95] ^ t[59]);
  assign t[56] = x[62] ^ x[63];
  assign t[57] = t[20] ? x[63] : x[62];
  assign t[58] = ~(t[96] ^ t[60]);
  assign t[59] = ~(t[97] ^ t[98]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = ~(t[99] ^ t[100]);
  assign t[61] = t[1] ? t[62] : t[101];
  assign t[62] = x[6] ? t[64] : t[63];
  assign t[63] = x[7] ? t[66] : t[65];
  assign t[64] = t[67] ^ x[70];
  assign t[65] = t[68] ^ t[69];
  assign t[66] = ~(t[102] ^ t[70]);
  assign t[67] = x[72] ^ x[73];
  assign t[68] = t[20] ? x[73] : x[72];
  assign t[69] = ~(t[103] ^ t[71]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = ~(t[104] ^ t[105]);
  assign t[71] = ~(t[106] ^ t[107]);
  assign t[72] = t[1] ? t[73] : t[108];
  assign t[73] = x[6] ? t[75] : t[74];
  assign t[74] = x[7] ? t[77] : t[76];
  assign t[75] = t[78] ^ x[80];
  assign t[76] = t[79] ^ t[80];
  assign t[77] = ~(t[109] ^ t[81]);
  assign t[78] = x[82] ^ x[83];
  assign t[79] = t[20] ? x[83] : x[82];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = ~(t[110] ^ t[82]);
  assign t[81] = ~(t[111] ^ t[112]);
  assign t[82] = ~(t[113] ^ t[114]);
  assign t[83] = (t[115]);
  assign t[84] = (t[116]);
  assign t[85] = (t[117]);
  assign t[86] = (t[118]);
  assign t[87] = (t[119]);
  assign t[88] = (t[120]);
  assign t[89] = (t[121]);
  assign t[8] = ~(t[84] ^ t[14]);
  assign t[90] = (t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[50] & ~t[61] & ~t[72]) | (~t[0] & t[50] & ~t[61] & ~t[72]) | (~t[0] & ~t[50] & t[61] & ~t[72]) | (~t[0] & ~t[50] & ~t[61] & t[72]) | (t[0] & t[50] & t[61] & ~t[72]) | (t[0] & t[50] & ~t[61] & t[72]) | (t[0] & ~t[50] & t[61] & t[72]) | (~t[0] & t[50] & t[61] & t[72]);
endmodule

module R2ind176(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[2]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[11]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[19]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[25]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[49]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[1]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[10]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[18]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[48]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[54]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [58:0] x;
 output y;

 wire [126:0] t;
  assign t[0] = t[1] ? t[2] : t[50];
  assign t[100] = t[122] ^ x[46];
  assign t[101] = t[123] ^ x[51];
  assign t[102] = t[124] ^ x[52];
  assign t[103] = t[125] ^ x[57];
  assign t[104] = t[126] ^ x[58];
  assign t[105] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[106] = (x[0]);
  assign t[107] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[108] = (x[9]);
  assign t[109] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (x[17]);
  assign t[111] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[112] = (x[23]);
  assign t[113] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[114] = (x[29]);
  assign t[115] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[116] = (x[35]);
  assign t[117] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[118] = (x[38]);
  assign t[119] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[41]);
  assign t[121] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[122] = (x[44]);
  assign t[123] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[124] = (x[47]);
  assign t[125] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[126] = (x[53]);
  assign t[12] = ~(t[52] ^ t[17]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[53] ^ t[54]);
  assign t[15] = ~(t[55] & t[56]);
  assign t[16] = ~(t[57] & t[58]);
  assign t[17] = ~(t[59] ^ t[60]);
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[57]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[25] = ~(t[28] | t[30]);
  assign t[26] = t[58] & t[31];
  assign t[27] = ~(t[32]);
  assign t[28] = ~(t[33]);
  assign t[29] = t[55] ? t[35] : t[34];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[55] ? t[37] : t[36];
  assign t[31] = ~(t[33] | t[55]);
  assign t[32] = ~(t[38] | t[39]);
  assign t[33] = ~(t[57]);
  assign t[34] = ~(t[58] & t[40]);
  assign t[35] = ~(x[7] & t[41]);
  assign t[36] = ~(t[42] & t[58]);
  assign t[37] = ~(t[43] & t[44]);
  assign t[38] = ~(t[33] | t[45]);
  assign t[39] = ~(t[33] | t[46]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(x[7] | t[47]);
  assign t[41] = ~(t[56] | t[58]);
  assign t[42] = ~(x[7] | t[56]);
  assign t[43] = x[7] & t[56];
  assign t[44] = ~(t[58]);
  assign t[45] = t[55] ? t[37] : t[48];
  assign t[46] = t[55] ? t[49] : t[35];
  assign t[47] = ~(t[56]);
  assign t[48] = ~(t[42] & t[44]);
  assign t[49] = ~(t[40] & t[44]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (t[61]);
  assign t[51] = (t[62]);
  assign t[52] = (t[63]);
  assign t[53] = (t[64]);
  assign t[54] = (t[65]);
  assign t[55] = (t[66]);
  assign t[56] = (t[67]);
  assign t[57] = (t[68]);
  assign t[58] = (t[69]);
  assign t[59] = (t[70]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = t[72] ^ x[5];
  assign t[62] = t[73] ^ x[14];
  assign t[63] = t[74] ^ x[22];
  assign t[64] = t[75] ^ x[28];
  assign t[65] = t[76] ^ x[34];
  assign t[66] = t[77] ^ x[37];
  assign t[67] = t[78] ^ x[40];
  assign t[68] = t[79] ^ x[43];
  assign t[69] = t[80] ^ x[46];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[81] ^ x[52];
  assign t[71] = t[82] ^ x[58];
  assign t[72] = (~t[83] & t[84]);
  assign t[73] = (~t[85] & t[86]);
  assign t[74] = (~t[87] & t[88]);
  assign t[75] = (~t[89] & t[90]);
  assign t[76] = (~t[91] & t[92]);
  assign t[77] = (~t[93] & t[94]);
  assign t[78] = (~t[95] & t[96]);
  assign t[79] = (~t[97] & t[98]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[99] & t[100]);
  assign t[81] = (~t[101] & t[102]);
  assign t[82] = (~t[103] & t[104]);
  assign t[83] = t[105] ^ x[4];
  assign t[84] = t[106] ^ x[5];
  assign t[85] = t[107] ^ x[13];
  assign t[86] = t[108] ^ x[14];
  assign t[87] = t[109] ^ x[21];
  assign t[88] = t[110] ^ x[22];
  assign t[89] = t[111] ^ x[27];
  assign t[8] = ~(t[51] ^ t[14]);
  assign t[90] = t[112] ^ x[28];
  assign t[91] = t[113] ^ x[33];
  assign t[92] = t[114] ^ x[34];
  assign t[93] = t[115] ^ x[36];
  assign t[94] = t[116] ^ x[37];
  assign t[95] = t[117] ^ x[39];
  assign t[96] = t[118] ^ x[40];
  assign t[97] = t[119] ^ x[42];
  assign t[98] = t[120] ^ x[43];
  assign t[99] = t[121] ^ x[45];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [88:0] x;
 output y;

 wire [272:0] t;
  assign t[0] = t[1] ? t[2] : t[91];
  assign t[100] = (t[132]);
  assign t[101] = (t[133]);
  assign t[102] = (t[134]);
  assign t[103] = (t[135]);
  assign t[104] = (t[136]);
  assign t[105] = (t[137]);
  assign t[106] = (t[138]);
  assign t[107] = (t[139]);
  assign t[108] = (t[140]);
  assign t[109] = (t[141]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = (t[142]);
  assign t[111] = (t[143]);
  assign t[112] = (t[144]);
  assign t[113] = (t[145]);
  assign t[114] = (t[146]);
  assign t[115] = (t[147]);
  assign t[116] = (t[148]);
  assign t[117] = (t[149]);
  assign t[118] = (t[150]);
  assign t[119] = (t[151]);
  assign t[11] = ~(x[6]);
  assign t[120] = (t[152]);
  assign t[121] = (t[153]);
  assign t[122] = (t[154]);
  assign t[123] = t[155] ^ x[5];
  assign t[124] = t[156] ^ x[14];
  assign t[125] = t[157] ^ x[22];
  assign t[126] = t[158] ^ x[28];
  assign t[127] = t[159] ^ x[34];
  assign t[128] = t[160] ^ x[37];
  assign t[129] = t[161] ^ x[40];
  assign t[12] = ~(t[93] ^ t[17]);
  assign t[130] = t[162] ^ x[43];
  assign t[131] = t[163] ^ x[46];
  assign t[132] = t[164] ^ x[52];
  assign t[133] = t[165] ^ x[58];
  assign t[134] = t[166] ^ x[59];
  assign t[135] = t[167] ^ x[61];
  assign t[136] = t[168] ^ x[64];
  assign t[137] = t[169] ^ x[65];
  assign t[138] = t[170] ^ x[66];
  assign t[139] = t[171] ^ x[67];
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[140] = t[172] ^ x[68];
  assign t[141] = t[173] ^ x[69];
  assign t[142] = t[174] ^ x[71];
  assign t[143] = t[175] ^ x[74];
  assign t[144] = t[176] ^ x[75];
  assign t[145] = t[177] ^ x[76];
  assign t[146] = t[178] ^ x[77];
  assign t[147] = t[179] ^ x[78];
  assign t[148] = t[180] ^ x[79];
  assign t[149] = t[181] ^ x[81];
  assign t[14] = ~(t[94] ^ t[95]);
  assign t[150] = t[182] ^ x[84];
  assign t[151] = t[183] ^ x[85];
  assign t[152] = t[184] ^ x[86];
  assign t[153] = t[185] ^ x[87];
  assign t[154] = t[186] ^ x[88];
  assign t[155] = (~t[187] & t[188]);
  assign t[156] = (~t[189] & t[190]);
  assign t[157] = (~t[191] & t[192]);
  assign t[158] = (~t[193] & t[194]);
  assign t[159] = (~t[195] & t[196]);
  assign t[15] = ~(t[96] & t[97]);
  assign t[160] = (~t[197] & t[198]);
  assign t[161] = (~t[199] & t[200]);
  assign t[162] = (~t[201] & t[202]);
  assign t[163] = (~t[203] & t[204]);
  assign t[164] = (~t[205] & t[206]);
  assign t[165] = (~t[207] & t[208]);
  assign t[166] = (~t[187] & t[209]);
  assign t[167] = (~t[189] & t[210]);
  assign t[168] = (~t[191] & t[211]);
  assign t[169] = (~t[195] & t[212]);
  assign t[16] = ~(t[98] & t[99]);
  assign t[170] = (~t[193] & t[213]);
  assign t[171] = (~t[207] & t[214]);
  assign t[172] = (~t[205] & t[215]);
  assign t[173] = (~t[187] & t[216]);
  assign t[174] = (~t[189] & t[217]);
  assign t[175] = (~t[191] & t[218]);
  assign t[176] = (~t[193] & t[219]);
  assign t[177] = (~t[195] & t[220]);
  assign t[178] = (~t[207] & t[221]);
  assign t[179] = (~t[205] & t[222]);
  assign t[17] = ~(t[100] ^ t[101]);
  assign t[180] = (~t[187] & t[223]);
  assign t[181] = (~t[189] & t[224]);
  assign t[182] = (~t[191] & t[225]);
  assign t[183] = (~t[193] & t[226]);
  assign t[184] = (~t[195] & t[227]);
  assign t[185] = (~t[207] & t[228]);
  assign t[186] = (~t[205] & t[229]);
  assign t[187] = t[230] ^ x[4];
  assign t[188] = t[231] ^ x[5];
  assign t[189] = t[232] ^ x[13];
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[190] = t[233] ^ x[14];
  assign t[191] = t[234] ^ x[21];
  assign t[192] = t[235] ^ x[22];
  assign t[193] = t[236] ^ x[27];
  assign t[194] = t[237] ^ x[28];
  assign t[195] = t[238] ^ x[33];
  assign t[196] = t[239] ^ x[34];
  assign t[197] = t[240] ^ x[36];
  assign t[198] = t[241] ^ x[37];
  assign t[199] = t[242] ^ x[39];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[200] = t[243] ^ x[40];
  assign t[201] = t[244] ^ x[42];
  assign t[202] = t[245] ^ x[43];
  assign t[203] = t[246] ^ x[45];
  assign t[204] = t[247] ^ x[46];
  assign t[205] = t[248] ^ x[51];
  assign t[206] = t[249] ^ x[52];
  assign t[207] = t[250] ^ x[57];
  assign t[208] = t[251] ^ x[58];
  assign t[209] = t[252] ^ x[59];
  assign t[20] = ~(t[23]);
  assign t[210] = t[253] ^ x[61];
  assign t[211] = t[254] ^ x[64];
  assign t[212] = t[255] ^ x[65];
  assign t[213] = t[256] ^ x[66];
  assign t[214] = t[257] ^ x[67];
  assign t[215] = t[258] ^ x[68];
  assign t[216] = t[259] ^ x[69];
  assign t[217] = t[260] ^ x[71];
  assign t[218] = t[261] ^ x[74];
  assign t[219] = t[262] ^ x[75];
  assign t[21] = ~(t[24] | t[25]);
  assign t[220] = t[263] ^ x[76];
  assign t[221] = t[264] ^ x[77];
  assign t[222] = t[265] ^ x[78];
  assign t[223] = t[266] ^ x[79];
  assign t[224] = t[267] ^ x[81];
  assign t[225] = t[268] ^ x[84];
  assign t[226] = t[269] ^ x[85];
  assign t[227] = t[270] ^ x[86];
  assign t[228] = t[271] ^ x[87];
  assign t[229] = t[272] ^ x[88];
  assign t[22] = ~(t[26] | t[27]);
  assign t[230] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[231] = (x[0]);
  assign t[232] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[233] = (x[9]);
  assign t[234] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[235] = (x[17]);
  assign t[236] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[237] = (x[23]);
  assign t[238] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[239] = (x[29]);
  assign t[23] = ~(t[98]);
  assign t[240] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[241] = (x[35]);
  assign t[242] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[243] = (x[38]);
  assign t[244] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[245] = (x[41]);
  assign t[246] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[247] = (x[44]);
  assign t[248] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[249] = (x[47]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[250] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[251] = (x[53]);
  assign t[252] = (x[1]);
  assign t[253] = (x[10]);
  assign t[254] = (x[18]);
  assign t[255] = (x[30]);
  assign t[256] = (x[24]);
  assign t[257] = (x[54]);
  assign t[258] = (x[48]);
  assign t[259] = (x[2]);
  assign t[25] = ~(t[28] | t[30]);
  assign t[260] = (x[11]);
  assign t[261] = (x[19]);
  assign t[262] = (x[25]);
  assign t[263] = (x[31]);
  assign t[264] = (x[55]);
  assign t[265] = (x[49]);
  assign t[266] = (x[3]);
  assign t[267] = (x[12]);
  assign t[268] = (x[20]);
  assign t[269] = (x[26]);
  assign t[26] = ~(t[31] & t[32]);
  assign t[270] = (x[32]);
  assign t[271] = (x[56]);
  assign t[272] = (x[50]);
  assign t[27] = ~(t[33] & t[34]);
  assign t[28] = ~(t[98]);
  assign t[29] = t[96] ? t[36] : t[35];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[96] ? t[38] : t[37];
  assign t[31] = ~(t[39] | t[40]);
  assign t[32] = ~(t[28] & t[41]);
  assign t[33] = ~(t[42] & t[43]);
  assign t[34] = t[28] | t[44];
  assign t[35] = ~(t[45] & t[46]);
  assign t[36] = ~(t[47] & t[46]);
  assign t[37] = ~(x[7] & t[48]);
  assign t[38] = ~(t[49] & t[46]);
  assign t[39] = ~(t[28] | t[50]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[51] | t[52]);
  assign t[41] = ~(t[37] & t[53]);
  assign t[42] = t[99] & t[54];
  assign t[43] = t[45] | t[47];
  assign t[44] = t[96] ? t[37] : t[38];
  assign t[45] = ~(x[7] | t[97]);
  assign t[46] = ~(t[99]);
  assign t[47] = x[7] & t[97];
  assign t[48] = ~(t[97] | t[99]);
  assign t[49] = ~(x[7] | t[55]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[96] ? t[35] : t[36];
  assign t[51] = ~(t[28]);
  assign t[52] = t[96] ? t[38] : t[56];
  assign t[53] = ~(t[99] & t[49]);
  assign t[54] = ~(t[28] | t[96]);
  assign t[55] = ~(t[97]);
  assign t[56] = ~(x[7] & t[57]);
  assign t[57] = ~(t[97] | t[46]);
  assign t[58] = t[1] ? t[59] : t[102];
  assign t[59] = x[6] ? t[61] : t[60];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = x[7] ? t[63] : t[62];
  assign t[61] = t[64] ^ x[60];
  assign t[62] = t[65] ^ t[66];
  assign t[63] = ~(t[103] ^ t[67]);
  assign t[64] = x[62] ^ x[63];
  assign t[65] = t[20] ? x[63] : x[62];
  assign t[66] = ~(t[104] ^ t[68]);
  assign t[67] = ~(t[105] ^ t[106]);
  assign t[68] = ~(t[107] ^ t[108]);
  assign t[69] = t[1] ? t[70] : t[109];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = x[6] ? t[72] : t[71];
  assign t[71] = x[7] ? t[74] : t[73];
  assign t[72] = t[75] ^ x[70];
  assign t[73] = t[76] ^ t[77];
  assign t[74] = ~(t[110] ^ t[78]);
  assign t[75] = x[72] ^ x[73];
  assign t[76] = t[20] ? x[73] : x[72];
  assign t[77] = ~(t[111] ^ t[79]);
  assign t[78] = ~(t[112] ^ t[113]);
  assign t[79] = ~(t[114] ^ t[115]);
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = t[1] ? t[81] : t[116];
  assign t[81] = x[6] ? t[83] : t[82];
  assign t[82] = x[7] ? t[85] : t[84];
  assign t[83] = t[86] ^ x[80];
  assign t[84] = t[87] ^ t[88];
  assign t[85] = ~(t[117] ^ t[89]);
  assign t[86] = x[82] ^ x[83];
  assign t[87] = t[20] ? x[83] : x[82];
  assign t[88] = ~(t[118] ^ t[90]);
  assign t[89] = ~(t[119] ^ t[120]);
  assign t[8] = ~(t[92] ^ t[14]);
  assign t[90] = ~(t[121] ^ t[122]);
  assign t[91] = (t[123]);
  assign t[92] = (t[124]);
  assign t[93] = (t[125]);
  assign t[94] = (t[126]);
  assign t[95] = (t[127]);
  assign t[96] = (t[128]);
  assign t[97] = (t[129]);
  assign t[98] = (t[130]);
  assign t[99] = (t[131]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[58] & ~t[69] & ~t[80]) | (~t[0] & t[58] & ~t[69] & ~t[80]) | (~t[0] & ~t[58] & t[69] & ~t[80]) | (~t[0] & ~t[58] & ~t[69] & t[80]) | (t[0] & t[58] & t[69] & ~t[80]) | (t[0] & t[58] & ~t[69] & t[80]) | (t[0] & ~t[58] & t[69] & t[80]) | (~t[0] & t[58] & t[69] & t[80]);
endmodule

module R2ind181(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[3]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[12]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[20]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[26]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[32]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[50]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[56]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[2]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[11]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[19]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[25]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[31]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[49]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[55]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [58:0] x;
 output y;

 wire [96:0] t;
  assign t[0] = t[1] ? t[2] : t[20];
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[17] ? x[16] : x[15];
  assign t[13] = ~(t[22] ^ t[18]);
  assign t[14] = ~(t[23] ^ t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = ~(t[19]);
  assign t[18] = ~(t[29] ^ t[30]);
  assign t[19] = ~(t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = (t[41]);
  assign t[31] = t[42] ^ x[5];
  assign t[32] = t[43] ^ x[14];
  assign t[33] = t[44] ^ x[22];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[34];
  assign t[36] = t[47] ^ x[37];
  assign t[37] = t[48] ^ x[40];
  assign t[38] = t[49] ^ x[43];
  assign t[39] = t[50] ^ x[46];
  assign t[3] = ~(t[6]);
  assign t[40] = t[51] ^ x[52];
  assign t[41] = t[52] ^ x[58];
  assign t[42] = (~t[53] & t[54]);
  assign t[43] = (~t[55] & t[56]);
  assign t[44] = (~t[57] & t[58]);
  assign t[45] = (~t[59] & t[60]);
  assign t[46] = (~t[61] & t[62]);
  assign t[47] = (~t[63] & t[64]);
  assign t[48] = (~t[65] & t[66]);
  assign t[49] = (~t[67] & t[68]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (~t[69] & t[70]);
  assign t[51] = (~t[71] & t[72]);
  assign t[52] = (~t[73] & t[74]);
  assign t[53] = t[75] ^ x[4];
  assign t[54] = t[76] ^ x[5];
  assign t[55] = t[77] ^ x[13];
  assign t[56] = t[78] ^ x[14];
  assign t[57] = t[79] ^ x[21];
  assign t[58] = t[80] ^ x[22];
  assign t[59] = t[81] ^ x[27];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[82] ^ x[28];
  assign t[61] = t[83] ^ x[33];
  assign t[62] = t[84] ^ x[34];
  assign t[63] = t[85] ^ x[36];
  assign t[64] = t[86] ^ x[37];
  assign t[65] = t[87] ^ x[39];
  assign t[66] = t[88] ^ x[40];
  assign t[67] = t[89] ^ x[42];
  assign t[68] = t[90] ^ x[43];
  assign t[69] = t[91] ^ x[45];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[92] ^ x[46];
  assign t[71] = t[93] ^ x[51];
  assign t[72] = t[94] ^ x[52];
  assign t[73] = t[95] ^ x[57];
  assign t[74] = t[96] ^ x[58];
  assign t[75] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[76] = (x[1]);
  assign t[77] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[78] = (x[10]);
  assign t[79] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[7] = t[12] ^ t[13];
  assign t[80] = (x[18]);
  assign t[81] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[82] = (x[24]);
  assign t[83] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[84] = (x[30]);
  assign t[85] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[35]);
  assign t[87] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[38]);
  assign t[89] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[21] ^ t[14]);
  assign t[90] = (x[41]);
  assign t[91] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[44]);
  assign t[93] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[94] = (x[48]);
  assign t[95] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[96] = (x[54]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [58:0] x;
 output y;

 wire [134:0] t;
  assign t[0] = t[1] ? t[2] : t[58];
  assign t[100] = t[122] ^ x[34];
  assign t[101] = t[123] ^ x[36];
  assign t[102] = t[124] ^ x[37];
  assign t[103] = t[125] ^ x[39];
  assign t[104] = t[126] ^ x[40];
  assign t[105] = t[127] ^ x[42];
  assign t[106] = t[128] ^ x[43];
  assign t[107] = t[129] ^ x[45];
  assign t[108] = t[130] ^ x[46];
  assign t[109] = t[131] ^ x[51];
  assign t[10] = ~(t[15] | t[16]);
  assign t[110] = t[132] ^ x[52];
  assign t[111] = t[133] ^ x[57];
  assign t[112] = t[134] ^ x[58];
  assign t[113] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[114] = (x[0]);
  assign t[115] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[116] = (x[9]);
  assign t[117] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[118] = (x[17]);
  assign t[119] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[11] = ~(x[6]);
  assign t[120] = (x[23]);
  assign t[121] = (x[29] & ~x[30] & ~x[31] & ~x[32]) | (~x[29] & x[30] & ~x[31] & ~x[32]) | (~x[29] & ~x[30] & x[31] & ~x[32]) | (~x[29] & ~x[30] & ~x[31] & x[32]) | (x[29] & x[30] & x[31] & ~x[32]) | (x[29] & x[30] & ~x[31] & x[32]) | (x[29] & ~x[30] & x[31] & x[32]) | (~x[29] & x[30] & x[31] & x[32]);
  assign t[122] = (x[29]);
  assign t[123] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[124] = (x[35]);
  assign t[125] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[126] = (x[38]);
  assign t[127] = (x[41] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[41] & 1'b0 & ~1'b0 & ~1'b0) | (~x[41] & ~1'b0 & 1'b0 & ~1'b0) | (~x[41] & ~1'b0 & ~1'b0 & 1'b0) | (x[41] & 1'b0 & 1'b0 & ~1'b0) | (x[41] & 1'b0 & ~1'b0 & 1'b0) | (x[41] & ~1'b0 & 1'b0 & 1'b0) | (~x[41] & 1'b0 & 1'b0 & 1'b0);
  assign t[128] = (x[41]);
  assign t[129] = (x[44] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[44] & 1'b0 & ~1'b0 & ~1'b0) | (~x[44] & ~1'b0 & 1'b0 & ~1'b0) | (~x[44] & ~1'b0 & ~1'b0 & 1'b0) | (x[44] & 1'b0 & 1'b0 & ~1'b0) | (x[44] & 1'b0 & ~1'b0 & 1'b0) | (x[44] & ~1'b0 & 1'b0 & 1'b0) | (~x[44] & 1'b0 & 1'b0 & 1'b0);
  assign t[12] = ~(t[60] ^ t[17]);
  assign t[130] = (x[44]);
  assign t[131] = (x[47] & ~x[48] & ~x[49] & ~x[50]) | (~x[47] & x[48] & ~x[49] & ~x[50]) | (~x[47] & ~x[48] & x[49] & ~x[50]) | (~x[47] & ~x[48] & ~x[49] & x[50]) | (x[47] & x[48] & x[49] & ~x[50]) | (x[47] & x[48] & ~x[49] & x[50]) | (x[47] & ~x[48] & x[49] & x[50]) | (~x[47] & x[48] & x[49] & x[50]);
  assign t[132] = (x[47]);
  assign t[133] = (x[53] & ~x[54] & ~x[55] & ~x[56]) | (~x[53] & x[54] & ~x[55] & ~x[56]) | (~x[53] & ~x[54] & x[55] & ~x[56]) | (~x[53] & ~x[54] & ~x[55] & x[56]) | (x[53] & x[54] & x[55] & ~x[56]) | (x[53] & x[54] & ~x[55] & x[56]) | (x[53] & ~x[54] & x[55] & x[56]) | (~x[53] & x[54] & x[55] & x[56]);
  assign t[134] = (x[53]);
  assign t[13] = ~(t[18] ^ t[19]);
  assign t[14] = ~(t[61] ^ t[62]);
  assign t[15] = ~(t[63] & t[64]);
  assign t[16] = ~(t[65] & t[66]);
  assign t[17] = ~(t[67] ^ t[68]);
  assign t[18] = t[20] ? x[16] : x[15];
  assign t[19] = ~(t[21] & t[22]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[23]);
  assign t[21] = ~(t[24] | t[25]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[65]);
  assign t[24] = ~(t[28] | t[29]);
  assign t[25] = ~(t[28] | t[30]);
  assign t[26] = ~(t[31] & t[32]);
  assign t[27] = ~(t[33] & t[34]);
  assign t[28] = ~(t[65]);
  assign t[29] = t[63] ? t[36] : t[35];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[63] ? t[38] : t[37];
  assign t[31] = ~(t[39] | t[40]);
  assign t[32] = ~(t[28] & t[41]);
  assign t[33] = ~(t[42] & t[43]);
  assign t[34] = t[28] | t[44];
  assign t[35] = ~(t[45] & t[46]);
  assign t[36] = ~(t[47] & t[46]);
  assign t[37] = ~(x[7] & t[48]);
  assign t[38] = ~(t[49] & t[46]);
  assign t[39] = ~(t[28] | t[50]);
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[51] | t[52]);
  assign t[41] = ~(t[37] & t[53]);
  assign t[42] = t[66] & t[54];
  assign t[43] = t[45] | t[47];
  assign t[44] = t[63] ? t[37] : t[38];
  assign t[45] = ~(x[7] | t[64]);
  assign t[46] = ~(t[66]);
  assign t[47] = x[7] & t[64];
  assign t[48] = ~(t[64] | t[66]);
  assign t[49] = ~(x[7] | t[55]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[63] ? t[35] : t[36];
  assign t[51] = ~(t[28]);
  assign t[52] = t[63] ? t[38] : t[56];
  assign t[53] = ~(t[66] & t[49]);
  assign t[54] = ~(t[28] | t[63]);
  assign t[55] = ~(t[64]);
  assign t[56] = ~(x[7] & t[57]);
  assign t[57] = ~(t[64] | t[46]);
  assign t[58] = (t[69]);
  assign t[59] = (t[70]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (t[71]);
  assign t[61] = (t[72]);
  assign t[62] = (t[73]);
  assign t[63] = (t[74]);
  assign t[64] = (t[75]);
  assign t[65] = (t[76]);
  assign t[66] = (t[77]);
  assign t[67] = (t[78]);
  assign t[68] = (t[79]);
  assign t[69] = t[80] ^ x[5];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[81] ^ x[14];
  assign t[71] = t[82] ^ x[22];
  assign t[72] = t[83] ^ x[28];
  assign t[73] = t[84] ^ x[34];
  assign t[74] = t[85] ^ x[37];
  assign t[75] = t[86] ^ x[40];
  assign t[76] = t[87] ^ x[43];
  assign t[77] = t[88] ^ x[46];
  assign t[78] = t[89] ^ x[52];
  assign t[79] = t[90] ^ x[58];
  assign t[7] = ~(t[12] ^ t[13]);
  assign t[80] = (~t[91] & t[92]);
  assign t[81] = (~t[93] & t[94]);
  assign t[82] = (~t[95] & t[96]);
  assign t[83] = (~t[97] & t[98]);
  assign t[84] = (~t[99] & t[100]);
  assign t[85] = (~t[101] & t[102]);
  assign t[86] = (~t[103] & t[104]);
  assign t[87] = (~t[105] & t[106]);
  assign t[88] = (~t[107] & t[108]);
  assign t[89] = (~t[109] & t[110]);
  assign t[8] = ~(t[59] ^ t[14]);
  assign t[90] = (~t[111] & t[112]);
  assign t[91] = t[113] ^ x[4];
  assign t[92] = t[114] ^ x[5];
  assign t[93] = t[115] ^ x[13];
  assign t[94] = t[116] ^ x[14];
  assign t[95] = t[117] ^ x[21];
  assign t[96] = t[118] ^ x[22];
  assign t[97] = t[119] ^ x[27];
  assign t[98] = t[120] ^ x[28];
  assign t[99] = t[121] ^ x[33];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [61:0] x;
 output y;

 wire [192:0] t;
  assign t[0] = t[1] ? t[2] : t[77];
  assign t[100] = t[120] ^ x[28];
  assign t[101] = t[121] ^ x[31];
  assign t[102] = t[122] ^ x[34];
  assign t[103] = t[123] ^ x[37];
  assign t[104] = t[124] ^ x[40];
  assign t[105] = t[125] ^ x[41];
  assign t[106] = t[126] ^ x[43];
  assign t[107] = t[127] ^ x[46];
  assign t[108] = t[128] ^ x[47];
  assign t[109] = t[129] ^ x[48];
  assign t[10] = ~(t[14] | t[15]);
  assign t[110] = t[130] ^ x[50];
  assign t[111] = t[131] ^ x[53];
  assign t[112] = t[132] ^ x[54];
  assign t[113] = t[133] ^ x[55];
  assign t[114] = t[134] ^ x[57];
  assign t[115] = t[135] ^ x[60];
  assign t[116] = t[136] ^ x[61];
  assign t[117] = (~t[137] & t[138]);
  assign t[118] = (~t[139] & t[140]);
  assign t[119] = (~t[141] & t[142]);
  assign t[11] = ~(x[6]);
  assign t[120] = (~t[143] & t[144]);
  assign t[121] = (~t[145] & t[146]);
  assign t[122] = (~t[147] & t[148]);
  assign t[123] = (~t[149] & t[150]);
  assign t[124] = (~t[151] & t[152]);
  assign t[125] = (~t[137] & t[153]);
  assign t[126] = (~t[139] & t[154]);
  assign t[127] = (~t[143] & t[155]);
  assign t[128] = (~t[141] & t[156]);
  assign t[129] = (~t[137] & t[157]);
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[130] = (~t[139] & t[158]);
  assign t[131] = (~t[143] & t[159]);
  assign t[132] = (~t[141] & t[160]);
  assign t[133] = (~t[137] & t[161]);
  assign t[134] = (~t[139] & t[162]);
  assign t[135] = (~t[143] & t[163]);
  assign t[136] = (~t[141] & t[164]);
  assign t[137] = t[165] ^ x[4];
  assign t[138] = t[166] ^ x[5];
  assign t[139] = t[167] ^ x[13];
  assign t[13] = ~(t[79] ^ t[80]);
  assign t[140] = t[168] ^ x[14];
  assign t[141] = t[169] ^ x[21];
  assign t[142] = t[170] ^ x[22];
  assign t[143] = t[171] ^ x[27];
  assign t[144] = t[172] ^ x[28];
  assign t[145] = t[173] ^ x[30];
  assign t[146] = t[174] ^ x[31];
  assign t[147] = t[175] ^ x[33];
  assign t[148] = t[176] ^ x[34];
  assign t[149] = t[177] ^ x[36];
  assign t[14] = ~(t[81] & t[82]);
  assign t[150] = t[178] ^ x[37];
  assign t[151] = t[179] ^ x[39];
  assign t[152] = t[180] ^ x[40];
  assign t[153] = t[181] ^ x[41];
  assign t[154] = t[182] ^ x[43];
  assign t[155] = t[183] ^ x[46];
  assign t[156] = t[184] ^ x[47];
  assign t[157] = t[185] ^ x[48];
  assign t[158] = t[186] ^ x[50];
  assign t[159] = t[187] ^ x[53];
  assign t[15] = ~(t[83] & t[84]);
  assign t[160] = t[188] ^ x[54];
  assign t[161] = t[189] ^ x[55];
  assign t[162] = t[190] ^ x[57];
  assign t[163] = t[191] ^ x[60];
  assign t[164] = t[192] ^ x[61];
  assign t[165] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[166] = (x[0]);
  assign t[167] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[168] = (x[9]);
  assign t[169] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[16] = t[18] ? x[16] : x[15];
  assign t[170] = (x[17]);
  assign t[171] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[172] = (x[23]);
  assign t[173] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[174] = (x[29]);
  assign t[175] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[176] = (x[32]);
  assign t[177] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[178] = (x[35]);
  assign t[179] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = ~(t[19] & t[20]);
  assign t[180] = (x[38]);
  assign t[181] = (x[1]);
  assign t[182] = (x[10]);
  assign t[183] = (x[24]);
  assign t[184] = (x[18]);
  assign t[185] = (x[2]);
  assign t[186] = (x[11]);
  assign t[187] = (x[25]);
  assign t[188] = (x[19]);
  assign t[189] = (x[3]);
  assign t[18] = ~(t[21]);
  assign t[190] = (x[12]);
  assign t[191] = (x[26]);
  assign t[192] = (x[20]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[83]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[26] | t[28]);
  assign t[24] = ~(t[29]);
  assign t[25] = ~(t[30] | t[31]);
  assign t[26] = ~(t[83]);
  assign t[27] = t[81] ? t[33] : t[32];
  assign t[28] = t[81] ? t[35] : t[34];
  assign t[29] = ~(t[36] | t[37]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[26]);
  assign t[31] = t[81] ? t[38] : t[34];
  assign t[32] = ~(t[39] & t[40]);
  assign t[33] = ~(t[41] & t[40]);
  assign t[34] = ~(x[7] & t[42]);
  assign t[35] = ~(t[43] & t[40]);
  assign t[36] = ~(t[30] | t[44]);
  assign t[37] = ~(t[30] | t[45]);
  assign t[38] = ~(t[84] & t[43]);
  assign t[39] = x[7] & t[82];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[84]);
  assign t[41] = ~(x[7] | t[82]);
  assign t[42] = ~(t[82] | t[84]);
  assign t[43] = ~(x[7] | t[46]);
  assign t[44] = t[81] ? t[47] : t[35];
  assign t[45] = t[81] ? t[32] : t[48];
  assign t[46] = ~(t[82]);
  assign t[47] = ~(x[7] & t[49]);
  assign t[48] = ~(t[41] & t[84]);
  assign t[49] = ~(t[82] | t[40]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[1] ? t[51] : t[85];
  assign t[51] = x[6] ? t[53] : t[52];
  assign t[52] = x[7] ? t[55] : t[54];
  assign t[53] = t[56] ^ x[42];
  assign t[54] = t[57] ^ t[55];
  assign t[55] = ~(t[86] ^ t[58]);
  assign t[56] = x[44] ^ x[45];
  assign t[57] = t[18] ? x[45] : x[44];
  assign t[58] = ~(t[87] ^ t[88]);
  assign t[59] = t[1] ? t[60] : t[89];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = x[6] ? t[62] : t[61];
  assign t[61] = x[7] ? t[64] : t[63];
  assign t[62] = t[65] ^ x[49];
  assign t[63] = t[66] ^ t[64];
  assign t[64] = ~(t[90] ^ t[67]);
  assign t[65] = x[51] ^ x[52];
  assign t[66] = t[18] ? x[52] : x[51];
  assign t[67] = ~(t[91] ^ t[92]);
  assign t[68] = t[1] ? t[69] : t[93];
  assign t[69] = x[6] ? t[71] : t[70];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = x[7] ? t[73] : t[72];
  assign t[71] = t[74] ^ x[56];
  assign t[72] = t[75] ^ t[73];
  assign t[73] = ~(t[94] ^ t[76]);
  assign t[74] = x[58] ^ x[59];
  assign t[75] = t[18] ? x[59] : x[58];
  assign t[76] = ~(t[95] ^ t[96]);
  assign t[77] = (t[97]);
  assign t[78] = (t[98]);
  assign t[79] = (t[99]);
  assign t[7] = ~(t[8] ^ t[12]);
  assign t[80] = (t[100]);
  assign t[81] = (t[101]);
  assign t[82] = (t[102]);
  assign t[83] = (t[103]);
  assign t[84] = (t[104]);
  assign t[85] = (t[105]);
  assign t[86] = (t[106]);
  assign t[87] = (t[107]);
  assign t[88] = (t[108]);
  assign t[89] = (t[109]);
  assign t[8] = ~(t[78] ^ t[13]);
  assign t[90] = (t[110]);
  assign t[91] = (t[111]);
  assign t[92] = (t[112]);
  assign t[93] = (t[113]);
  assign t[94] = (t[114]);
  assign t[95] = (t[115]);
  assign t[96] = (t[116]);
  assign t[97] = t[117] ^ x[5];
  assign t[98] = t[118] ^ x[14];
  assign t[99] = t[119] ^ x[22];
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0] & ~t[50] & ~t[59] & ~t[68]) | (~t[0] & t[50] & ~t[59] & ~t[68]) | (~t[0] & ~t[50] & t[59] & ~t[68]) | (~t[0] & ~t[50] & ~t[59] & t[68]) | (t[0] & t[50] & t[59] & ~t[68]) | (t[0] & t[50] & ~t[59] & t[68]) | (t[0] & ~t[50] & t[59] & t[68]) | (~t[0] & t[50] & t[59] & t[68]);
endmodule

module R2ind186(x, y);
 input [40:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[16] ? x[16] : x[15];
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[14] = ~(t[22] & t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[24]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[14];
  assign t[28] = t[36] ^ x[22];
  assign t[29] = t[37] ^ x[28];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[38] ^ x[31];
  assign t[31] = t[39] ^ x[34];
  assign t[32] = t[40] ^ x[37];
  assign t[33] = t[41] ^ x[40];
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[46] & t[47]);
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = t[58] ^ x[4];
  assign t[43] = t[59] ^ x[5];
  assign t[44] = t[60] ^ x[13];
  assign t[45] = t[61] ^ x[14];
  assign t[46] = t[62] ^ x[21];
  assign t[47] = t[63] ^ x[22];
  assign t[48] = t[64] ^ x[27];
  assign t[49] = t[65] ^ x[28];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[66] ^ x[30];
  assign t[51] = t[67] ^ x[31];
  assign t[52] = t[68] ^ x[33];
  assign t[53] = t[69] ^ x[34];
  assign t[54] = t[70] ^ x[36];
  assign t[55] = t[71] ^ x[37];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[40];
  assign t[58] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[59] = (x[3]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[61] = (x[12]);
  assign t[62] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[63] = (x[20]);
  assign t[64] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[65] = (x[26]);
  assign t[66] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[29]);
  assign t[68] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[32]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[35]);
  assign t[72] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[38]);
  assign t[7] = t[12] ^ t[8];
  assign t[8] = ~(t[19] ^ t[13]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [40:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[16] ? x[16] : x[15];
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[14] = ~(t[22] & t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[24]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[14];
  assign t[28] = t[36] ^ x[22];
  assign t[29] = t[37] ^ x[28];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[38] ^ x[31];
  assign t[31] = t[39] ^ x[34];
  assign t[32] = t[40] ^ x[37];
  assign t[33] = t[41] ^ x[40];
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[46] & t[47]);
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = t[58] ^ x[4];
  assign t[43] = t[59] ^ x[5];
  assign t[44] = t[60] ^ x[13];
  assign t[45] = t[61] ^ x[14];
  assign t[46] = t[62] ^ x[21];
  assign t[47] = t[63] ^ x[22];
  assign t[48] = t[64] ^ x[27];
  assign t[49] = t[65] ^ x[28];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[66] ^ x[30];
  assign t[51] = t[67] ^ x[31];
  assign t[52] = t[68] ^ x[33];
  assign t[53] = t[69] ^ x[34];
  assign t[54] = t[70] ^ x[36];
  assign t[55] = t[71] ^ x[37];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[40];
  assign t[58] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[59] = (x[2]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[61] = (x[11]);
  assign t[62] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[63] = (x[19]);
  assign t[64] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[65] = (x[25]);
  assign t[66] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[29]);
  assign t[68] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[32]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[35]);
  assign t[72] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[38]);
  assign t[7] = t[12] ^ t[8];
  assign t[8] = ~(t[19] ^ t[13]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [40:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = t[1] ? t[2] : t[18];
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(x[6]);
  assign t[12] = t[16] ? x[16] : x[15];
  assign t[13] = ~(t[20] ^ t[21]);
  assign t[14] = ~(t[22] & t[23]);
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[17]);
  assign t[17] = ~(t[24]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = t[34] ^ x[5];
  assign t[27] = t[35] ^ x[14];
  assign t[28] = t[36] ^ x[22];
  assign t[29] = t[37] ^ x[28];
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = t[38] ^ x[31];
  assign t[31] = t[39] ^ x[34];
  assign t[32] = t[40] ^ x[37];
  assign t[33] = t[41] ^ x[40];
  assign t[34] = (~t[42] & t[43]);
  assign t[35] = (~t[44] & t[45]);
  assign t[36] = (~t[46] & t[47]);
  assign t[37] = (~t[48] & t[49]);
  assign t[38] = (~t[50] & t[51]);
  assign t[39] = (~t[52] & t[53]);
  assign t[3] = ~(t[6]);
  assign t[40] = (~t[54] & t[55]);
  assign t[41] = (~t[56] & t[57]);
  assign t[42] = t[58] ^ x[4];
  assign t[43] = t[59] ^ x[5];
  assign t[44] = t[60] ^ x[13];
  assign t[45] = t[61] ^ x[14];
  assign t[46] = t[62] ^ x[21];
  assign t[47] = t[63] ^ x[22];
  assign t[48] = t[64] ^ x[27];
  assign t[49] = t[65] ^ x[28];
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = t[66] ^ x[30];
  assign t[51] = t[67] ^ x[31];
  assign t[52] = t[68] ^ x[33];
  assign t[53] = t[69] ^ x[34];
  assign t[54] = t[70] ^ x[36];
  assign t[55] = t[71] ^ x[37];
  assign t[56] = t[72] ^ x[39];
  assign t[57] = t[73] ^ x[40];
  assign t[58] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[59] = (x[1]);
  assign t[5] = t[9] ^ x[8];
  assign t[60] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[61] = (x[10]);
  assign t[62] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[63] = (x[18]);
  assign t[64] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[65] = (x[24]);
  assign t[66] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[29]);
  assign t[68] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[32]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[35]);
  assign t[72] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[38]);
  assign t[7] = t[12] ^ t[8];
  assign t[8] = ~(t[19] ^ t[13]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [40:0] x;
 output y;

 wire [105:0] t;
  assign t[0] = t[1] ? t[2] : t[50];
  assign t[100] = (x[32] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[32] & 1'b0 & ~1'b0 & ~1'b0) | (~x[32] & ~1'b0 & 1'b0 & ~1'b0) | (~x[32] & ~1'b0 & ~1'b0 & 1'b0) | (x[32] & 1'b0 & 1'b0 & ~1'b0) | (x[32] & 1'b0 & ~1'b0 & 1'b0) | (x[32] & ~1'b0 & 1'b0 & 1'b0) | (~x[32] & 1'b0 & 1'b0 & 1'b0);
  assign t[101] = (x[32]);
  assign t[102] = (x[35] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[35] & 1'b0 & ~1'b0 & ~1'b0) | (~x[35] & ~1'b0 & 1'b0 & ~1'b0) | (~x[35] & ~1'b0 & ~1'b0 & 1'b0) | (x[35] & 1'b0 & 1'b0 & ~1'b0) | (x[35] & 1'b0 & ~1'b0 & 1'b0) | (x[35] & ~1'b0 & 1'b0 & 1'b0) | (~x[35] & 1'b0 & 1'b0 & 1'b0);
  assign t[103] = (x[35]);
  assign t[104] = (x[38] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[38] & 1'b0 & ~1'b0 & ~1'b0) | (~x[38] & ~1'b0 & 1'b0 & ~1'b0) | (~x[38] & ~1'b0 & ~1'b0 & 1'b0) | (x[38] & 1'b0 & 1'b0 & ~1'b0) | (x[38] & 1'b0 & ~1'b0 & 1'b0) | (x[38] & ~1'b0 & 1'b0 & 1'b0) | (~x[38] & 1'b0 & 1'b0 & 1'b0);
  assign t[105] = (x[38]);
  assign t[10] = ~(t[14] | t[15]);
  assign t[11] = ~(x[6]);
  assign t[12] = ~(t[16] ^ t[17]);
  assign t[13] = ~(t[52] ^ t[53]);
  assign t[14] = ~(t[54] & t[55]);
  assign t[15] = ~(t[56] & t[57]);
  assign t[16] = t[18] ? x[16] : x[15];
  assign t[17] = ~(t[19] & t[20]);
  assign t[18] = ~(t[21]);
  assign t[19] = ~(t[22] | t[23]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[24] | t[25]);
  assign t[21] = ~(t[56]);
  assign t[22] = ~(t[26] | t[27]);
  assign t[23] = ~(t[26] | t[28]);
  assign t[24] = ~(t[29]);
  assign t[25] = ~(t[30] | t[31]);
  assign t[26] = ~(t[56]);
  assign t[27] = t[54] ? t[33] : t[32];
  assign t[28] = t[54] ? t[35] : t[34];
  assign t[29] = ~(t[36] | t[37]);
  assign t[2] = x[6] ? t[5] : t[4];
  assign t[30] = ~(t[26]);
  assign t[31] = t[54] ? t[38] : t[34];
  assign t[32] = ~(t[39] & t[40]);
  assign t[33] = ~(t[41] & t[40]);
  assign t[34] = ~(x[7] & t[42]);
  assign t[35] = ~(t[43] & t[40]);
  assign t[36] = ~(t[30] | t[44]);
  assign t[37] = ~(t[30] | t[45]);
  assign t[38] = ~(t[57] & t[43]);
  assign t[39] = x[7] & t[55];
  assign t[3] = ~(t[6]);
  assign t[40] = ~(t[57]);
  assign t[41] = ~(x[7] | t[55]);
  assign t[42] = ~(t[55] | t[57]);
  assign t[43] = ~(x[7] | t[46]);
  assign t[44] = t[54] ? t[47] : t[35];
  assign t[45] = t[54] ? t[32] : t[48];
  assign t[46] = ~(t[55]);
  assign t[47] = ~(x[7] & t[49]);
  assign t[48] = ~(t[41] & t[57]);
  assign t[49] = ~(t[55] | t[40]);
  assign t[4] = x[7] ? t[8] : t[7];
  assign t[50] = (t[58]);
  assign t[51] = (t[59]);
  assign t[52] = (t[60]);
  assign t[53] = (t[61]);
  assign t[54] = (t[62]);
  assign t[55] = (t[63]);
  assign t[56] = (t[64]);
  assign t[57] = (t[65]);
  assign t[58] = t[66] ^ x[5];
  assign t[59] = t[67] ^ x[14];
  assign t[5] = t[9] ^ x[8];
  assign t[60] = t[68] ^ x[22];
  assign t[61] = t[69] ^ x[28];
  assign t[62] = t[70] ^ x[31];
  assign t[63] = t[71] ^ x[34];
  assign t[64] = t[72] ^ x[37];
  assign t[65] = t[73] ^ x[40];
  assign t[66] = (~t[74] & t[75]);
  assign t[67] = (~t[76] & t[77]);
  assign t[68] = (~t[78] & t[79]);
  assign t[69] = (~t[80] & t[81]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (~t[82] & t[83]);
  assign t[71] = (~t[84] & t[85]);
  assign t[72] = (~t[86] & t[87]);
  assign t[73] = (~t[88] & t[89]);
  assign t[74] = t[90] ^ x[4];
  assign t[75] = t[91] ^ x[5];
  assign t[76] = t[92] ^ x[13];
  assign t[77] = t[93] ^ x[14];
  assign t[78] = t[94] ^ x[21];
  assign t[79] = t[95] ^ x[22];
  assign t[7] = ~(t[8] ^ t[12]);
  assign t[80] = t[96] ^ x[27];
  assign t[81] = t[97] ^ x[28];
  assign t[82] = t[98] ^ x[30];
  assign t[83] = t[99] ^ x[31];
  assign t[84] = t[100] ^ x[33];
  assign t[85] = t[101] ^ x[34];
  assign t[86] = t[102] ^ x[36];
  assign t[87] = t[103] ^ x[37];
  assign t[88] = t[104] ^ x[39];
  assign t[89] = t[105] ^ x[40];
  assign t[8] = ~(t[51] ^ t[13]);
  assign t[90] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[91] = (x[0]);
  assign t[92] = (x[9] & ~x[10] & ~x[11] & ~x[12]) | (~x[9] & x[10] & ~x[11] & ~x[12]) | (~x[9] & ~x[10] & x[11] & ~x[12]) | (~x[9] & ~x[10] & ~x[11] & x[12]) | (x[9] & x[10] & x[11] & ~x[12]) | (x[9] & x[10] & ~x[11] & x[12]) | (x[9] & ~x[10] & x[11] & x[12]) | (~x[9] & x[10] & x[11] & x[12]);
  assign t[93] = (x[9]);
  assign t[94] = (x[17] & ~x[18] & ~x[19] & ~x[20]) | (~x[17] & x[18] & ~x[19] & ~x[20]) | (~x[17] & ~x[18] & x[19] & ~x[20]) | (~x[17] & ~x[18] & ~x[19] & x[20]) | (x[17] & x[18] & x[19] & ~x[20]) | (x[17] & x[18] & ~x[19] & x[20]) | (x[17] & ~x[18] & x[19] & x[20]) | (~x[17] & x[18] & x[19] & x[20]);
  assign t[95] = (x[17]);
  assign t[96] = (x[23] & ~x[24] & ~x[25] & ~x[26]) | (~x[23] & x[24] & ~x[25] & ~x[26]) | (~x[23] & ~x[24] & x[25] & ~x[26]) | (~x[23] & ~x[24] & ~x[25] & x[26]) | (x[23] & x[24] & x[25] & ~x[26]) | (x[23] & x[24] & ~x[25] & x[26]) | (x[23] & ~x[24] & x[25] & x[26]) | (~x[23] & x[24] & x[25] & x[26]);
  assign t[97] = (x[23]);
  assign t[98] = (x[29] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[29] & 1'b0 & ~1'b0 & ~1'b0) | (~x[29] & ~1'b0 & 1'b0 & ~1'b0) | (~x[29] & ~1'b0 & ~1'b0 & 1'b0) | (x[29] & 1'b0 & 1'b0 & ~1'b0) | (x[29] & 1'b0 & ~1'b0 & 1'b0) | (x[29] & ~1'b0 & 1'b0 & 1'b0) | (~x[29] & 1'b0 & 1'b0 & 1'b0);
  assign t[99] = (x[29]);
  assign t[9] = x[15] ^ x[16];
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind191(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind196(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind201(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind206(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind211(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind216(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind221(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind226(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind231(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind236(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind241(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind246(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind251(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind255(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind256(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind257(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind258(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind259(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind260(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind261(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind262(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind263(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind264(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind265(x, y);
 input [8:0] x;
 output y;

 wire [40:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[22] & t[11]);
  assign t[11] = ~(t[21] & t[3]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[4] & t[6]);
  assign t[14] = ~(t[15] & t[19]);
  assign t[15] = ~(t[16] & t[3]);
  assign t[16] = ~(t[22] & t[21]);
  assign t[17] = ~(t[13] & t[18]);
  assign t[18] = t[1] | t[19];
  assign t[19] = (t[23]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = (t[24]);
  assign t[21] = (t[25]);
  assign t[22] = (t[26]);
  assign t[23] = t[27] ^ x[5];
  assign t[24] = t[28] ^ x[6];
  assign t[25] = t[29] ^ x[7];
  assign t[26] = t[30] ^ x[8];
  assign t[27] = (~t[31] & t[32]);
  assign t[28] = (~t[31] & t[33]);
  assign t[29] = (~t[31] & t[34]);
  assign t[2] = ~(t[19] | t[5]);
  assign t[30] = (~t[31] & t[35]);
  assign t[31] = t[36] ^ x[4];
  assign t[32] = t[37] ^ x[5];
  assign t[33] = t[38] ^ x[6];
  assign t[34] = t[39] ^ x[7];
  assign t[35] = t[40] ^ x[8];
  assign t[36] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[37] = (x[1]);
  assign t[38] = (x[2]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[20]);
  assign t[40] = (x[0]);
  assign t[4] = ~(t[21]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[22]);
  assign t[7] = ~(t[20] | t[21]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[20] & t[4]);
  assign y = (t[0] & ~t[8] & ~t[12] & ~t[17]) | (~t[0] & t[8] & ~t[12] & ~t[17]) | (~t[0] & ~t[8] & t[12] & ~t[17]) | (~t[0] & ~t[8] & ~t[12] & t[17]) | (t[0] & t[8] & t[12] & ~t[17]) | (t[0] & t[8] & ~t[12] & t[17]) | (t[0] & ~t[8] & t[12] & t[17]) | (~t[0] & t[8] & t[12] & t[17]);
endmodule

module R2ind266(x, y);
 input [8:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[6];
  assign t[13] = t[17] ^ x[7];
  assign t[14] = t[18] ^ x[8];
  assign t[15] = (~t[19] & t[20]);
  assign t[16] = (~t[19] & t[21]);
  assign t[17] = (~t[19] & t[22]);
  assign t[18] = (~t[19] & t[23]);
  assign t[19] = t[24] ^ x[4];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[5];
  assign t[21] = t[26] ^ x[6];
  assign t[22] = t[27] ^ x[7];
  assign t[23] = t[28] ^ x[8];
  assign t[24] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[25] = (x[1]);
  assign t[26] = (x[3]);
  assign t[27] = (x[0]);
  assign t[28] = (x[2]);
  assign t[2] = t[5] | t[7];
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[9]);
  assign t[5] = ~(t[6] | t[3]);
  assign t[6] = ~(t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind267(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[3]);
  assign t[28] = (x[0]);
  assign t[29] = (x[2]);
  assign t[2] = ~(t[5] & t[8]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] & t[7]);
  assign t[6] = ~(t[10] & t[9]);
  assign t[7] = ~(t[11]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind268(x, y);
 input [7:0] x;
 output y;

 wire [22:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[13] ^ x[6];
  assign t[11] = t[14] ^ x[7];
  assign t[12] = (~t[15] & t[16]);
  assign t[13] = (~t[15] & t[17]);
  assign t[14] = (~t[15] & t[18]);
  assign t[15] = t[19] ^ x[4];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[6];
  assign t[18] = t[22] ^ x[7];
  assign t[19] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[1] = ~(t[6] & t[3]);
  assign t[20] = (x[2]);
  assign t[21] = (x[0]);
  assign t[22] = (x[3]);
  assign t[2] = ~(t[7] & t[4]);
  assign t[3] = ~(t[8]);
  assign t[4] = ~(t[8] & t[5]);
  assign t[5] = ~(t[6]);
  assign t[6] = (t[9]);
  assign t[7] = (t[10]);
  assign t[8] = (t[11]);
  assign t[9] = t[12] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind269(x, y);
 input [8:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = t[16] ^ x[5];
  assign t[13] = t[17] ^ x[6];
  assign t[14] = t[18] ^ x[7];
  assign t[15] = t[19] ^ x[8];
  assign t[16] = (~t[20] & t[21]);
  assign t[17] = (~t[20] & t[22]);
  assign t[18] = (~t[20] & t[23]);
  assign t[19] = (~t[20] & t[24]);
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[25] ^ x[4];
  assign t[21] = t[26] ^ x[5];
  assign t[22] = t[27] ^ x[6];
  assign t[23] = t[28] ^ x[7];
  assign t[24] = t[29] ^ x[8];
  assign t[25] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[26] = (x[1]);
  assign t[27] = (x[2]);
  assign t[28] = (x[3]);
  assign t[29] = (x[0]);
  assign t[2] = ~(t[8] | t[5]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[11]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = (t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind270(x, y);
 input [29:0] x;
 output y;

 wire [94:0] t;
  assign t[0] = ~(t[45] ^ t[1]);
  assign t[10] = ~(t[16]);
  assign t[11] = t[47] ? t[18] : t[17];
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = t[47] ? t[24] : t[23];
  assign t[15] = t[47] ? t[26] : t[25];
  assign t[16] = ~(t[46]);
  assign t[17] = ~(t[27] & t[48]);
  assign t[18] = ~(t[28] & t[29]);
  assign t[19] = ~(t[10] | t[30]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[10] | t[31]);
  assign t[21] = t[48] & t[32];
  assign t[22] = t[28] | t[27];
  assign t[23] = ~(t[33] & t[29]);
  assign t[24] = ~(x[17] & t[34]);
  assign t[25] = ~(t[28] & t[48]);
  assign t[26] = ~(t[27] & t[29]);
  assign t[27] = x[17] & t[49];
  assign t[28] = ~(x[17] | t[49]);
  assign t[29] = ~(t[48]);
  assign t[2] = t[46] ? x[10] : x[9];
  assign t[30] = t[47] ? t[17] : t[18];
  assign t[31] = t[47] ? t[36] : t[35];
  assign t[32] = ~(t[16] | t[47]);
  assign t[33] = ~(x[17] | t[37]);
  assign t[34] = ~(t[49] | t[29]);
  assign t[35] = ~(t[48] & t[33]);
  assign t[36] = ~(x[17] & t[38]);
  assign t[37] = ~(t[49]);
  assign t[38] = ~(t[49] | t[48]);
  assign t[39] = t[40] ^ t[50];
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = t[46] ? x[23] : x[22];
  assign t[41] = t[42] ^ t[51];
  assign t[42] = t[46] ? x[26] : x[25];
  assign t[43] = t[44] ^ t[52];
  assign t[44] = t[46] ? x[29] : x[28];
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = (t[57]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[50] = (t[58]);
  assign t[51] = (t[59]);
  assign t[52] = (t[60]);
  assign t[53] = t[61] ^ x[5];
  assign t[54] = t[62] ^ x[8];
  assign t[55] = t[63] ^ x[13];
  assign t[56] = t[64] ^ x[16];
  assign t[57] = t[65] ^ x[20];
  assign t[58] = t[66] ^ x[21];
  assign t[59] = t[67] ^ x[24];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[68] ^ x[27];
  assign t[61] = (~t[69] & t[70]);
  assign t[62] = (~t[71] & t[72]);
  assign t[63] = (~t[73] & t[74]);
  assign t[64] = (~t[75] & t[76]);
  assign t[65] = (~t[77] & t[78]);
  assign t[66] = (~t[69] & t[79]);
  assign t[67] = (~t[69] & t[80]);
  assign t[68] = (~t[69] & t[81]);
  assign t[69] = t[82] ^ x[4];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[83] ^ x[5];
  assign t[71] = t[84] ^ x[7];
  assign t[72] = t[85] ^ x[8];
  assign t[73] = t[86] ^ x[12];
  assign t[74] = t[87] ^ x[13];
  assign t[75] = t[88] ^ x[15];
  assign t[76] = t[89] ^ x[16];
  assign t[77] = t[90] ^ x[19];
  assign t[78] = t[91] ^ x[20];
  assign t[79] = t[92] ^ x[21];
  assign t[7] = ~(t[12] & t[13]);
  assign t[80] = t[93] ^ x[24];
  assign t[81] = t[94] ^ x[27];
  assign t[82] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[83] = (x[0]);
  assign t[84] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[6]);
  assign t[86] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[11]);
  assign t[88] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[14]);
  assign t[8] = ~(t[10] | t[14]);
  assign t[90] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[18]);
  assign t[92] = (x[1]);
  assign t[93] = (x[2]);
  assign t[94] = (x[3]);
  assign t[9] = ~(t[10] | t[15]);
  assign y = (t[0] & ~t[39] & ~t[41] & ~t[43]) | (~t[0] & t[39] & ~t[41] & ~t[43]) | (~t[0] & ~t[39] & t[41] & ~t[43]) | (~t[0] & ~t[39] & ~t[41] & t[43]) | (t[0] & t[39] & t[41] & ~t[43]) | (t[0] & t[39] & ~t[41] & t[43]) | (t[0] & ~t[39] & t[41] & t[43]) | (~t[0] & t[39] & t[41] & t[43]);
endmodule

module R2ind271(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[3]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind272(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[2]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind273(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[1]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind274(x, y);
 input [20:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = ~(t[39] ^ t[1]);
  assign t[10] = ~(t[16]);
  assign t[11] = t[41] ? t[18] : t[17];
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = t[41] ? t[24] : t[23];
  assign t[15] = t[41] ? t[26] : t[25];
  assign t[16] = ~(t[40]);
  assign t[17] = ~(t[27] & t[42]);
  assign t[18] = ~(t[28] & t[29]);
  assign t[19] = ~(t[10] | t[30]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[10] | t[31]);
  assign t[21] = t[42] & t[32];
  assign t[22] = t[28] | t[27];
  assign t[23] = ~(t[33] & t[29]);
  assign t[24] = ~(x[17] & t[34]);
  assign t[25] = ~(t[28] & t[42]);
  assign t[26] = ~(t[27] & t[29]);
  assign t[27] = x[17] & t[43];
  assign t[28] = ~(x[17] | t[43]);
  assign t[29] = ~(t[42]);
  assign t[2] = t[40] ? x[10] : x[9];
  assign t[30] = t[41] ? t[17] : t[18];
  assign t[31] = t[41] ? t[36] : t[35];
  assign t[32] = ~(t[16] | t[41]);
  assign t[33] = ~(x[17] | t[37]);
  assign t[34] = ~(t[43] | t[29]);
  assign t[35] = ~(t[42] & t[33]);
  assign t[36] = ~(x[17] & t[38]);
  assign t[37] = ~(t[43]);
  assign t[38] = ~(t[43] | t[42]);
  assign t[39] = (t[44]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = (t[48]);
  assign t[44] = t[49] ^ x[5];
  assign t[45] = t[50] ^ x[8];
  assign t[46] = t[51] ^ x[13];
  assign t[47] = t[52] ^ x[16];
  assign t[48] = t[53] ^ x[20];
  assign t[49] = (~t[54] & t[55]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[50] = (~t[56] & t[57]);
  assign t[51] = (~t[58] & t[59]);
  assign t[52] = (~t[60] & t[61]);
  assign t[53] = (~t[62] & t[63]);
  assign t[54] = t[64] ^ x[4];
  assign t[55] = t[65] ^ x[5];
  assign t[56] = t[66] ^ x[7];
  assign t[57] = t[67] ^ x[8];
  assign t[58] = t[68] ^ x[12];
  assign t[59] = t[69] ^ x[13];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[15];
  assign t[61] = t[71] ^ x[16];
  assign t[62] = t[72] ^ x[19];
  assign t[63] = t[73] ^ x[20];
  assign t[64] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[65] = (x[0]);
  assign t[66] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[6]);
  assign t[68] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[11]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[14]);
  assign t[72] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[18]);
  assign t[7] = ~(t[12] & t[13]);
  assign t[8] = ~(t[10] | t[14]);
  assign t[9] = ~(t[10] | t[15]);
  assign y = (t[0]);
endmodule

module R2ind275(x, y);
 input [29:0] x;
 output y;

 wire [102:0] t;
  assign t[0] = ~(t[53] ^ t[1]);
  assign t[100] = (x[1]);
  assign t[101] = (x[2]);
  assign t[102] = (x[3]);
  assign t[10] = ~(t[14]);
  assign t[11] = t[55] ? t[19] : t[18];
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[54]);
  assign t[15] = t[55] ? t[25] : t[24];
  assign t[16] = ~(t[10] | t[26]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[28] & t[56]);
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[10] | t[31]);
  assign t[21] = ~(t[10] | t[32]);
  assign t[22] = t[56] & t[33];
  assign t[23] = t[29] | t[28];
  assign t[24] = ~(x[17] & t[34]);
  assign t[25] = ~(t[35] & t[30]);
  assign t[26] = t[55] ? t[37] : t[36];
  assign t[27] = ~(t[33] & t[38]);
  assign t[28] = x[17] & t[57];
  assign t[29] = ~(x[17] | t[57]);
  assign t[2] = t[54] ? x[10] : x[9];
  assign t[30] = ~(t[56]);
  assign t[31] = t[55] ? t[18] : t[19];
  assign t[32] = t[55] ? t[24] : t[39];
  assign t[33] = ~(t[14] | t[55]);
  assign t[34] = ~(t[57] | t[56]);
  assign t[35] = ~(x[17] | t[40]);
  assign t[36] = ~(t[28] & t[30]);
  assign t[37] = ~(t[29] & t[56]);
  assign t[38] = ~(t[39] & t[41]);
  assign t[39] = ~(t[56] & t[35]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = ~(t[57]);
  assign t[41] = ~(x[17] & t[42]);
  assign t[42] = ~(t[57] | t[30]);
  assign t[43] = t[44] ^ t[58];
  assign t[44] = t[45] ? x[23] : x[22];
  assign t[45] = ~(t[46]);
  assign t[46] = ~(t[54]);
  assign t[47] = t[48] ^ t[59];
  assign t[48] = t[49] ? x[26] : x[25];
  assign t[49] = ~(t[46]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[50] = t[51] ^ t[60];
  assign t[51] = t[52] ? x[29] : x[28];
  assign t[52] = ~(t[46]);
  assign t[53] = (t[61]);
  assign t[54] = (t[62]);
  assign t[55] = (t[63]);
  assign t[56] = (t[64]);
  assign t[57] = (t[65]);
  assign t[58] = (t[66]);
  assign t[59] = (t[67]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (t[68]);
  assign t[61] = t[69] ^ x[5];
  assign t[62] = t[70] ^ x[8];
  assign t[63] = t[71] ^ x[13];
  assign t[64] = t[72] ^ x[16];
  assign t[65] = t[73] ^ x[20];
  assign t[66] = t[74] ^ x[21];
  assign t[67] = t[75] ^ x[24];
  assign t[68] = t[76] ^ x[27];
  assign t[69] = (~t[77] & t[78]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (~t[79] & t[80]);
  assign t[71] = (~t[81] & t[82]);
  assign t[72] = (~t[83] & t[84]);
  assign t[73] = (~t[85] & t[86]);
  assign t[74] = (~t[77] & t[87]);
  assign t[75] = (~t[77] & t[88]);
  assign t[76] = (~t[77] & t[89]);
  assign t[77] = t[90] ^ x[4];
  assign t[78] = t[91] ^ x[5];
  assign t[79] = t[92] ^ x[7];
  assign t[7] = ~(t[12] & t[13]);
  assign t[80] = t[93] ^ x[8];
  assign t[81] = t[94] ^ x[12];
  assign t[82] = t[95] ^ x[13];
  assign t[83] = t[96] ^ x[15];
  assign t[84] = t[97] ^ x[16];
  assign t[85] = t[98] ^ x[19];
  assign t[86] = t[99] ^ x[20];
  assign t[87] = t[100] ^ x[21];
  assign t[88] = t[101] ^ x[24];
  assign t[89] = t[102] ^ x[27];
  assign t[8] = ~(t[14] | t[15]);
  assign t[90] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[91] = (x[0]);
  assign t[92] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[6]);
  assign t[94] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[95] = (x[11]);
  assign t[96] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[97] = (x[14]);
  assign t[98] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[99] = (x[18]);
  assign t[9] = t[16] | t[17];
  assign y = (t[0] & ~t[43] & ~t[47] & ~t[50]) | (~t[0] & t[43] & ~t[47] & ~t[50]) | (~t[0] & ~t[43] & t[47] & ~t[50]) | (~t[0] & ~t[43] & ~t[47] & t[50]) | (t[0] & t[43] & t[47] & ~t[50]) | (t[0] & t[43] & ~t[47] & t[50]) | (t[0] & ~t[43] & t[47] & t[50]) | (~t[0] & t[43] & t[47] & t[50]);
endmodule

module R2ind276(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind277(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind278(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind279(x, y);
 input [20:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[43] ^ t[1]);
  assign t[10] = ~(t[14]);
  assign t[11] = t[45] ? t[19] : t[18];
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[44]);
  assign t[15] = t[45] ? t[25] : t[24];
  assign t[16] = ~(t[10] | t[26]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[28] & t[46]);
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[10] | t[31]);
  assign t[21] = ~(t[10] | t[32]);
  assign t[22] = t[46] & t[33];
  assign t[23] = t[29] | t[28];
  assign t[24] = ~(x[17] & t[34]);
  assign t[25] = ~(t[35] & t[30]);
  assign t[26] = t[45] ? t[37] : t[36];
  assign t[27] = ~(t[33] & t[38]);
  assign t[28] = x[17] & t[47];
  assign t[29] = ~(x[17] | t[47]);
  assign t[2] = t[44] ? x[10] : x[9];
  assign t[30] = ~(t[46]);
  assign t[31] = t[45] ? t[18] : t[19];
  assign t[32] = t[45] ? t[24] : t[39];
  assign t[33] = ~(t[14] | t[45]);
  assign t[34] = ~(t[47] | t[46]);
  assign t[35] = ~(x[17] | t[40]);
  assign t[36] = ~(t[28] & t[30]);
  assign t[37] = ~(t[29] & t[46]);
  assign t[38] = ~(t[39] & t[41]);
  assign t[39] = ~(t[46] & t[35]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[40] = ~(t[47]);
  assign t[41] = ~(x[17] & t[42]);
  assign t[42] = ~(t[47] | t[30]);
  assign t[43] = (t[48]);
  assign t[44] = (t[49]);
  assign t[45] = (t[50]);
  assign t[46] = (t[51]);
  assign t[47] = (t[52]);
  assign t[48] = t[53] ^ x[5];
  assign t[49] = t[54] ^ x[8];
  assign t[4] = ~(t[6] | t[7]);
  assign t[50] = t[55] ^ x[13];
  assign t[51] = t[56] ^ x[16];
  assign t[52] = t[57] ^ x[20];
  assign t[53] = (~t[58] & t[59]);
  assign t[54] = (~t[60] & t[61]);
  assign t[55] = (~t[62] & t[63]);
  assign t[56] = (~t[64] & t[65]);
  assign t[57] = (~t[66] & t[67]);
  assign t[58] = t[68] ^ x[4];
  assign t[59] = t[69] ^ x[5];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[7];
  assign t[61] = t[71] ^ x[8];
  assign t[62] = t[72] ^ x[12];
  assign t[63] = t[73] ^ x[13];
  assign t[64] = t[74] ^ x[15];
  assign t[65] = t[75] ^ x[16];
  assign t[66] = t[76] ^ x[19];
  assign t[67] = t[77] ^ x[20];
  assign t[68] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[69] = (x[0]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[6]);
  assign t[72] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[11]);
  assign t[74] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[14]);
  assign t[76] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[18]);
  assign t[7] = ~(t[12] & t[13]);
  assign t[8] = ~(t[14] | t[15]);
  assign t[9] = t[16] | t[17];
  assign y = (t[0]);
endmodule

module R2ind280(x, y);
 input [29:0] x;
 output y;

 wire [92:0] t;
  assign t[0] = ~(t[43] ^ t[1]);
  assign t[10] = ~(t[18] | t[45]);
  assign t[11] = ~(t[19] & t[20]);
  assign t[12] = ~(t[46] | t[21]);
  assign t[13] = t[22] & t[45];
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = ~(t[22] | t[24]);
  assign t[16] = ~(t[22] | t[25]);
  assign t[17] = ~(t[22] | t[26]);
  assign t[18] = ~(t[44]);
  assign t[19] = ~(t[47] & t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(x[20] & t[12]);
  assign t[21] = ~(t[47]);
  assign t[22] = ~(t[18]);
  assign t[23] = t[45] ? t[29] : t[28];
  assign t[24] = t[45] ? t[31] : t[30];
  assign t[25] = t[45] ? t[32] : t[19];
  assign t[26] = t[45] ? t[30] : t[31];
  assign t[27] = ~(x[20] | t[33]);
  assign t[28] = ~(t[34] & t[47]);
  assign t[29] = ~(t[35] & t[21]);
  assign t[2] = t[44] ? x[10] : x[9];
  assign t[30] = ~(t[34] & t[21]);
  assign t[31] = ~(t[35] & t[47]);
  assign t[32] = ~(x[20] & t[36]);
  assign t[33] = ~(t[46]);
  assign t[34] = x[20] & t[46];
  assign t[35] = ~(x[20] | t[46]);
  assign t[36] = ~(t[46] | t[47]);
  assign t[37] = t[38] ^ t[48];
  assign t[38] = t[44] ? x[23] : x[22];
  assign t[39] = t[40] ^ t[49];
  assign t[3] = t[4] | t[5];
  assign t[40] = t[44] ? x[26] : x[25];
  assign t[41] = t[42] ^ t[50];
  assign t[42] = t[44] ? x[29] : x[28];
  assign t[43] = (t[51]);
  assign t[44] = (t[52]);
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = (t[57]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[50] = (t[58]);
  assign t[51] = t[59] ^ x[5];
  assign t[52] = t[60] ^ x[8];
  assign t[53] = t[61] ^ x[13];
  assign t[54] = t[62] ^ x[16];
  assign t[55] = t[63] ^ x[19];
  assign t[56] = t[64] ^ x[21];
  assign t[57] = t[65] ^ x[24];
  assign t[58] = t[66] ^ x[27];
  assign t[59] = (~t[67] & t[68]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (~t[69] & t[70]);
  assign t[61] = (~t[71] & t[72]);
  assign t[62] = (~t[73] & t[74]);
  assign t[63] = (~t[75] & t[76]);
  assign t[64] = (~t[67] & t[77]);
  assign t[65] = (~t[67] & t[78]);
  assign t[66] = (~t[67] & t[79]);
  assign t[67] = t[80] ^ x[4];
  assign t[68] = t[81] ^ x[5];
  assign t[69] = t[82] ^ x[7];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[83] ^ x[8];
  assign t[71] = t[84] ^ x[12];
  assign t[72] = t[85] ^ x[13];
  assign t[73] = t[86] ^ x[15];
  assign t[74] = t[87] ^ x[16];
  assign t[75] = t[88] ^ x[18];
  assign t[76] = t[89] ^ x[19];
  assign t[77] = t[90] ^ x[21];
  assign t[78] = t[91] ^ x[24];
  assign t[79] = t[92] ^ x[27];
  assign t[7] = ~(t[12] & t[13]);
  assign t[80] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[81] = (x[0]);
  assign t[82] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[6]);
  assign t[84] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[11]);
  assign t[86] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[14]);
  assign t[88] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[17]);
  assign t[8] = ~(t[14] | t[15]);
  assign t[90] = (x[1]);
  assign t[91] = (x[2]);
  assign t[92] = (x[3]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = (t[0] & ~t[37] & ~t[39] & ~t[41]) | (~t[0] & t[37] & ~t[39] & ~t[41]) | (~t[0] & ~t[37] & t[39] & ~t[41]) | (~t[0] & ~t[37] & ~t[39] & t[41]) | (t[0] & t[37] & t[39] & ~t[41]) | (t[0] & t[37] & ~t[39] & t[41]) | (t[0] & ~t[37] & t[39] & t[41]) | (~t[0] & t[37] & t[39] & t[41]);
endmodule

module R2ind281(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[3]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind282(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[2]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind283(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[1]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind284(x, y);
 input [20:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[37] ^ t[1]);
  assign t[10] = ~(t[18] | t[39]);
  assign t[11] = ~(t[19] & t[20]);
  assign t[12] = ~(t[40] | t[21]);
  assign t[13] = t[22] & t[39];
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = ~(t[22] | t[24]);
  assign t[16] = ~(t[22] | t[25]);
  assign t[17] = ~(t[22] | t[26]);
  assign t[18] = ~(t[38]);
  assign t[19] = ~(t[41] & t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(x[20] & t[12]);
  assign t[21] = ~(t[41]);
  assign t[22] = ~(t[18]);
  assign t[23] = t[39] ? t[29] : t[28];
  assign t[24] = t[39] ? t[31] : t[30];
  assign t[25] = t[39] ? t[32] : t[19];
  assign t[26] = t[39] ? t[30] : t[31];
  assign t[27] = ~(x[20] | t[33]);
  assign t[28] = ~(t[34] & t[41]);
  assign t[29] = ~(t[35] & t[21]);
  assign t[2] = t[38] ? x[10] : x[9];
  assign t[30] = ~(t[34] & t[21]);
  assign t[31] = ~(t[35] & t[41]);
  assign t[32] = ~(x[20] & t[36]);
  assign t[33] = ~(t[40]);
  assign t[34] = x[20] & t[40];
  assign t[35] = ~(x[20] | t[40]);
  assign t[36] = ~(t[40] | t[41]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = t[4] | t[5];
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = t[47] ^ x[5];
  assign t[43] = t[48] ^ x[8];
  assign t[44] = t[49] ^ x[13];
  assign t[45] = t[50] ^ x[16];
  assign t[46] = t[51] ^ x[19];
  assign t[47] = (~t[52] & t[53]);
  assign t[48] = (~t[54] & t[55]);
  assign t[49] = (~t[56] & t[57]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[50] = (~t[58] & t[59]);
  assign t[51] = (~t[60] & t[61]);
  assign t[52] = t[62] ^ x[4];
  assign t[53] = t[63] ^ x[5];
  assign t[54] = t[64] ^ x[7];
  assign t[55] = t[65] ^ x[8];
  assign t[56] = t[66] ^ x[12];
  assign t[57] = t[67] ^ x[13];
  assign t[58] = t[68] ^ x[15];
  assign t[59] = t[69] ^ x[16];
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[70] ^ x[18];
  assign t[61] = t[71] ^ x[19];
  assign t[62] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[63] = (x[0]);
  assign t[64] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[6]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[11]);
  assign t[68] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[14]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[17]);
  assign t[7] = ~(t[12] & t[13]);
  assign t[8] = ~(t[14] | t[15]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = (t[0]);
endmodule

module R2ind285(x, y);
 input [29:0] x;
 output y;

 wire [92:0] t;
  assign t[0] = ~(t[43] ^ t[1]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[19] & t[20]);
  assign t[13] = ~(t[21]);
  assign t[14] = t[22] | t[23];
  assign t[15] = ~(t[22]);
  assign t[16] = t[45] ? t[25] : t[24];
  assign t[17] = ~(t[22] | t[45]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[46] | t[28]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[15] & t[45];
  assign t[21] = ~(t[22] | t[29]);
  assign t[22] = ~(t[44]);
  assign t[23] = t[45] ? t[31] : t[30];
  assign t[24] = ~(t[32] & t[47]);
  assign t[25] = ~(t[33] & t[28]);
  assign t[26] = ~(t[47] & t[34]);
  assign t[27] = ~(x[20] & t[19]);
  assign t[28] = ~(t[47]);
  assign t[29] = t[45] ? t[30] : t[31];
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[34] & t[28]);
  assign t[31] = ~(x[20] & t[35]);
  assign t[32] = x[20] & t[46];
  assign t[33] = ~(x[20] | t[46]);
  assign t[34] = ~(x[20] | t[36]);
  assign t[35] = ~(t[46] | t[47]);
  assign t[36] = ~(t[46]);
  assign t[37] = t[38] ^ t[48];
  assign t[38] = t[44] ? x[23] : x[22];
  assign t[39] = t[40] ^ t[49];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[44] ? x[26] : x[25];
  assign t[41] = t[42] ^ t[50];
  assign t[42] = t[44] ? x[29] : x[28];
  assign t[43] = (t[51]);
  assign t[44] = (t[52]);
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = (t[57]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[58]);
  assign t[51] = t[59] ^ x[5];
  assign t[52] = t[60] ^ x[10];
  assign t[53] = t[61] ^ x[13];
  assign t[54] = t[62] ^ x[16];
  assign t[55] = t[63] ^ x[19];
  assign t[56] = t[64] ^ x[21];
  assign t[57] = t[65] ^ x[24];
  assign t[58] = t[66] ^ x[27];
  assign t[59] = (~t[67] & t[68]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (~t[69] & t[70]);
  assign t[61] = (~t[71] & t[72]);
  assign t[62] = (~t[73] & t[74]);
  assign t[63] = (~t[75] & t[76]);
  assign t[64] = (~t[67] & t[77]);
  assign t[65] = (~t[67] & t[78]);
  assign t[66] = (~t[67] & t[79]);
  assign t[67] = t[80] ^ x[4];
  assign t[68] = t[81] ^ x[5];
  assign t[69] = t[82] ^ x[9];
  assign t[6] = ~(t[10]);
  assign t[70] = t[83] ^ x[10];
  assign t[71] = t[84] ^ x[12];
  assign t[72] = t[85] ^ x[13];
  assign t[73] = t[86] ^ x[15];
  assign t[74] = t[87] ^ x[16];
  assign t[75] = t[88] ^ x[18];
  assign t[76] = t[89] ^ x[19];
  assign t[77] = t[90] ^ x[21];
  assign t[78] = t[91] ^ x[24];
  assign t[79] = t[92] ^ x[27];
  assign t[7] = ~(t[44]);
  assign t[80] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[81] = (x[0]);
  assign t[82] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[8]);
  assign t[84] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[11]);
  assign t[86] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[14]);
  assign t[88] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[89] = (x[17]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[90] = (x[1]);
  assign t[91] = (x[2]);
  assign t[92] = (x[3]);
  assign t[9] = ~(t[13] & t[14]);
  assign y = (t[0] & ~t[37] & ~t[39] & ~t[41]) | (~t[0] & t[37] & ~t[39] & ~t[41]) | (~t[0] & ~t[37] & t[39] & ~t[41]) | (~t[0] & ~t[37] & ~t[39] & t[41]) | (t[0] & t[37] & t[39] & ~t[41]) | (t[0] & t[37] & ~t[39] & t[41]) | (t[0] & ~t[37] & t[39] & t[41]) | (~t[0] & t[37] & t[39] & t[41]);
endmodule

module R2ind286(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[3]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind287(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[2]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind288(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[1]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind289(x, y);
 input [20:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[37] ^ t[1]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[19] & t[20]);
  assign t[13] = ~(t[21]);
  assign t[14] = t[22] | t[23];
  assign t[15] = ~(t[22]);
  assign t[16] = t[39] ? t[25] : t[24];
  assign t[17] = ~(t[22] | t[39]);
  assign t[18] = ~(t[26] & t[27]);
  assign t[19] = ~(t[40] | t[28]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[15] & t[39];
  assign t[21] = ~(t[22] | t[29]);
  assign t[22] = ~(t[38]);
  assign t[23] = t[39] ? t[31] : t[30];
  assign t[24] = ~(t[32] & t[41]);
  assign t[25] = ~(t[33] & t[28]);
  assign t[26] = ~(t[41] & t[34]);
  assign t[27] = ~(x[20] & t[19]);
  assign t[28] = ~(t[41]);
  assign t[29] = t[39] ? t[30] : t[31];
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[34] & t[28]);
  assign t[31] = ~(x[20] & t[35]);
  assign t[32] = x[20] & t[40];
  assign t[33] = ~(x[20] | t[40]);
  assign t[34] = ~(x[20] | t[36]);
  assign t[35] = ~(t[40] | t[41]);
  assign t[36] = ~(t[40]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = t[47] ^ x[5];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = t[49] ^ x[13];
  assign t[45] = t[50] ^ x[16];
  assign t[46] = t[51] ^ x[19];
  assign t[47] = (~t[52] & t[53]);
  assign t[48] = (~t[54] & t[55]);
  assign t[49] = (~t[56] & t[57]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[58] & t[59]);
  assign t[51] = (~t[60] & t[61]);
  assign t[52] = t[62] ^ x[4];
  assign t[53] = t[63] ^ x[5];
  assign t[54] = t[64] ^ x[9];
  assign t[55] = t[65] ^ x[10];
  assign t[56] = t[66] ^ x[12];
  assign t[57] = t[67] ^ x[13];
  assign t[58] = t[68] ^ x[15];
  assign t[59] = t[69] ^ x[16];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[18];
  assign t[61] = t[71] ^ x[19];
  assign t[62] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[63] = (x[0]);
  assign t[64] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[8]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[11]);
  assign t[68] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[14]);
  assign t[6] = ~(t[10]);
  assign t[70] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[17]);
  assign t[7] = ~(t[38]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = ~(t[13] & t[14]);
  assign y = (t[0]);
endmodule

module R2ind290(x, y);
 input [29:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[51] ^ t[1]);
  assign t[100] = (x[3]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = ~(t[16] | t[18]);
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = t[21] | t[25];
  assign t[16] = ~(t[21]);
  assign t[17] = t[53] ? t[27] : t[26];
  assign t[18] = t[53] ? t[29] : t[28];
  assign t[19] = ~(t[21] | t[30]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[16] | t[31]);
  assign t[21] = ~(t[52]);
  assign t[22] = ~(t[32] & t[33]);
  assign t[23] = t[54] & t[34];
  assign t[24] = t[35] | t[36];
  assign t[25] = t[53] ? t[32] : t[37];
  assign t[26] = ~(t[35] & t[38]);
  assign t[27] = ~(t[36] & t[54]);
  assign t[28] = ~(t[35] & t[54]);
  assign t[29] = ~(t[36] & t[38]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[53] ? t[26] : t[29];
  assign t[31] = t[53] ? t[37] : t[39];
  assign t[32] = ~(x[17] & t[40]);
  assign t[33] = ~(t[54] & t[41]);
  assign t[34] = ~(t[21] | t[53]);
  assign t[35] = ~(x[17] | t[55]);
  assign t[36] = x[17] & t[55];
  assign t[37] = ~(t[41] & t[38]);
  assign t[38] = ~(t[54]);
  assign t[39] = ~(x[17] & t[42]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = ~(t[55] | t[54]);
  assign t[41] = ~(x[17] | t[43]);
  assign t[42] = ~(t[55] | t[38]);
  assign t[43] = ~(t[55]);
  assign t[44] = t[45] ^ t[56];
  assign t[45] = t[46] ? x[23] : x[22];
  assign t[46] = ~(t[7]);
  assign t[47] = t[48] ^ t[57];
  assign t[48] = t[4] ? x[26] : x[25];
  assign t[49] = t[50] ^ t[58];
  assign t[4] = ~(t[7]);
  assign t[50] = t[4] ? x[29] : x[28];
  assign t[51] = (t[59]);
  assign t[52] = (t[60]);
  assign t[53] = (t[61]);
  assign t[54] = (t[62]);
  assign t[55] = (t[63]);
  assign t[56] = (t[64]);
  assign t[57] = (t[65]);
  assign t[58] = (t[66]);
  assign t[59] = t[67] ^ x[5];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[68] ^ x[10];
  assign t[61] = t[69] ^ x[13];
  assign t[62] = t[70] ^ x[16];
  assign t[63] = t[71] ^ x[20];
  assign t[64] = t[72] ^ x[21];
  assign t[65] = t[73] ^ x[24];
  assign t[66] = t[74] ^ x[27];
  assign t[67] = (~t[75] & t[76]);
  assign t[68] = (~t[77] & t[78]);
  assign t[69] = (~t[79] & t[80]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (~t[81] & t[82]);
  assign t[71] = (~t[83] & t[84]);
  assign t[72] = (~t[75] & t[85]);
  assign t[73] = (~t[75] & t[86]);
  assign t[74] = (~t[75] & t[87]);
  assign t[75] = t[88] ^ x[4];
  assign t[76] = t[89] ^ x[5];
  assign t[77] = t[90] ^ x[9];
  assign t[78] = t[91] ^ x[10];
  assign t[79] = t[92] ^ x[12];
  assign t[7] = ~(t[52]);
  assign t[80] = t[93] ^ x[13];
  assign t[81] = t[94] ^ x[15];
  assign t[82] = t[95] ^ x[16];
  assign t[83] = t[96] ^ x[19];
  assign t[84] = t[97] ^ x[20];
  assign t[85] = t[98] ^ x[21];
  assign t[86] = t[99] ^ x[24];
  assign t[87] = t[100] ^ x[27];
  assign t[88] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[89] = (x[0]);
  assign t[8] = ~(t[12] & t[13]);
  assign t[90] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[8]);
  assign t[92] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[11]);
  assign t[94] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[95] = (x[14]);
  assign t[96] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[97] = (x[18]);
  assign t[98] = (x[1]);
  assign t[99] = (x[2]);
  assign t[9] = ~(t[14] & t[15]);
  assign y = (t[0] & ~t[44] & ~t[47] & ~t[49]) | (~t[0] & t[44] & ~t[47] & ~t[49]) | (~t[0] & ~t[44] & t[47] & ~t[49]) | (~t[0] & ~t[44] & ~t[47] & t[49]) | (t[0] & t[44] & t[47] & ~t[49]) | (t[0] & t[44] & ~t[47] & t[49]) | (t[0] & ~t[44] & t[47] & t[49]) | (~t[0] & t[44] & t[47] & t[49]);
endmodule

module R2ind291(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind292(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind293(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind294(x, y);
 input [20:0] x;
 output y;

 wire [78:0] t;
  assign t[0] = ~(t[44] ^ t[1]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = ~(t[16] | t[18]);
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = ~(t[23] & t[24]);
  assign t[15] = t[21] | t[25];
  assign t[16] = ~(t[21]);
  assign t[17] = t[46] ? t[27] : t[26];
  assign t[18] = t[46] ? t[29] : t[28];
  assign t[19] = ~(t[21] | t[30]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[16] | t[31]);
  assign t[21] = ~(t[45]);
  assign t[22] = ~(t[32] & t[33]);
  assign t[23] = t[47] & t[34];
  assign t[24] = t[35] | t[36];
  assign t[25] = t[46] ? t[32] : t[37];
  assign t[26] = ~(t[35] & t[38]);
  assign t[27] = ~(t[36] & t[47]);
  assign t[28] = ~(t[35] & t[47]);
  assign t[29] = ~(t[36] & t[38]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[46] ? t[26] : t[29];
  assign t[31] = t[46] ? t[37] : t[39];
  assign t[32] = ~(x[17] & t[40]);
  assign t[33] = ~(t[47] & t[41]);
  assign t[34] = ~(t[21] | t[46]);
  assign t[35] = ~(x[17] | t[48]);
  assign t[36] = x[17] & t[48];
  assign t[37] = ~(t[41] & t[38]);
  assign t[38] = ~(t[47]);
  assign t[39] = ~(x[17] & t[42]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = ~(t[48] | t[47]);
  assign t[41] = ~(x[17] | t[43]);
  assign t[42] = ~(t[48] | t[38]);
  assign t[43] = ~(t[48]);
  assign t[44] = (t[49]);
  assign t[45] = (t[50]);
  assign t[46] = (t[51]);
  assign t[47] = (t[52]);
  assign t[48] = (t[53]);
  assign t[49] = t[54] ^ x[5];
  assign t[4] = ~(t[7]);
  assign t[50] = t[55] ^ x[10];
  assign t[51] = t[56] ^ x[13];
  assign t[52] = t[57] ^ x[16];
  assign t[53] = t[58] ^ x[20];
  assign t[54] = (~t[59] & t[60]);
  assign t[55] = (~t[61] & t[62]);
  assign t[56] = (~t[63] & t[64]);
  assign t[57] = (~t[65] & t[66]);
  assign t[58] = (~t[67] & t[68]);
  assign t[59] = t[69] ^ x[4];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[5];
  assign t[61] = t[71] ^ x[9];
  assign t[62] = t[72] ^ x[10];
  assign t[63] = t[73] ^ x[12];
  assign t[64] = t[74] ^ x[13];
  assign t[65] = t[75] ^ x[15];
  assign t[66] = t[76] ^ x[16];
  assign t[67] = t[77] ^ x[19];
  assign t[68] = t[78] ^ x[20];
  assign t[69] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (x[0]);
  assign t[71] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[8]);
  assign t[73] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[11]);
  assign t[75] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[14]);
  assign t[77] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[18]);
  assign t[7] = ~(t[45]);
  assign t[8] = ~(t[12] & t[13]);
  assign t[9] = ~(t[14] & t[15]);
  assign y = (t[0]);
endmodule

module R2ind295(x, y);
 input [29:0] x;
 output y;

 wire [95:0] t;
  assign t[0] = ~(t[46] ^ t[1]);
  assign t[10] = ~(t[14] | t[16]);
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[47]);
  assign t[13] = t[48] ? t[20] : t[19];
  assign t[14] = ~(t[12]);
  assign t[15] = t[48] ? t[22] : t[21];
  assign t[16] = t[48] ? t[23] : t[19];
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = t[12] | t[26];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[29] & t[28]);
  assign t[21] = ~(x[14] & t[30]);
  assign t[22] = ~(t[31] & t[28]);
  assign t[23] = ~(t[29] & t[49]);
  assign t[24] = ~(t[14] | t[32]);
  assign t[25] = ~(t[14] | t[33]);
  assign t[26] = t[48] ? t[34] : t[22];
  assign t[27] = x[14] & t[50];
  assign t[28] = ~(t[49]);
  assign t[29] = ~(x[14] | t[50]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[50] | t[28]);
  assign t[31] = ~(x[14] | t[35]);
  assign t[32] = t[48] ? t[36] : t[20];
  assign t[33] = t[48] ? t[19] : t[23];
  assign t[34] = ~(x[14] & t[37]);
  assign t[35] = ~(t[50]);
  assign t[36] = ~(t[27] & t[49]);
  assign t[37] = ~(t[50] | t[49]);
  assign t[38] = t[39] ^ t[51];
  assign t[39] = t[4] ? x[23] : x[22];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[41] ^ t[52];
  assign t[41] = t[42] ? x[26] : x[25];
  assign t[42] = ~(t[7]);
  assign t[43] = t[44] ^ t[53];
  assign t[44] = t[45] ? x[29] : x[28];
  assign t[45] = ~(t[7]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = (t[57]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[58]);
  assign t[51] = (t[59]);
  assign t[52] = (t[60]);
  assign t[53] = (t[61]);
  assign t[54] = t[62] ^ x[5];
  assign t[55] = t[63] ^ x[10];
  assign t[56] = t[64] ^ x[13];
  assign t[57] = t[65] ^ x[17];
  assign t[58] = t[66] ^ x[20];
  assign t[59] = t[67] ^ x[21];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[68] ^ x[24];
  assign t[61] = t[69] ^ x[27];
  assign t[62] = (~t[70] & t[71]);
  assign t[63] = (~t[72] & t[73]);
  assign t[64] = (~t[74] & t[75]);
  assign t[65] = (~t[76] & t[77]);
  assign t[66] = (~t[78] & t[79]);
  assign t[67] = (~t[70] & t[80]);
  assign t[68] = (~t[70] & t[81]);
  assign t[69] = (~t[70] & t[82]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[83] ^ x[4];
  assign t[71] = t[84] ^ x[5];
  assign t[72] = t[85] ^ x[9];
  assign t[73] = t[86] ^ x[10];
  assign t[74] = t[87] ^ x[12];
  assign t[75] = t[88] ^ x[13];
  assign t[76] = t[89] ^ x[16];
  assign t[77] = t[90] ^ x[17];
  assign t[78] = t[91] ^ x[19];
  assign t[79] = t[92] ^ x[20];
  assign t[7] = ~(t[47]);
  assign t[80] = t[93] ^ x[21];
  assign t[81] = t[94] ^ x[24];
  assign t[82] = t[95] ^ x[27];
  assign t[83] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[84] = (x[0]);
  assign t[85] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[8]);
  assign t[87] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[11]);
  assign t[89] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[12] | t[13]);
  assign t[90] = (x[15]);
  assign t[91] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[18]);
  assign t[93] = (x[1]);
  assign t[94] = (x[2]);
  assign t[95] = (x[3]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = (t[0] & ~t[38] & ~t[40] & ~t[43]) | (~t[0] & t[38] & ~t[40] & ~t[43]) | (~t[0] & ~t[38] & t[40] & ~t[43]) | (~t[0] & ~t[38] & ~t[40] & t[43]) | (t[0] & t[38] & t[40] & ~t[43]) | (t[0] & t[38] & ~t[40] & t[43]) | (t[0] & ~t[38] & t[40] & t[43]) | (~t[0] & t[38] & t[40] & t[43]);
endmodule

module R2ind296(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind297(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind298(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind299(x, y);
 input [20:0] x;
 output y;

 wire [72:0] t;
  assign t[0] = ~(t[38] ^ t[1]);
  assign t[10] = ~(t[14] | t[16]);
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[39]);
  assign t[13] = t[40] ? t[20] : t[19];
  assign t[14] = ~(t[12]);
  assign t[15] = t[40] ? t[22] : t[21];
  assign t[16] = t[40] ? t[23] : t[19];
  assign t[17] = ~(t[24] | t[25]);
  assign t[18] = t[12] | t[26];
  assign t[19] = ~(t[27] & t[28]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[29] & t[28]);
  assign t[21] = ~(x[14] & t[30]);
  assign t[22] = ~(t[31] & t[28]);
  assign t[23] = ~(t[29] & t[41]);
  assign t[24] = ~(t[14] | t[32]);
  assign t[25] = ~(t[14] | t[33]);
  assign t[26] = t[40] ? t[34] : t[22];
  assign t[27] = x[14] & t[42];
  assign t[28] = ~(t[41]);
  assign t[29] = ~(x[14] | t[42]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[42] | t[28]);
  assign t[31] = ~(x[14] | t[35]);
  assign t[32] = t[40] ? t[36] : t[20];
  assign t[33] = t[40] ? t[19] : t[23];
  assign t[34] = ~(x[14] & t[37]);
  assign t[35] = ~(t[42]);
  assign t[36] = ~(t[27] & t[41]);
  assign t[37] = ~(t[42] | t[41]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = (t[47]);
  assign t[43] = t[48] ^ x[5];
  assign t[44] = t[49] ^ x[10];
  assign t[45] = t[50] ^ x[13];
  assign t[46] = t[51] ^ x[17];
  assign t[47] = t[52] ^ x[20];
  assign t[48] = (~t[53] & t[54]);
  assign t[49] = (~t[55] & t[56]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[57] & t[58]);
  assign t[51] = (~t[59] & t[60]);
  assign t[52] = (~t[61] & t[62]);
  assign t[53] = t[63] ^ x[4];
  assign t[54] = t[64] ^ x[5];
  assign t[55] = t[65] ^ x[9];
  assign t[56] = t[66] ^ x[10];
  assign t[57] = t[67] ^ x[12];
  assign t[58] = t[68] ^ x[13];
  assign t[59] = t[69] ^ x[16];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[17];
  assign t[61] = t[71] ^ x[19];
  assign t[62] = t[72] ^ x[20];
  assign t[63] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[64] = (x[0]);
  assign t[65] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[8]);
  assign t[67] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[11]);
  assign t[69] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (x[15]);
  assign t[71] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[18]);
  assign t[7] = ~(t[39]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[14] | t[15]);
  assign y = (t[0]);
endmodule

module R2ind300(x, y);
 input [29:0] x;
 output y;

 wire [93:0] t;
  assign t[0] = ~(t[44] ^ t[1]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[15]);
  assign t[13] = t[46] ? t[20] : t[19];
  assign t[14] = t[46] ? t[22] : t[21];
  assign t[15] = ~(t[45]);
  assign t[16] = t[46] ? t[20] : t[21];
  assign t[17] = ~(t[23] | t[24]);
  assign t[18] = ~(t[25] & t[26]);
  assign t[19] = ~(t[27] & t[47]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[28] & t[29]);
  assign t[21] = ~(t[27] & t[29]);
  assign t[22] = ~(t[28] & t[47]);
  assign t[23] = ~(t[15] | t[30]);
  assign t[24] = ~(t[15] | t[31]);
  assign t[25] = ~(t[48] | t[29]);
  assign t[26] = t[12] & t[46];
  assign t[27] = x[20] & t[48];
  assign t[28] = ~(x[20] | t[48]);
  assign t[29] = ~(t[47]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[46] ? t[21] : t[20];
  assign t[31] = t[46] ? t[33] : t[32];
  assign t[32] = ~(x[20] & t[34]);
  assign t[33] = ~(t[35] & t[29]);
  assign t[34] = ~(t[48] | t[47]);
  assign t[35] = ~(x[20] | t[36]);
  assign t[36] = ~(t[48]);
  assign t[37] = t[38] ^ t[49];
  assign t[38] = t[39] ? x[23] : x[22];
  assign t[39] = ~(t[7]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[41] ^ t[50];
  assign t[41] = t[45] ? x[26] : x[25];
  assign t[42] = t[43] ^ t[51];
  assign t[43] = t[4] ? x[29] : x[28];
  assign t[44] = (t[52]);
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = (t[57]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[58]);
  assign t[51] = (t[59]);
  assign t[52] = t[60] ^ x[5];
  assign t[53] = t[61] ^ x[10];
  assign t[54] = t[62] ^ x[13];
  assign t[55] = t[63] ^ x[16];
  assign t[56] = t[64] ^ x[19];
  assign t[57] = t[65] ^ x[21];
  assign t[58] = t[66] ^ x[24];
  assign t[59] = t[67] ^ x[27];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (~t[68] & t[69]);
  assign t[61] = (~t[70] & t[71]);
  assign t[62] = (~t[72] & t[73]);
  assign t[63] = (~t[74] & t[75]);
  assign t[64] = (~t[76] & t[77]);
  assign t[65] = (~t[68] & t[78]);
  assign t[66] = (~t[68] & t[79]);
  assign t[67] = (~t[68] & t[80]);
  assign t[68] = t[81] ^ x[4];
  assign t[69] = t[82] ^ x[5];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[83] ^ x[9];
  assign t[71] = t[84] ^ x[10];
  assign t[72] = t[85] ^ x[12];
  assign t[73] = t[86] ^ x[13];
  assign t[74] = t[87] ^ x[15];
  assign t[75] = t[88] ^ x[16];
  assign t[76] = t[89] ^ x[18];
  assign t[77] = t[90] ^ x[19];
  assign t[78] = t[91] ^ x[21];
  assign t[79] = t[92] ^ x[24];
  assign t[7] = ~(t[45]);
  assign t[80] = t[93] ^ x[27];
  assign t[81] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[82] = (x[0]);
  assign t[83] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[8]);
  assign t[85] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[11]);
  assign t[87] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[14]);
  assign t[89] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[12] | t[13]);
  assign t[90] = (x[17]);
  assign t[91] = (x[1]);
  assign t[92] = (x[2]);
  assign t[93] = (x[3]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0] & ~t[37] & ~t[40] & ~t[42]) | (~t[0] & t[37] & ~t[40] & ~t[42]) | (~t[0] & ~t[37] & t[40] & ~t[42]) | (~t[0] & ~t[37] & ~t[40] & t[42]) | (t[0] & t[37] & t[40] & ~t[42]) | (t[0] & t[37] & ~t[40] & t[42]) | (t[0] & ~t[37] & t[40] & t[42]) | (~t[0] & t[37] & t[40] & t[42]);
endmodule

module R2ind301(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind302(x, y);
 input [10:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = t[1] ^ t[2];
  assign t[10] = t[14] ^ x[7];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[13] = (x[2]);
  assign t[14] = (x[6] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[6] & 1'b0 & ~1'b0 & ~1'b0) | (~x[6] & ~1'b0 & 1'b0 & ~1'b0) | (~x[6] & ~1'b0 & ~1'b0 & 1'b0) | (x[6] & 1'b0 & 1'b0 & ~1'b0) | (x[6] & 1'b0 & ~1'b0 & 1'b0) | (x[6] & ~1'b0 & 1'b0 & 1'b0) | (~x[6] & 1'b0 & 1'b0 & 1'b0);
  assign t[15] = (x[6]);
  assign t[1] = t[3] ? x[10] : x[9];
  assign t[2] = (t[4]);
  assign t[3] = (t[5]);
  assign t[4] = t[6] ^ x[5];
  assign t[5] = t[7] ^ x[8];
  assign t[6] = (~t[8] & t[9]);
  assign t[7] = (~t[10] & t[11]);
  assign t[8] = t[12] ^ x[4];
  assign t[9] = t[13] ^ x[5];
  assign y = (t[0]);
endmodule

module R2ind303(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind304(x, y);
 input [20:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[37] ^ t[1]);
  assign t[10] = ~(t[15] | t[16]);
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[15]);
  assign t[13] = t[39] ? t[20] : t[19];
  assign t[14] = t[39] ? t[22] : t[21];
  assign t[15] = ~(t[38]);
  assign t[16] = t[39] ? t[20] : t[21];
  assign t[17] = ~(t[23] | t[24]);
  assign t[18] = ~(t[25] & t[26]);
  assign t[19] = ~(t[27] & t[40]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[28] & t[29]);
  assign t[21] = ~(t[27] & t[29]);
  assign t[22] = ~(t[28] & t[40]);
  assign t[23] = ~(t[15] | t[30]);
  assign t[24] = ~(t[15] | t[31]);
  assign t[25] = ~(t[41] | t[29]);
  assign t[26] = t[12] & t[39];
  assign t[27] = x[20] & t[41];
  assign t[28] = ~(x[20] | t[41]);
  assign t[29] = ~(t[40]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[39] ? t[21] : t[20];
  assign t[31] = t[39] ? t[33] : t[32];
  assign t[32] = ~(x[20] & t[34]);
  assign t[33] = ~(t[35] & t[29]);
  assign t[34] = ~(t[41] | t[40]);
  assign t[35] = ~(x[20] | t[36]);
  assign t[36] = ~(t[41]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[45]);
  assign t[41] = (t[46]);
  assign t[42] = t[47] ^ x[5];
  assign t[43] = t[48] ^ x[10];
  assign t[44] = t[49] ^ x[13];
  assign t[45] = t[50] ^ x[16];
  assign t[46] = t[51] ^ x[19];
  assign t[47] = (~t[52] & t[53]);
  assign t[48] = (~t[54] & t[55]);
  assign t[49] = (~t[56] & t[57]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[58] & t[59]);
  assign t[51] = (~t[60] & t[61]);
  assign t[52] = t[62] ^ x[4];
  assign t[53] = t[63] ^ x[5];
  assign t[54] = t[64] ^ x[9];
  assign t[55] = t[65] ^ x[10];
  assign t[56] = t[66] ^ x[12];
  assign t[57] = t[67] ^ x[13];
  assign t[58] = t[68] ^ x[15];
  assign t[59] = t[69] ^ x[16];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[18];
  assign t[61] = t[71] ^ x[19];
  assign t[62] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[63] = (x[0]);
  assign t[64] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[8]);
  assign t[66] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[11]);
  assign t[68] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[14]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[71] = (x[17]);
  assign t[7] = ~(t[38]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0]);
endmodule

module R2ind305(x, y);
 input [29:0] x;
 output y;

 wire [104:0] t;
  assign t[0] = ~(t[55] ^ t[1]);
  assign t[100] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[101] = (x[18]);
  assign t[102] = (x[1]);
  assign t[103] = (x[2]);
  assign t[104] = (x[3]);
  assign t[10] = t[15] | t[16];
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[19]);
  assign t[13] = t[57] ? t[21] : t[20];
  assign t[14] = t[57] ? t[23] : t[22];
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[12] | t[26]);
  assign t[17] = ~(t[27] | t[28]);
  assign t[18] = t[19] | t[29];
  assign t[19] = ~(t[56]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[30] & t[31]);
  assign t[21] = ~(t[32] & t[58]);
  assign t[22] = ~(t[58] & t[33]);
  assign t[23] = ~(x[17] & t[34]);
  assign t[24] = ~(t[35] | t[36]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[57] ? t[22] : t[23];
  assign t[27] = ~(t[39]);
  assign t[28] = ~(t[12] | t[40]);
  assign t[29] = t[57] ? t[23] : t[41];
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(x[17] | t[59]);
  assign t[31] = ~(t[58]);
  assign t[32] = x[17] & t[59];
  assign t[33] = ~(x[17] | t[42]);
  assign t[34] = ~(t[59] | t[58]);
  assign t[35] = ~(t[19] | t[43]);
  assign t[36] = ~(t[19] | t[44]);
  assign t[37] = ~(t[59] | t[31]);
  assign t[38] = t[12] & t[57];
  assign t[39] = ~(t[45] & t[46]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[57] ? t[47] : t[41];
  assign t[41] = ~(t[33] & t[31]);
  assign t[42] = ~(t[59]);
  assign t[43] = t[57] ? t[48] : t[20];
  assign t[44] = t[57] ? t[41] : t[23];
  assign t[45] = ~(t[19] | t[57]);
  assign t[46] = ~(t[22] & t[47]);
  assign t[47] = ~(x[17] & t[37]);
  assign t[48] = ~(t[32] & t[31]);
  assign t[49] = t[50] ^ t[60];
  assign t[4] = ~(t[7]);
  assign t[50] = t[4] ? x[23] : x[22];
  assign t[51] = t[52] ^ t[61];
  assign t[52] = t[4] ? x[26] : x[25];
  assign t[53] = t[54] ^ t[62];
  assign t[54] = t[4] ? x[29] : x[28];
  assign t[55] = (t[63]);
  assign t[56] = (t[64]);
  assign t[57] = (t[65]);
  assign t[58] = (t[66]);
  assign t[59] = (t[67]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (t[68]);
  assign t[61] = (t[69]);
  assign t[62] = (t[70]);
  assign t[63] = t[71] ^ x[5];
  assign t[64] = t[72] ^ x[10];
  assign t[65] = t[73] ^ x[13];
  assign t[66] = t[74] ^ x[16];
  assign t[67] = t[75] ^ x[20];
  assign t[68] = t[76] ^ x[21];
  assign t[69] = t[77] ^ x[24];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[78] ^ x[27];
  assign t[71] = (~t[79] & t[80]);
  assign t[72] = (~t[81] & t[82]);
  assign t[73] = (~t[83] & t[84]);
  assign t[74] = (~t[85] & t[86]);
  assign t[75] = (~t[87] & t[88]);
  assign t[76] = (~t[79] & t[89]);
  assign t[77] = (~t[79] & t[90]);
  assign t[78] = (~t[79] & t[91]);
  assign t[79] = t[92] ^ x[4];
  assign t[7] = ~(t[56]);
  assign t[80] = t[93] ^ x[5];
  assign t[81] = t[94] ^ x[9];
  assign t[82] = t[95] ^ x[10];
  assign t[83] = t[96] ^ x[12];
  assign t[84] = t[97] ^ x[13];
  assign t[85] = t[98] ^ x[15];
  assign t[86] = t[99] ^ x[16];
  assign t[87] = t[100] ^ x[19];
  assign t[88] = t[101] ^ x[20];
  assign t[89] = t[102] ^ x[21];
  assign t[8] = ~(t[12] | t[13]);
  assign t[90] = t[103] ^ x[24];
  assign t[91] = t[104] ^ x[27];
  assign t[92] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[93] = (x[0]);
  assign t[94] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[95] = (x[8]);
  assign t[96] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[97] = (x[11]);
  assign t[98] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[99] = (x[14]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0] & ~t[49] & ~t[51] & ~t[53]) | (~t[0] & t[49] & ~t[51] & ~t[53]) | (~t[0] & ~t[49] & t[51] & ~t[53]) | (~t[0] & ~t[49] & ~t[51] & t[53]) | (t[0] & t[49] & t[51] & ~t[53]) | (t[0] & t[49] & ~t[51] & t[53]) | (t[0] & ~t[49] & t[51] & t[53]) | (~t[0] & t[49] & t[51] & t[53]);
endmodule

module R2ind306(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind307(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind308(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind309(x, y);
 input [20:0] x;
 output y;

 wire [83:0] t;
  assign t[0] = ~(t[49] ^ t[1]);
  assign t[10] = t[15] | t[16];
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[19]);
  assign t[13] = t[51] ? t[21] : t[20];
  assign t[14] = t[51] ? t[23] : t[22];
  assign t[15] = ~(t[24] & t[25]);
  assign t[16] = ~(t[12] | t[26]);
  assign t[17] = ~(t[27] | t[28]);
  assign t[18] = t[19] | t[29];
  assign t[19] = ~(t[50]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[30] & t[31]);
  assign t[21] = ~(t[32] & t[52]);
  assign t[22] = ~(t[52] & t[33]);
  assign t[23] = ~(x[17] & t[34]);
  assign t[24] = ~(t[35] | t[36]);
  assign t[25] = ~(t[37] & t[38]);
  assign t[26] = t[51] ? t[22] : t[23];
  assign t[27] = ~(t[39]);
  assign t[28] = ~(t[12] | t[40]);
  assign t[29] = t[51] ? t[23] : t[41];
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(x[17] | t[53]);
  assign t[31] = ~(t[52]);
  assign t[32] = x[17] & t[53];
  assign t[33] = ~(x[17] | t[42]);
  assign t[34] = ~(t[53] | t[52]);
  assign t[35] = ~(t[19] | t[43]);
  assign t[36] = ~(t[19] | t[44]);
  assign t[37] = ~(t[53] | t[31]);
  assign t[38] = t[12] & t[51];
  assign t[39] = ~(t[45] & t[46]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[51] ? t[47] : t[41];
  assign t[41] = ~(t[33] & t[31]);
  assign t[42] = ~(t[53]);
  assign t[43] = t[51] ? t[48] : t[20];
  assign t[44] = t[51] ? t[41] : t[23];
  assign t[45] = ~(t[19] | t[51]);
  assign t[46] = ~(t[22] & t[47]);
  assign t[47] = ~(x[17] & t[37]);
  assign t[48] = ~(t[32] & t[31]);
  assign t[49] = (t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[55]);
  assign t[51] = (t[56]);
  assign t[52] = (t[57]);
  assign t[53] = (t[58]);
  assign t[54] = t[59] ^ x[5];
  assign t[55] = t[60] ^ x[10];
  assign t[56] = t[61] ^ x[13];
  assign t[57] = t[62] ^ x[16];
  assign t[58] = t[63] ^ x[20];
  assign t[59] = (~t[64] & t[65]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (~t[66] & t[67]);
  assign t[61] = (~t[68] & t[69]);
  assign t[62] = (~t[70] & t[71]);
  assign t[63] = (~t[72] & t[73]);
  assign t[64] = t[74] ^ x[4];
  assign t[65] = t[75] ^ x[5];
  assign t[66] = t[76] ^ x[9];
  assign t[67] = t[77] ^ x[10];
  assign t[68] = t[78] ^ x[12];
  assign t[69] = t[79] ^ x[13];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[80] ^ x[15];
  assign t[71] = t[81] ^ x[16];
  assign t[72] = t[82] ^ x[19];
  assign t[73] = t[83] ^ x[20];
  assign t[74] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[75] = (x[0]);
  assign t[76] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[8]);
  assign t[78] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[11]);
  assign t[7] = ~(t[50]);
  assign t[80] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[14]);
  assign t[82] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[18]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0]);
endmodule

module R2ind310(x, y);
 input [29:0] x;
 output y;

 wire [90:0] t;
  assign t[0] = ~(t[41] ^ t[1]);
  assign t[10] = ~(t[43] | t[16]);
  assign t[11] = t[12] & t[44];
  assign t[12] = ~(t[17]);
  assign t[13] = t[44] ? t[19] : t[18];
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[17] & t[22]);
  assign t[16] = ~(t[45]);
  assign t[17] = ~(t[42]);
  assign t[18] = ~(t[23] & t[16]);
  assign t[19] = ~(t[24] & t[45]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[17] | t[25]);
  assign t[21] = ~(t[12] | t[26]);
  assign t[22] = ~(t[27] & t[28]);
  assign t[23] = ~(x[20] | t[43]);
  assign t[24] = x[20] & t[43];
  assign t[25] = t[44] ? t[18] : t[29];
  assign t[26] = t[44] ? t[31] : t[30];
  assign t[27] = ~(x[20] & t[32]);
  assign t[28] = ~(t[45] & t[33]);
  assign t[29] = ~(t[24] & t[16]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(x[20] & t[10]);
  assign t[31] = ~(t[33] & t[16]);
  assign t[32] = ~(t[43] | t[45]);
  assign t[33] = ~(x[20] | t[34]);
  assign t[34] = ~(t[43]);
  assign t[35] = t[36] ^ t[46];
  assign t[36] = t[4] ? x[23] : x[22];
  assign t[37] = t[38] ^ t[47];
  assign t[38] = t[4] ? x[26] : x[25];
  assign t[39] = t[40] ^ t[48];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[4] ? x[29] : x[28];
  assign t[41] = (t[49]);
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = (t[52]);
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = t[57] ^ x[5];
  assign t[4] = ~(t[7]);
  assign t[50] = t[58] ^ x[10];
  assign t[51] = t[59] ^ x[13];
  assign t[52] = t[60] ^ x[16];
  assign t[53] = t[61] ^ x[19];
  assign t[54] = t[62] ^ x[21];
  assign t[55] = t[63] ^ x[24];
  assign t[56] = t[64] ^ x[27];
  assign t[57] = (~t[65] & t[66]);
  assign t[58] = (~t[67] & t[68]);
  assign t[59] = (~t[69] & t[70]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[73] & t[74]);
  assign t[62] = (~t[65] & t[75]);
  assign t[63] = (~t[65] & t[76]);
  assign t[64] = (~t[65] & t[77]);
  assign t[65] = t[78] ^ x[4];
  assign t[66] = t[79] ^ x[5];
  assign t[67] = t[80] ^ x[9];
  assign t[68] = t[81] ^ x[10];
  assign t[69] = t[82] ^ x[12];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[83] ^ x[13];
  assign t[71] = t[84] ^ x[15];
  assign t[72] = t[85] ^ x[16];
  assign t[73] = t[86] ^ x[18];
  assign t[74] = t[87] ^ x[19];
  assign t[75] = t[88] ^ x[21];
  assign t[76] = t[89] ^ x[24];
  assign t[77] = t[90] ^ x[27];
  assign t[78] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[79] = (x[0]);
  assign t[7] = ~(t[42]);
  assign t[80] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[8]);
  assign t[82] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[11]);
  assign t[84] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[14]);
  assign t[86] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[17]);
  assign t[88] = (x[1]);
  assign t[89] = (x[2]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[90] = (x[3]);
  assign t[9] = ~(t[14] & t[15]);
  assign y = (t[0] & ~t[35] & ~t[37] & ~t[39]) | (~t[0] & t[35] & ~t[37] & ~t[39]) | (~t[0] & ~t[35] & t[37] & ~t[39]) | (~t[0] & ~t[35] & ~t[37] & t[39]) | (t[0] & t[35] & t[37] & ~t[39]) | (t[0] & t[35] & ~t[37] & t[39]) | (t[0] & ~t[35] & t[37] & t[39]) | (~t[0] & t[35] & t[37] & t[39]);
endmodule

module R2ind311(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind312(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind313(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind314(x, y);
 input [20:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[35] ^ t[1]);
  assign t[10] = ~(t[37] | t[16]);
  assign t[11] = t[12] & t[38];
  assign t[12] = ~(t[17]);
  assign t[13] = t[38] ? t[19] : t[18];
  assign t[14] = ~(t[20] | t[21]);
  assign t[15] = ~(t[17] & t[22]);
  assign t[16] = ~(t[39]);
  assign t[17] = ~(t[36]);
  assign t[18] = ~(t[23] & t[16]);
  assign t[19] = ~(t[24] & t[39]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[17] | t[25]);
  assign t[21] = ~(t[12] | t[26]);
  assign t[22] = ~(t[27] & t[28]);
  assign t[23] = ~(x[20] | t[37]);
  assign t[24] = x[20] & t[37];
  assign t[25] = t[38] ? t[18] : t[29];
  assign t[26] = t[38] ? t[31] : t[30];
  assign t[27] = ~(x[20] & t[32]);
  assign t[28] = ~(t[39] & t[33]);
  assign t[29] = ~(t[24] & t[16]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(x[20] & t[10]);
  assign t[31] = ~(t[33] & t[16]);
  assign t[32] = ~(t[37] | t[39]);
  assign t[33] = ~(x[20] | t[34]);
  assign t[34] = ~(t[37]);
  assign t[35] = (t[40]);
  assign t[36] = (t[41]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[45] ^ x[5];
  assign t[41] = t[46] ^ x[10];
  assign t[42] = t[47] ^ x[13];
  assign t[43] = t[48] ^ x[16];
  assign t[44] = t[49] ^ x[19];
  assign t[45] = (~t[50] & t[51]);
  assign t[46] = (~t[52] & t[53]);
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[7]);
  assign t[50] = t[60] ^ x[4];
  assign t[51] = t[61] ^ x[5];
  assign t[52] = t[62] ^ x[9];
  assign t[53] = t[63] ^ x[10];
  assign t[54] = t[64] ^ x[12];
  assign t[55] = t[65] ^ x[13];
  assign t[56] = t[66] ^ x[15];
  assign t[57] = t[67] ^ x[16];
  assign t[58] = t[68] ^ x[18];
  assign t[59] = t[69] ^ x[19];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[61] = (x[0]);
  assign t[62] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[8]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[11]);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[14]);
  assign t[68] = (x[17] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[17] & 1'b0 & ~1'b0 & ~1'b0) | (~x[17] & ~1'b0 & 1'b0 & ~1'b0) | (~x[17] & ~1'b0 & ~1'b0 & 1'b0) | (x[17] & 1'b0 & 1'b0 & ~1'b0) | (x[17] & 1'b0 & ~1'b0 & 1'b0) | (x[17] & ~1'b0 & 1'b0 & 1'b0) | (~x[17] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[17]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[7] = ~(t[36]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[14] & t[15]);
  assign y = (t[0]);
endmodule

module R2ind315(x, y);
 input [29:0] x;
 output y;

 wire [90:0] t;
  assign t[0] = ~(t[41] ^ t[1]);
  assign t[10] = t[43] & t[16];
  assign t[11] = t[17] | t[18];
  assign t[12] = ~(t[16] & t[19]);
  assign t[13] = ~(t[20] & t[21]);
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = ~(t[22] | t[24]);
  assign t[16] = ~(t[25] | t[44]);
  assign t[17] = ~(x[17] | t[45]);
  assign t[18] = x[17] & t[45];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[45] | t[28]);
  assign t[21] = t[22] & t[44];
  assign t[22] = ~(t[25]);
  assign t[23] = t[44] ? t[26] : t[29];
  assign t[24] = t[44] ? t[31] : t[30];
  assign t[25] = ~(t[42]);
  assign t[26] = ~(t[43] & t[32]);
  assign t[27] = ~(x[17] & t[20]);
  assign t[28] = ~(t[43]);
  assign t[29] = ~(x[17] & t[33]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[18] & t[28]);
  assign t[31] = ~(t[17] & t[43]);
  assign t[32] = ~(x[17] | t[34]);
  assign t[33] = ~(t[45] | t[43]);
  assign t[34] = ~(t[45]);
  assign t[35] = t[36] ^ t[46];
  assign t[36] = t[4] ? x[23] : x[22];
  assign t[37] = t[38] ^ t[47];
  assign t[38] = t[4] ? x[26] : x[25];
  assign t[39] = t[40] ^ t[48];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[4] ? x[29] : x[28];
  assign t[41] = (t[49]);
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = (t[52]);
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = t[57] ^ x[5];
  assign t[4] = ~(t[7]);
  assign t[50] = t[58] ^ x[10];
  assign t[51] = t[59] ^ x[13];
  assign t[52] = t[60] ^ x[16];
  assign t[53] = t[61] ^ x[20];
  assign t[54] = t[62] ^ x[21];
  assign t[55] = t[63] ^ x[24];
  assign t[56] = t[64] ^ x[27];
  assign t[57] = (~t[65] & t[66]);
  assign t[58] = (~t[67] & t[68]);
  assign t[59] = (~t[69] & t[70]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[73] & t[74]);
  assign t[62] = (~t[65] & t[75]);
  assign t[63] = (~t[65] & t[76]);
  assign t[64] = (~t[65] & t[77]);
  assign t[65] = t[78] ^ x[4];
  assign t[66] = t[79] ^ x[5];
  assign t[67] = t[80] ^ x[9];
  assign t[68] = t[81] ^ x[10];
  assign t[69] = t[82] ^ x[12];
  assign t[6] = ~(t[10] & t[11]);
  assign t[70] = t[83] ^ x[13];
  assign t[71] = t[84] ^ x[15];
  assign t[72] = t[85] ^ x[16];
  assign t[73] = t[86] ^ x[19];
  assign t[74] = t[87] ^ x[20];
  assign t[75] = t[88] ^ x[21];
  assign t[76] = t[89] ^ x[24];
  assign t[77] = t[90] ^ x[27];
  assign t[78] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[79] = (x[0]);
  assign t[7] = ~(t[42]);
  assign t[80] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[8]);
  assign t[82] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[11]);
  assign t[84] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[14]);
  assign t[86] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[18]);
  assign t[88] = (x[1]);
  assign t[89] = (x[2]);
  assign t[8] = ~(t[12] & t[13]);
  assign t[90] = (x[3]);
  assign t[9] = t[14] | t[15];
  assign y = (t[0] & ~t[35] & ~t[37] & ~t[39]) | (~t[0] & t[35] & ~t[37] & ~t[39]) | (~t[0] & ~t[35] & t[37] & ~t[39]) | (~t[0] & ~t[35] & ~t[37] & t[39]) | (t[0] & t[35] & t[37] & ~t[39]) | (t[0] & t[35] & ~t[37] & t[39]) | (t[0] & ~t[35] & t[37] & t[39]) | (~t[0] & t[35] & t[37] & t[39]);
endmodule

module R2ind316(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind317(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind318(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind319(x, y);
 input [20:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[35] ^ t[1]);
  assign t[10] = t[37] & t[16];
  assign t[11] = t[17] | t[18];
  assign t[12] = ~(t[16] & t[19]);
  assign t[13] = ~(t[20] & t[21]);
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = ~(t[22] | t[24]);
  assign t[16] = ~(t[25] | t[38]);
  assign t[17] = ~(x[17] | t[39]);
  assign t[18] = x[17] & t[39];
  assign t[19] = ~(t[26] & t[27]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[39] | t[28]);
  assign t[21] = t[22] & t[38];
  assign t[22] = ~(t[25]);
  assign t[23] = t[38] ? t[26] : t[29];
  assign t[24] = t[38] ? t[31] : t[30];
  assign t[25] = ~(t[36]);
  assign t[26] = ~(t[37] & t[32]);
  assign t[27] = ~(x[17] & t[20]);
  assign t[28] = ~(t[37]);
  assign t[29] = ~(x[17] & t[33]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[18] & t[28]);
  assign t[31] = ~(t[17] & t[37]);
  assign t[32] = ~(x[17] | t[34]);
  assign t[33] = ~(t[39] | t[37]);
  assign t[34] = ~(t[39]);
  assign t[35] = (t[40]);
  assign t[36] = (t[41]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[45] ^ x[5];
  assign t[41] = t[46] ^ x[10];
  assign t[42] = t[47] ^ x[13];
  assign t[43] = t[48] ^ x[16];
  assign t[44] = t[49] ^ x[20];
  assign t[45] = (~t[50] & t[51]);
  assign t[46] = (~t[52] & t[53]);
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[7]);
  assign t[50] = t[60] ^ x[4];
  assign t[51] = t[61] ^ x[5];
  assign t[52] = t[62] ^ x[9];
  assign t[53] = t[63] ^ x[10];
  assign t[54] = t[64] ^ x[12];
  assign t[55] = t[65] ^ x[13];
  assign t[56] = t[66] ^ x[15];
  assign t[57] = t[67] ^ x[16];
  assign t[58] = t[68] ^ x[19];
  assign t[59] = t[69] ^ x[20];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[61] = (x[0]);
  assign t[62] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[8]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[11]);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[14]);
  assign t[68] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[18]);
  assign t[6] = ~(t[10] & t[11]);
  assign t[7] = ~(t[36]);
  assign t[8] = ~(t[12] & t[13]);
  assign t[9] = t[14] | t[15];
  assign y = (t[0]);
endmodule

module R2ind320(x, y);
 input [29:0] x;
 output y;

 wire [90:0] t;
  assign t[0] = ~(t[41] ^ t[1]);
  assign t[10] = ~(t[11] | t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = t[43] ? t[17] : t[16];
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = t[43] ? t[21] : t[20];
  assign t[15] = ~(t[42]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[17] = ~(t[24] & t[44]);
  assign t[18] = ~(t[11] | t[25]);
  assign t[19] = ~(t[11] | t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(x[17] & t[27]);
  assign t[21] = ~(t[44] & t[28]);
  assign t[22] = ~(x[17] | t[45]);
  assign t[23] = ~(t[44]);
  assign t[24] = x[17] & t[45];
  assign t[25] = t[43] ? t[30] : t[29];
  assign t[26] = t[43] ? t[32] : t[31];
  assign t[27] = ~(t[45] | t[44]);
  assign t[28] = ~(x[17] | t[33]);
  assign t[29] = ~(t[28] & t[23]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(x[17] & t[34]);
  assign t[31] = ~(t[22] & t[44]);
  assign t[32] = ~(t[24] & t[23]);
  assign t[33] = ~(t[45]);
  assign t[34] = ~(t[45] | t[23]);
  assign t[35] = t[36] ^ t[46];
  assign t[36] = t[4] ? x[23] : x[22];
  assign t[37] = t[38] ^ t[47];
  assign t[38] = t[4] ? x[26] : x[25];
  assign t[39] = t[40] ^ t[48];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[4] ? x[29] : x[28];
  assign t[41] = (t[49]);
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = (t[52]);
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = t[57] ^ x[5];
  assign t[4] = ~(t[7]);
  assign t[50] = t[58] ^ x[10];
  assign t[51] = t[59] ^ x[13];
  assign t[52] = t[60] ^ x[16];
  assign t[53] = t[61] ^ x[20];
  assign t[54] = t[62] ^ x[21];
  assign t[55] = t[63] ^ x[24];
  assign t[56] = t[64] ^ x[27];
  assign t[57] = (~t[65] & t[66]);
  assign t[58] = (~t[67] & t[68]);
  assign t[59] = (~t[69] & t[70]);
  assign t[5] = ~(t[8]);
  assign t[60] = (~t[71] & t[72]);
  assign t[61] = (~t[73] & t[74]);
  assign t[62] = (~t[65] & t[75]);
  assign t[63] = (~t[65] & t[76]);
  assign t[64] = (~t[65] & t[77]);
  assign t[65] = t[78] ^ x[4];
  assign t[66] = t[79] ^ x[5];
  assign t[67] = t[80] ^ x[9];
  assign t[68] = t[81] ^ x[10];
  assign t[69] = t[82] ^ x[12];
  assign t[6] = ~(t[9] | t[10]);
  assign t[70] = t[83] ^ x[13];
  assign t[71] = t[84] ^ x[15];
  assign t[72] = t[85] ^ x[16];
  assign t[73] = t[86] ^ x[19];
  assign t[74] = t[87] ^ x[20];
  assign t[75] = t[88] ^ x[21];
  assign t[76] = t[89] ^ x[24];
  assign t[77] = t[90] ^ x[27];
  assign t[78] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[79] = (x[0]);
  assign t[7] = ~(t[42]);
  assign t[80] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[81] = (x[8]);
  assign t[82] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[83] = (x[11]);
  assign t[84] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[85] = (x[14]);
  assign t[86] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[87] = (x[18]);
  assign t[88] = (x[1]);
  assign t[89] = (x[2]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[90] = (x[3]);
  assign t[9] = ~(t[13]);
  assign y = (t[0] & ~t[35] & ~t[37] & ~t[39]) | (~t[0] & t[35] & ~t[37] & ~t[39]) | (~t[0] & ~t[35] & t[37] & ~t[39]) | (~t[0] & ~t[35] & ~t[37] & t[39]) | (t[0] & t[35] & t[37] & ~t[39]) | (t[0] & t[35] & ~t[37] & t[39]) | (t[0] & ~t[35] & t[37] & t[39]) | (~t[0] & t[35] & t[37] & t[39]);
endmodule

module R2ind321(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind322(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind323(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind324(x, y);
 input [20:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[35] ^ t[1]);
  assign t[10] = ~(t[11] | t[14]);
  assign t[11] = ~(t[15]);
  assign t[12] = t[37] ? t[17] : t[16];
  assign t[13] = ~(t[18] | t[19]);
  assign t[14] = t[37] ? t[21] : t[20];
  assign t[15] = ~(t[36]);
  assign t[16] = ~(t[22] & t[23]);
  assign t[17] = ~(t[24] & t[38]);
  assign t[18] = ~(t[11] | t[25]);
  assign t[19] = ~(t[11] | t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(x[17] & t[27]);
  assign t[21] = ~(t[38] & t[28]);
  assign t[22] = ~(x[17] | t[39]);
  assign t[23] = ~(t[38]);
  assign t[24] = x[17] & t[39];
  assign t[25] = t[37] ? t[30] : t[29];
  assign t[26] = t[37] ? t[32] : t[31];
  assign t[27] = ~(t[39] | t[38]);
  assign t[28] = ~(x[17] | t[33]);
  assign t[29] = ~(t[28] & t[23]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(x[17] & t[34]);
  assign t[31] = ~(t[22] & t[38]);
  assign t[32] = ~(t[24] & t[23]);
  assign t[33] = ~(t[39]);
  assign t[34] = ~(t[39] | t[23]);
  assign t[35] = (t[40]);
  assign t[36] = (t[41]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[45] ^ x[5];
  assign t[41] = t[46] ^ x[10];
  assign t[42] = t[47] ^ x[13];
  assign t[43] = t[48] ^ x[16];
  assign t[44] = t[49] ^ x[20];
  assign t[45] = (~t[50] & t[51]);
  assign t[46] = (~t[52] & t[53]);
  assign t[47] = (~t[54] & t[55]);
  assign t[48] = (~t[56] & t[57]);
  assign t[49] = (~t[58] & t[59]);
  assign t[4] = ~(t[7]);
  assign t[50] = t[60] ^ x[4];
  assign t[51] = t[61] ^ x[5];
  assign t[52] = t[62] ^ x[9];
  assign t[53] = t[63] ^ x[10];
  assign t[54] = t[64] ^ x[12];
  assign t[55] = t[65] ^ x[13];
  assign t[56] = t[66] ^ x[15];
  assign t[57] = t[67] ^ x[16];
  assign t[58] = t[68] ^ x[19];
  assign t[59] = t[69] ^ x[20];
  assign t[5] = ~(t[8]);
  assign t[60] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[61] = (x[0]);
  assign t[62] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[63] = (x[8]);
  assign t[64] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[65] = (x[11]);
  assign t[66] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[67] = (x[14]);
  assign t[68] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[69] = (x[18]);
  assign t[6] = ~(t[9] | t[10]);
  assign t[7] = ~(t[36]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind325(x, y);
 input [29:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[36] ^ t[1]);
  assign t[10] = ~(t[16]);
  assign t[11] = t[38] ? t[18] : t[17];
  assign t[12] = ~(t[16] | t[19]);
  assign t[13] = ~(t[16] | t[20]);
  assign t[14] = ~(t[39] | t[21]);
  assign t[15] = t[10] & t[38];
  assign t[16] = ~(t[37]);
  assign t[17] = ~(x[17] & t[22]);
  assign t[18] = ~(t[40] & t[23]);
  assign t[19] = t[38] ? t[25] : t[24];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[38] ? t[26] : t[17];
  assign t[21] = ~(t[40]);
  assign t[22] = ~(t[39] | t[40]);
  assign t[23] = ~(x[17] | t[27]);
  assign t[24] = ~(t[28] & t[21]);
  assign t[25] = ~(t[29] & t[21]);
  assign t[26] = ~(t[23] & t[21]);
  assign t[27] = ~(t[39]);
  assign t[28] = ~(x[17] | t[39]);
  assign t[29] = x[17] & t[39];
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[31] ^ t[41];
  assign t[31] = t[4] ? x[23] : x[22];
  assign t[32] = t[33] ^ t[42];
  assign t[33] = t[4] ? x[26] : x[25];
  assign t[34] = t[35] ^ t[43];
  assign t[35] = t[4] ? x[29] : x[28];
  assign t[36] = (t[44]);
  assign t[37] = (t[45]);
  assign t[38] = (t[46]);
  assign t[39] = (t[47]);
  assign t[3] = t[5] | t[6];
  assign t[40] = (t[48]);
  assign t[41] = (t[49]);
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = t[52] ^ x[5];
  assign t[45] = t[53] ^ x[10];
  assign t[46] = t[54] ^ x[13];
  assign t[47] = t[55] ^ x[16];
  assign t[48] = t[56] ^ x[20];
  assign t[49] = t[57] ^ x[21];
  assign t[4] = ~(t[7]);
  assign t[50] = t[58] ^ x[24];
  assign t[51] = t[59] ^ x[27];
  assign t[52] = (~t[60] & t[61]);
  assign t[53] = (~t[62] & t[63]);
  assign t[54] = (~t[64] & t[65]);
  assign t[55] = (~t[66] & t[67]);
  assign t[56] = (~t[68] & t[69]);
  assign t[57] = (~t[60] & t[70]);
  assign t[58] = (~t[60] & t[71]);
  assign t[59] = (~t[60] & t[72]);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = t[73] ^ x[4];
  assign t[61] = t[74] ^ x[5];
  assign t[62] = t[75] ^ x[9];
  assign t[63] = t[76] ^ x[10];
  assign t[64] = t[77] ^ x[12];
  assign t[65] = t[78] ^ x[13];
  assign t[66] = t[79] ^ x[15];
  assign t[67] = t[80] ^ x[16];
  assign t[68] = t[81] ^ x[19];
  assign t[69] = t[82] ^ x[20];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[83] ^ x[21];
  assign t[71] = t[84] ^ x[24];
  assign t[72] = t[85] ^ x[27];
  assign t[73] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[74] = (x[0]);
  assign t[75] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[8]);
  assign t[77] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[78] = (x[11]);
  assign t[79] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[37]);
  assign t[80] = (x[14]);
  assign t[81] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[18]);
  assign t[83] = (x[1]);
  assign t[84] = (x[2]);
  assign t[85] = (x[3]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[14] & t[15]);
  assign y = (t[0] & ~t[30] & ~t[32] & ~t[34]) | (~t[0] & t[30] & ~t[32] & ~t[34]) | (~t[0] & ~t[30] & t[32] & ~t[34]) | (~t[0] & ~t[30] & ~t[32] & t[34]) | (t[0] & t[30] & t[32] & ~t[34]) | (t[0] & t[30] & ~t[32] & t[34]) | (t[0] & ~t[30] & t[32] & t[34]) | (~t[0] & t[30] & t[32] & t[34]);
endmodule

module R2ind326(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind327(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind328(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind329(x, y);
 input [20:0] x;
 output y;

 wire [64:0] t;
  assign t[0] = ~(t[30] ^ t[1]);
  assign t[10] = ~(t[16]);
  assign t[11] = t[32] ? t[18] : t[17];
  assign t[12] = ~(t[16] | t[19]);
  assign t[13] = ~(t[16] | t[20]);
  assign t[14] = ~(t[33] | t[21]);
  assign t[15] = t[10] & t[32];
  assign t[16] = ~(t[31]);
  assign t[17] = ~(x[17] & t[22]);
  assign t[18] = ~(t[34] & t[23]);
  assign t[19] = t[32] ? t[25] : t[24];
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = t[32] ? t[26] : t[17];
  assign t[21] = ~(t[34]);
  assign t[22] = ~(t[33] | t[34]);
  assign t[23] = ~(x[17] | t[27]);
  assign t[24] = ~(t[28] & t[21]);
  assign t[25] = ~(t[29] & t[21]);
  assign t[26] = ~(t[23] & t[21]);
  assign t[27] = ~(t[33]);
  assign t[28] = ~(x[17] | t[33]);
  assign t[29] = x[17] & t[33];
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = (t[35]);
  assign t[31] = (t[36]);
  assign t[32] = (t[37]);
  assign t[33] = (t[38]);
  assign t[34] = (t[39]);
  assign t[35] = t[40] ^ x[5];
  assign t[36] = t[41] ^ x[10];
  assign t[37] = t[42] ^ x[13];
  assign t[38] = t[43] ^ x[16];
  assign t[39] = t[44] ^ x[20];
  assign t[3] = t[5] | t[6];
  assign t[40] = (~t[45] & t[46]);
  assign t[41] = (~t[47] & t[48]);
  assign t[42] = (~t[49] & t[50]);
  assign t[43] = (~t[51] & t[52]);
  assign t[44] = (~t[53] & t[54]);
  assign t[45] = t[55] ^ x[4];
  assign t[46] = t[56] ^ x[5];
  assign t[47] = t[57] ^ x[9];
  assign t[48] = t[58] ^ x[10];
  assign t[49] = t[59] ^ x[12];
  assign t[4] = ~(t[7]);
  assign t[50] = t[60] ^ x[13];
  assign t[51] = t[61] ^ x[15];
  assign t[52] = t[62] ^ x[16];
  assign t[53] = t[63] ^ x[19];
  assign t[54] = t[64] ^ x[20];
  assign t[55] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[56] = (x[0]);
  assign t[57] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[58] = (x[8]);
  assign t[59] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[5] = ~(t[8] & t[9]);
  assign t[60] = (x[11]);
  assign t[61] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[14]);
  assign t[63] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[18]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[7] = ~(t[31]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[14] & t[15]);
  assign y = (t[0]);
endmodule

module R2ind330(x, y);
 input [29:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[51] ^ t[1]);
  assign t[100] = (x[3]);
  assign t[10] = ~(t[11] | t[15]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[53] ? t[18] : t[17];
  assign t[13] = ~(t[19] | t[20]);
  assign t[14] = ~(t[21] | t[22]);
  assign t[15] = t[53] ? t[24] : t[23];
  assign t[16] = ~(t[52]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(x[14] & t[27]);
  assign t[19] = ~(t[11] | t[28]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = ~(t[16] | t[31]);
  assign t[22] = ~(t[16] | t[32]);
  assign t[23] = ~(t[33] & t[54]);
  assign t[24] = ~(t[34] & t[26]);
  assign t[25] = ~(x[14] | t[35]);
  assign t[26] = ~(t[54]);
  assign t[27] = ~(t[55] | t[26]);
  assign t[28] = t[53] ? t[23] : t[24];
  assign t[29] = ~(t[36] | t[37]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[16] & t[38]);
  assign t[31] = t[53] ? t[39] : t[24];
  assign t[32] = t[53] ? t[17] : t[40];
  assign t[33] = x[14] & t[55];
  assign t[34] = ~(x[14] | t[55]);
  assign t[35] = ~(t[55]);
  assign t[36] = ~(t[16] | t[41]);
  assign t[37] = ~(t[11] | t[42]);
  assign t[38] = ~(t[40] & t[43]);
  assign t[39] = ~(t[33] & t[26]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = ~(x[14] & t[44]);
  assign t[41] = t[53] ? t[24] : t[39];
  assign t[42] = t[53] ? t[17] : t[18];
  assign t[43] = ~(t[54] & t[25]);
  assign t[44] = ~(t[55] | t[54]);
  assign t[45] = t[46] ^ t[56];
  assign t[46] = t[4] ? x[23] : x[22];
  assign t[47] = t[48] ^ t[57];
  assign t[48] = t[4] ? x[26] : x[25];
  assign t[49] = t[50] ^ t[58];
  assign t[4] = ~(t[7]);
  assign t[50] = t[4] ? x[29] : x[28];
  assign t[51] = (t[59]);
  assign t[52] = (t[60]);
  assign t[53] = (t[61]);
  assign t[54] = (t[62]);
  assign t[55] = (t[63]);
  assign t[56] = (t[64]);
  assign t[57] = (t[65]);
  assign t[58] = (t[66]);
  assign t[59] = t[67] ^ x[5];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[68] ^ x[10];
  assign t[61] = t[69] ^ x[13];
  assign t[62] = t[70] ^ x[17];
  assign t[63] = t[71] ^ x[20];
  assign t[64] = t[72] ^ x[21];
  assign t[65] = t[73] ^ x[24];
  assign t[66] = t[74] ^ x[27];
  assign t[67] = (~t[75] & t[76]);
  assign t[68] = (~t[77] & t[78]);
  assign t[69] = (~t[79] & t[80]);
  assign t[6] = ~(t[10]);
  assign t[70] = (~t[81] & t[82]);
  assign t[71] = (~t[83] & t[84]);
  assign t[72] = (~t[75] & t[85]);
  assign t[73] = (~t[75] & t[86]);
  assign t[74] = (~t[75] & t[87]);
  assign t[75] = t[88] ^ x[4];
  assign t[76] = t[89] ^ x[5];
  assign t[77] = t[90] ^ x[9];
  assign t[78] = t[91] ^ x[10];
  assign t[79] = t[92] ^ x[12];
  assign t[7] = ~(t[52]);
  assign t[80] = t[93] ^ x[13];
  assign t[81] = t[94] ^ x[16];
  assign t[82] = t[95] ^ x[17];
  assign t[83] = t[96] ^ x[19];
  assign t[84] = t[97] ^ x[20];
  assign t[85] = t[98] ^ x[21];
  assign t[86] = t[99] ^ x[24];
  assign t[87] = t[100] ^ x[27];
  assign t[88] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[89] = (x[0]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[90] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[91] = (x[8]);
  assign t[92] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[93] = (x[11]);
  assign t[94] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[95] = (x[15]);
  assign t[96] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[97] = (x[18]);
  assign t[98] = (x[1]);
  assign t[99] = (x[2]);
  assign t[9] = ~(t[13] & t[14]);
  assign y = (t[0] & ~t[45] & ~t[47] & ~t[49]) | (~t[0] & t[45] & ~t[47] & ~t[49]) | (~t[0] & ~t[45] & t[47] & ~t[49]) | (~t[0] & ~t[45] & ~t[47] & t[49]) | (t[0] & t[45] & t[47] & ~t[49]) | (t[0] & t[45] & ~t[47] & t[49]) | (t[0] & ~t[45] & t[47] & t[49]) | (~t[0] & t[45] & t[47] & t[49]);
endmodule

module R2ind331(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind332(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind333(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind334(x, y);
 input [20:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[45] ^ t[1]);
  assign t[10] = ~(t[11] | t[15]);
  assign t[11] = ~(t[16]);
  assign t[12] = t[47] ? t[18] : t[17];
  assign t[13] = ~(t[19] | t[20]);
  assign t[14] = ~(t[21] | t[22]);
  assign t[15] = t[47] ? t[24] : t[23];
  assign t[16] = ~(t[46]);
  assign t[17] = ~(t[25] & t[26]);
  assign t[18] = ~(x[14] & t[27]);
  assign t[19] = ~(t[11] | t[28]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[29] & t[30]);
  assign t[21] = ~(t[16] | t[31]);
  assign t[22] = ~(t[16] | t[32]);
  assign t[23] = ~(t[33] & t[48]);
  assign t[24] = ~(t[34] & t[26]);
  assign t[25] = ~(x[14] | t[35]);
  assign t[26] = ~(t[48]);
  assign t[27] = ~(t[49] | t[26]);
  assign t[28] = t[47] ? t[23] : t[24];
  assign t[29] = ~(t[36] | t[37]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[16] & t[38]);
  assign t[31] = t[47] ? t[39] : t[24];
  assign t[32] = t[47] ? t[17] : t[40];
  assign t[33] = x[14] & t[49];
  assign t[34] = ~(x[14] | t[49]);
  assign t[35] = ~(t[49]);
  assign t[36] = ~(t[16] | t[41]);
  assign t[37] = ~(t[11] | t[42]);
  assign t[38] = ~(t[40] & t[43]);
  assign t[39] = ~(t[33] & t[26]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = ~(x[14] & t[44]);
  assign t[41] = t[47] ? t[24] : t[39];
  assign t[42] = t[47] ? t[17] : t[18];
  assign t[43] = ~(t[48] & t[25]);
  assign t[44] = ~(t[49] | t[48]);
  assign t[45] = (t[50]);
  assign t[46] = (t[51]);
  assign t[47] = (t[52]);
  assign t[48] = (t[53]);
  assign t[49] = (t[54]);
  assign t[4] = ~(t[7]);
  assign t[50] = t[55] ^ x[5];
  assign t[51] = t[56] ^ x[10];
  assign t[52] = t[57] ^ x[13];
  assign t[53] = t[58] ^ x[17];
  assign t[54] = t[59] ^ x[20];
  assign t[55] = (~t[60] & t[61]);
  assign t[56] = (~t[62] & t[63]);
  assign t[57] = (~t[64] & t[65]);
  assign t[58] = (~t[66] & t[67]);
  assign t[59] = (~t[68] & t[69]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[4];
  assign t[61] = t[71] ^ x[5];
  assign t[62] = t[72] ^ x[9];
  assign t[63] = t[73] ^ x[10];
  assign t[64] = t[74] ^ x[12];
  assign t[65] = t[75] ^ x[13];
  assign t[66] = t[76] ^ x[16];
  assign t[67] = t[77] ^ x[17];
  assign t[68] = t[78] ^ x[19];
  assign t[69] = t[79] ^ x[20];
  assign t[6] = ~(t[10]);
  assign t[70] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[71] = (x[0]);
  assign t[72] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[73] = (x[8]);
  assign t[74] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[75] = (x[11]);
  assign t[76] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[77] = (x[15]);
  assign t[78] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[79] = (x[18]);
  assign t[7] = ~(t[46]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = ~(t[13] & t[14]);
  assign y = (t[0]);
endmodule

module R2ind335(x, y);
 input [29:0] x;
 output y;

 wire [89:0] t;
  assign t[0] = ~(t[40] ^ t[1]);
  assign t[10] = t[42] & t[15];
  assign t[11] = ~(t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[43] ? t[19] : t[18];
  assign t[14] = t[43] ? t[21] : t[20];
  assign t[15] = ~(t[17] | t[43]);
  assign t[16] = ~(t[22] | t[23]);
  assign t[17] = ~(t[41]);
  assign t[18] = ~(t[42] & t[24]);
  assign t[19] = ~(x[17] & t[25]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[26] & t[42]);
  assign t[21] = ~(t[27] & t[28]);
  assign t[22] = ~(t[17] | t[29]);
  assign t[23] = ~(t[17] | t[30]);
  assign t[24] = ~(x[17] | t[31]);
  assign t[25] = ~(t[44] | t[42]);
  assign t[26] = ~(x[17] | t[44]);
  assign t[27] = x[17] & t[44];
  assign t[28] = ~(t[42]);
  assign t[29] = t[43] ? t[21] : t[32];
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[43] ? t[33] : t[19];
  assign t[31] = ~(t[44]);
  assign t[32] = ~(t[26] & t[28]);
  assign t[33] = ~(t[24] & t[28]);
  assign t[34] = t[35] ^ t[45];
  assign t[35] = t[4] ? x[23] : x[22];
  assign t[36] = t[37] ^ t[46];
  assign t[37] = t[4] ? x[26] : x[25];
  assign t[38] = t[39] ^ t[47];
  assign t[39] = t[4] ? x[29] : x[28];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[48]);
  assign t[41] = (t[49]);
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = (t[52]);
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = t[56] ^ x[5];
  assign t[49] = t[57] ^ x[10];
  assign t[4] = ~(t[7]);
  assign t[50] = t[58] ^ x[13];
  assign t[51] = t[59] ^ x[16];
  assign t[52] = t[60] ^ x[20];
  assign t[53] = t[61] ^ x[21];
  assign t[54] = t[62] ^ x[24];
  assign t[55] = t[63] ^ x[27];
  assign t[56] = (~t[64] & t[65]);
  assign t[57] = (~t[66] & t[67]);
  assign t[58] = (~t[68] & t[69]);
  assign t[59] = (~t[70] & t[71]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (~t[72] & t[73]);
  assign t[61] = (~t[64] & t[74]);
  assign t[62] = (~t[64] & t[75]);
  assign t[63] = (~t[64] & t[76]);
  assign t[64] = t[77] ^ x[4];
  assign t[65] = t[78] ^ x[5];
  assign t[66] = t[79] ^ x[9];
  assign t[67] = t[80] ^ x[10];
  assign t[68] = t[81] ^ x[12];
  assign t[69] = t[82] ^ x[13];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[83] ^ x[15];
  assign t[71] = t[84] ^ x[16];
  assign t[72] = t[85] ^ x[19];
  assign t[73] = t[86] ^ x[20];
  assign t[74] = t[87] ^ x[21];
  assign t[75] = t[88] ^ x[24];
  assign t[76] = t[89] ^ x[27];
  assign t[77] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[78] = (x[0]);
  assign t[79] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[7] = ~(t[41]);
  assign t[80] = (x[8]);
  assign t[81] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[11]);
  assign t[83] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[14]);
  assign t[85] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[18]);
  assign t[87] = (x[1]);
  assign t[88] = (x[2]);
  assign t[89] = (x[3]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0] & ~t[34] & ~t[36] & ~t[38]) | (~t[0] & t[34] & ~t[36] & ~t[38]) | (~t[0] & ~t[34] & t[36] & ~t[38]) | (~t[0] & ~t[34] & ~t[36] & t[38]) | (t[0] & t[34] & t[36] & ~t[38]) | (t[0] & t[34] & ~t[36] & t[38]) | (t[0] & ~t[34] & t[36] & t[38]) | (~t[0] & t[34] & t[36] & t[38]);
endmodule

module R2ind336(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind337(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind338(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind339(x, y);
 input [20:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[34] ^ t[1]);
  assign t[10] = t[36] & t[15];
  assign t[11] = ~(t[16]);
  assign t[12] = ~(t[17]);
  assign t[13] = t[37] ? t[19] : t[18];
  assign t[14] = t[37] ? t[21] : t[20];
  assign t[15] = ~(t[17] | t[37]);
  assign t[16] = ~(t[22] | t[23]);
  assign t[17] = ~(t[35]);
  assign t[18] = ~(t[36] & t[24]);
  assign t[19] = ~(x[17] & t[25]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[26] & t[36]);
  assign t[21] = ~(t[27] & t[28]);
  assign t[22] = ~(t[17] | t[29]);
  assign t[23] = ~(t[17] | t[30]);
  assign t[24] = ~(x[17] | t[31]);
  assign t[25] = ~(t[38] | t[36]);
  assign t[26] = ~(x[17] | t[38]);
  assign t[27] = x[17] & t[38];
  assign t[28] = ~(t[36]);
  assign t[29] = t[37] ? t[21] : t[32];
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[37] ? t[33] : t[19];
  assign t[31] = ~(t[38]);
  assign t[32] = ~(t[26] & t[28]);
  assign t[33] = ~(t[24] & t[28]);
  assign t[34] = (t[39]);
  assign t[35] = (t[40]);
  assign t[36] = (t[41]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = t[44] ^ x[5];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[45] ^ x[10];
  assign t[41] = t[46] ^ x[13];
  assign t[42] = t[47] ^ x[16];
  assign t[43] = t[48] ^ x[20];
  assign t[44] = (~t[49] & t[50]);
  assign t[45] = (~t[51] & t[52]);
  assign t[46] = (~t[53] & t[54]);
  assign t[47] = (~t[55] & t[56]);
  assign t[48] = (~t[57] & t[58]);
  assign t[49] = t[59] ^ x[4];
  assign t[4] = ~(t[7]);
  assign t[50] = t[60] ^ x[5];
  assign t[51] = t[61] ^ x[9];
  assign t[52] = t[62] ^ x[10];
  assign t[53] = t[63] ^ x[12];
  assign t[54] = t[64] ^ x[13];
  assign t[55] = t[65] ^ x[15];
  assign t[56] = t[66] ^ x[16];
  assign t[57] = t[67] ^ x[19];
  assign t[58] = t[68] ^ x[20];
  assign t[59] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (x[0]);
  assign t[61] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[62] = (x[8]);
  assign t[63] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[11]);
  assign t[65] = (x[14] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[14] & 1'b0 & ~1'b0 & ~1'b0) | (~x[14] & ~1'b0 & 1'b0 & ~1'b0) | (~x[14] & ~1'b0 & ~1'b0 & 1'b0) | (x[14] & 1'b0 & 1'b0 & ~1'b0) | (x[14] & 1'b0 & ~1'b0 & 1'b0) | (x[14] & ~1'b0 & 1'b0 & 1'b0) | (~x[14] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[14]);
  assign t[67] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[18]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[7] = ~(t[35]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0]);
endmodule

module R2ind340(x, y);
 input [29:0] x;
 output y;

 wire [97:0] t;
  assign t[0] = ~(t[48] ^ t[1]);
  assign t[10] = ~(t[15] & t[16]);
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[49]);
  assign t[13] = t[50] ? t[20] : t[19];
  assign t[14] = t[50] ? t[22] : t[21];
  assign t[15] = ~(t[23] | t[24]);
  assign t[16] = ~(t[12] & t[25]);
  assign t[17] = ~(t[26] & t[27]);
  assign t[18] = t[12] | t[28];
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] & t[30]);
  assign t[21] = ~(x[14] & t[32]);
  assign t[22] = ~(t[33] & t[30]);
  assign t[23] = ~(t[12] | t[34]);
  assign t[24] = ~(t[35] | t[36]);
  assign t[25] = ~(t[21] & t[37]);
  assign t[26] = t[51] & t[38];
  assign t[27] = t[29] | t[31];
  assign t[28] = t[50] ? t[21] : t[22];
  assign t[29] = ~(x[14] | t[52]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[51]);
  assign t[31] = x[14] & t[52];
  assign t[32] = ~(t[52] | t[51]);
  assign t[33] = ~(x[14] | t[39]);
  assign t[34] = t[50] ? t[19] : t[20];
  assign t[35] = ~(t[12]);
  assign t[36] = t[50] ? t[22] : t[40];
  assign t[37] = ~(t[51] & t[33]);
  assign t[38] = ~(t[12] | t[50]);
  assign t[39] = ~(t[52]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = ~(x[14] & t[41]);
  assign t[41] = ~(t[52] | t[30]);
  assign t[42] = t[43] ^ t[53];
  assign t[43] = t[4] ? x[23] : x[22];
  assign t[44] = t[45] ^ t[54];
  assign t[45] = t[4] ? x[26] : x[25];
  assign t[46] = t[47] ^ t[55];
  assign t[47] = t[4] ? x[29] : x[28];
  assign t[48] = (t[56]);
  assign t[49] = (t[57]);
  assign t[4] = ~(t[7]);
  assign t[50] = (t[58]);
  assign t[51] = (t[59]);
  assign t[52] = (t[60]);
  assign t[53] = (t[61]);
  assign t[54] = (t[62]);
  assign t[55] = (t[63]);
  assign t[56] = t[64] ^ x[5];
  assign t[57] = t[65] ^ x[10];
  assign t[58] = t[66] ^ x[13];
  assign t[59] = t[67] ^ x[17];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[68] ^ x[20];
  assign t[61] = t[69] ^ x[21];
  assign t[62] = t[70] ^ x[24];
  assign t[63] = t[71] ^ x[27];
  assign t[64] = (~t[72] & t[73]);
  assign t[65] = (~t[74] & t[75]);
  assign t[66] = (~t[76] & t[77]);
  assign t[67] = (~t[78] & t[79]);
  assign t[68] = (~t[80] & t[81]);
  assign t[69] = (~t[72] & t[82]);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (~t[72] & t[83]);
  assign t[71] = (~t[72] & t[84]);
  assign t[72] = t[85] ^ x[4];
  assign t[73] = t[86] ^ x[5];
  assign t[74] = t[87] ^ x[9];
  assign t[75] = t[88] ^ x[10];
  assign t[76] = t[89] ^ x[12];
  assign t[77] = t[90] ^ x[13];
  assign t[78] = t[91] ^ x[16];
  assign t[79] = t[92] ^ x[17];
  assign t[7] = ~(t[49]);
  assign t[80] = t[93] ^ x[19];
  assign t[81] = t[94] ^ x[20];
  assign t[82] = t[95] ^ x[21];
  assign t[83] = t[96] ^ x[24];
  assign t[84] = t[97] ^ x[27];
  assign t[85] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[86] = (x[0]);
  assign t[87] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[8]);
  assign t[89] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[8] = ~(t[12] | t[13]);
  assign t[90] = (x[11]);
  assign t[91] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[92] = (x[15]);
  assign t[93] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[94] = (x[18]);
  assign t[95] = (x[1]);
  assign t[96] = (x[2]);
  assign t[97] = (x[3]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0] & ~t[42] & ~t[44] & ~t[46]) | (~t[0] & t[42] & ~t[44] & ~t[46]) | (~t[0] & ~t[42] & t[44] & ~t[46]) | (~t[0] & ~t[42] & ~t[44] & t[46]) | (t[0] & t[42] & t[44] & ~t[46]) | (t[0] & t[42] & ~t[44] & t[46]) | (t[0] & ~t[42] & t[44] & t[46]) | (~t[0] & t[42] & t[44] & t[46]);
endmodule

module R2ind341(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind342(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind343(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind344(x, y);
 input [20:0] x;
 output y;

 wire [76:0] t;
  assign t[0] = ~(t[42] ^ t[1]);
  assign t[10] = ~(t[15] & t[16]);
  assign t[11] = ~(t[17] & t[18]);
  assign t[12] = ~(t[43]);
  assign t[13] = t[44] ? t[20] : t[19];
  assign t[14] = t[44] ? t[22] : t[21];
  assign t[15] = ~(t[23] | t[24]);
  assign t[16] = ~(t[12] & t[25]);
  assign t[17] = ~(t[26] & t[27]);
  assign t[18] = t[12] | t[28];
  assign t[19] = ~(t[29] & t[30]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(t[31] & t[30]);
  assign t[21] = ~(x[14] & t[32]);
  assign t[22] = ~(t[33] & t[30]);
  assign t[23] = ~(t[12] | t[34]);
  assign t[24] = ~(t[35] | t[36]);
  assign t[25] = ~(t[21] & t[37]);
  assign t[26] = t[45] & t[38];
  assign t[27] = t[29] | t[31];
  assign t[28] = t[44] ? t[21] : t[22];
  assign t[29] = ~(x[14] | t[46]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = ~(t[45]);
  assign t[31] = x[14] & t[46];
  assign t[32] = ~(t[46] | t[45]);
  assign t[33] = ~(x[14] | t[39]);
  assign t[34] = t[44] ? t[19] : t[20];
  assign t[35] = ~(t[12]);
  assign t[36] = t[44] ? t[22] : t[40];
  assign t[37] = ~(t[45] & t[33]);
  assign t[38] = ~(t[12] | t[44]);
  assign t[39] = ~(t[46]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = ~(x[14] & t[41]);
  assign t[41] = ~(t[46] | t[30]);
  assign t[42] = (t[47]);
  assign t[43] = (t[48]);
  assign t[44] = (t[49]);
  assign t[45] = (t[50]);
  assign t[46] = (t[51]);
  assign t[47] = t[52] ^ x[5];
  assign t[48] = t[53] ^ x[10];
  assign t[49] = t[54] ^ x[13];
  assign t[4] = ~(t[7]);
  assign t[50] = t[55] ^ x[17];
  assign t[51] = t[56] ^ x[20];
  assign t[52] = (~t[57] & t[58]);
  assign t[53] = (~t[59] & t[60]);
  assign t[54] = (~t[61] & t[62]);
  assign t[55] = (~t[63] & t[64]);
  assign t[56] = (~t[65] & t[66]);
  assign t[57] = t[67] ^ x[4];
  assign t[58] = t[68] ^ x[5];
  assign t[59] = t[69] ^ x[9];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[10];
  assign t[61] = t[71] ^ x[12];
  assign t[62] = t[72] ^ x[13];
  assign t[63] = t[73] ^ x[16];
  assign t[64] = t[74] ^ x[17];
  assign t[65] = t[75] ^ x[19];
  assign t[66] = t[76] ^ x[20];
  assign t[67] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[68] = (x[0]);
  assign t[69] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (x[8]);
  assign t[71] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[72] = (x[11]);
  assign t[73] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[74] = (x[15]);
  assign t[75] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[76] = (x[18]);
  assign t[7] = ~(t[43]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0]);
endmodule

module R2ind345(x, y);
 input [29:0] x;
 output y;

 wire [91:0] t;
  assign t[0] = ~(t[42] ^ t[1]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[16] | t[17]);
  assign t[12] = ~(t[43]);
  assign t[13] = t[44] ? t[19] : t[18];
  assign t[14] = t[44] ? t[21] : t[20];
  assign t[15] = ~(t[22] | t[23]);
  assign t[16] = ~(t[12]);
  assign t[17] = t[44] ? t[24] : t[20];
  assign t[18] = ~(t[25] & t[26]);
  assign t[19] = ~(t[27] & t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(x[14] & t[28]);
  assign t[21] = ~(t[29] & t[26]);
  assign t[22] = ~(t[16] | t[30]);
  assign t[23] = ~(t[16] | t[31]);
  assign t[24] = ~(t[45] & t[29]);
  assign t[25] = x[14] & t[46];
  assign t[26] = ~(t[45]);
  assign t[27] = ~(x[14] | t[46]);
  assign t[28] = ~(t[46] | t[45]);
  assign t[29] = ~(x[14] | t[32]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[44] ? t[33] : t[21];
  assign t[31] = t[44] ? t[18] : t[34];
  assign t[32] = ~(t[46]);
  assign t[33] = ~(x[14] & t[35]);
  assign t[34] = ~(t[27] & t[45]);
  assign t[35] = ~(t[46] | t[26]);
  assign t[36] = t[37] ^ t[47];
  assign t[37] = t[4] ? x[23] : x[22];
  assign t[38] = t[39] ^ t[48];
  assign t[39] = t[4] ? x[26] : x[25];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[41] ^ t[49];
  assign t[41] = t[4] ? x[29] : x[28];
  assign t[42] = (t[50]);
  assign t[43] = (t[51]);
  assign t[44] = (t[52]);
  assign t[45] = (t[53]);
  assign t[46] = (t[54]);
  assign t[47] = (t[55]);
  assign t[48] = (t[56]);
  assign t[49] = (t[57]);
  assign t[4] = ~(t[7]);
  assign t[50] = t[58] ^ x[5];
  assign t[51] = t[59] ^ x[10];
  assign t[52] = t[60] ^ x[13];
  assign t[53] = t[61] ^ x[17];
  assign t[54] = t[62] ^ x[20];
  assign t[55] = t[63] ^ x[21];
  assign t[56] = t[64] ^ x[24];
  assign t[57] = t[65] ^ x[27];
  assign t[58] = (~t[66] & t[67]);
  assign t[59] = (~t[68] & t[69]);
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = (~t[70] & t[71]);
  assign t[61] = (~t[72] & t[73]);
  assign t[62] = (~t[74] & t[75]);
  assign t[63] = (~t[66] & t[76]);
  assign t[64] = (~t[66] & t[77]);
  assign t[65] = (~t[66] & t[78]);
  assign t[66] = t[79] ^ x[4];
  assign t[67] = t[80] ^ x[5];
  assign t[68] = t[81] ^ x[9];
  assign t[69] = t[82] ^ x[10];
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = t[83] ^ x[12];
  assign t[71] = t[84] ^ x[13];
  assign t[72] = t[85] ^ x[16];
  assign t[73] = t[86] ^ x[17];
  assign t[74] = t[87] ^ x[19];
  assign t[75] = t[88] ^ x[20];
  assign t[76] = t[89] ^ x[21];
  assign t[77] = t[90] ^ x[24];
  assign t[78] = t[91] ^ x[27];
  assign t[79] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[7] = ~(t[43]);
  assign t[80] = (x[0]);
  assign t[81] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[82] = (x[8]);
  assign t[83] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[84] = (x[11]);
  assign t[85] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[86] = (x[15]);
  assign t[87] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[88] = (x[18]);
  assign t[89] = (x[1]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[90] = (x[2]);
  assign t[91] = (x[3]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0] & ~t[36] & ~t[38] & ~t[40]) | (~t[0] & t[36] & ~t[38] & ~t[40]) | (~t[0] & ~t[36] & t[38] & ~t[40]) | (~t[0] & ~t[36] & ~t[38] & t[40]) | (t[0] & t[36] & t[38] & ~t[40]) | (t[0] & t[36] & ~t[38] & t[40]) | (t[0] & ~t[36] & t[38] & t[40]) | (~t[0] & t[36] & t[38] & t[40]);
endmodule

module R2ind346(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[3]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind347(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[2]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind348(x, y);
 input [10:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[1] ^ t[4];
  assign t[10] = t[14] ^ x[4];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[9];
  assign t[13] = t[17] ^ x[10];
  assign t[14] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[15] = (x[1]);
  assign t[16] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[17] = (x[8]);
  assign t[1] = t[2] ? x[7] : x[6];
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[5]);
  assign t[4] = (t[6]);
  assign t[5] = (t[7]);
  assign t[6] = t[8] ^ x[5];
  assign t[7] = t[9] ^ x[10];
  assign t[8] = (~t[10] & t[11]);
  assign t[9] = (~t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind349(x, y);
 input [20:0] x;
 output y;

 wire [70:0] t;
  assign t[0] = ~(t[36] ^ t[1]);
  assign t[10] = ~(t[15]);
  assign t[11] = ~(t[16] | t[17]);
  assign t[12] = ~(t[37]);
  assign t[13] = t[38] ? t[19] : t[18];
  assign t[14] = t[38] ? t[21] : t[20];
  assign t[15] = ~(t[22] | t[23]);
  assign t[16] = ~(t[12]);
  assign t[17] = t[38] ? t[24] : t[20];
  assign t[18] = ~(t[25] & t[26]);
  assign t[19] = ~(t[27] & t[26]);
  assign t[1] = ~(t[2] ^ t[3]);
  assign t[20] = ~(x[14] & t[28]);
  assign t[21] = ~(t[29] & t[26]);
  assign t[22] = ~(t[16] | t[30]);
  assign t[23] = ~(t[16] | t[31]);
  assign t[24] = ~(t[39] & t[29]);
  assign t[25] = x[14] & t[40];
  assign t[26] = ~(t[39]);
  assign t[27] = ~(x[14] | t[40]);
  assign t[28] = ~(t[40] | t[39]);
  assign t[29] = ~(x[14] | t[32]);
  assign t[2] = t[4] ? x[7] : x[6];
  assign t[30] = t[38] ? t[33] : t[21];
  assign t[31] = t[38] ? t[18] : t[34];
  assign t[32] = ~(t[40]);
  assign t[33] = ~(x[14] & t[35]);
  assign t[34] = ~(t[27] & t[39]);
  assign t[35] = ~(t[40] | t[26]);
  assign t[36] = (t[41]);
  assign t[37] = (t[42]);
  assign t[38] = (t[43]);
  assign t[39] = (t[44]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = (t[45]);
  assign t[41] = t[46] ^ x[5];
  assign t[42] = t[47] ^ x[10];
  assign t[43] = t[48] ^ x[13];
  assign t[44] = t[49] ^ x[17];
  assign t[45] = t[50] ^ x[20];
  assign t[46] = (~t[51] & t[52]);
  assign t[47] = (~t[53] & t[54]);
  assign t[48] = (~t[55] & t[56]);
  assign t[49] = (~t[57] & t[58]);
  assign t[4] = ~(t[7]);
  assign t[50] = (~t[59] & t[60]);
  assign t[51] = t[61] ^ x[4];
  assign t[52] = t[62] ^ x[5];
  assign t[53] = t[63] ^ x[9];
  assign t[54] = t[64] ^ x[10];
  assign t[55] = t[65] ^ x[12];
  assign t[56] = t[66] ^ x[13];
  assign t[57] = t[67] ^ x[16];
  assign t[58] = t[68] ^ x[17];
  assign t[59] = t[69] ^ x[19];
  assign t[5] = ~(t[8] | t[9]);
  assign t[60] = t[70] ^ x[20];
  assign t[61] = (x[0] & ~x[1] & ~x[2] & ~x[3]) | (~x[0] & x[1] & ~x[2] & ~x[3]) | (~x[0] & ~x[1] & x[2] & ~x[3]) | (~x[0] & ~x[1] & ~x[2] & x[3]) | (x[0] & x[1] & x[2] & ~x[3]) | (x[0] & x[1] & ~x[2] & x[3]) | (x[0] & ~x[1] & x[2] & x[3]) | (~x[0] & x[1] & x[2] & x[3]);
  assign t[62] = (x[0]);
  assign t[63] = (x[8] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[8] & 1'b0 & ~1'b0 & ~1'b0) | (~x[8] & ~1'b0 & 1'b0 & ~1'b0) | (~x[8] & ~1'b0 & ~1'b0 & 1'b0) | (x[8] & 1'b0 & 1'b0 & ~1'b0) | (x[8] & 1'b0 & ~1'b0 & 1'b0) | (x[8] & ~1'b0 & 1'b0 & 1'b0) | (~x[8] & 1'b0 & 1'b0 & 1'b0);
  assign t[64] = (x[8]);
  assign t[65] = (x[11] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[11] & 1'b0 & ~1'b0 & ~1'b0) | (~x[11] & ~1'b0 & 1'b0 & ~1'b0) | (~x[11] & ~1'b0 & ~1'b0 & 1'b0) | (x[11] & 1'b0 & 1'b0 & ~1'b0) | (x[11] & 1'b0 & ~1'b0 & 1'b0) | (x[11] & ~1'b0 & 1'b0 & 1'b0) | (~x[11] & 1'b0 & 1'b0 & 1'b0);
  assign t[66] = (x[11]);
  assign t[67] = (x[15] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[15] & 1'b0 & ~1'b0 & ~1'b0) | (~x[15] & ~1'b0 & 1'b0 & ~1'b0) | (~x[15] & ~1'b0 & ~1'b0 & 1'b0) | (x[15] & 1'b0 & 1'b0 & ~1'b0) | (x[15] & 1'b0 & ~1'b0 & 1'b0) | (x[15] & ~1'b0 & 1'b0 & 1'b0) | (~x[15] & 1'b0 & 1'b0 & 1'b0);
  assign t[68] = (x[15]);
  assign t[69] = (x[18] & ~1'b0 & ~1'b0 & ~1'b0) | (~x[18] & 1'b0 & ~1'b0 & ~1'b0) | (~x[18] & ~1'b0 & 1'b0 & ~1'b0) | (~x[18] & ~1'b0 & ~1'b0 & 1'b0) | (x[18] & 1'b0 & 1'b0 & ~1'b0) | (x[18] & 1'b0 & ~1'b0 & 1'b0) | (x[18] & ~1'b0 & 1'b0 & 1'b0) | (~x[18] & 1'b0 & 1'b0 & 1'b0);
  assign t[6] = ~(t[10] | t[11]);
  assign t[70] = (x[18]);
  assign t[7] = ~(t[37]);
  assign t[8] = ~(t[12] | t[13]);
  assign t[9] = ~(t[12] | t[14]);
  assign y = (t[0]);
endmodule

module R2ind350(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind351(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind352(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind353(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind354(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind355(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind356(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind357(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind358(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind359(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind360(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind361(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind362(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind363(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind364(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind365(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind366(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind367(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind368(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind369(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind370(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind371(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind372(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind373(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind374(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind375(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind376(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind377(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind378(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind379(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind380(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind381(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind382(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind383(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind384(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind385(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind386(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind387(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind388(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind389(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind390(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind391(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind392(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind393(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind394(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind395(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind396(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind397(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind398(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind399(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind400(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind401(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind402(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind403(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind404(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind405(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind406(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind407(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind408(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind409(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind410(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind411(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind412(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind413(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind414(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind415(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind416(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind417(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind418(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind419(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind420(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind421(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind422(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind423(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind424(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind425(x, y);
 input [18:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = x[0] ? t[5] : t[4];
  assign t[10] = (t[18]);
  assign t[11] = (t[19]);
  assign t[12] = t[20] ^ x[6];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[13];
  assign t[15] = t[23] ^ x[14];
  assign t[16] = t[24] ^ x[15];
  assign t[17] = t[25] ^ x[16];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[18];
  assign t[1] = x[0] ? t[7] : t[6];
  assign t[20] = (~t[28] & t[29]);
  assign t[21] = (~t[30] & t[31]);
  assign t[22] = (~t[28] & t[32]);
  assign t[23] = (~t[30] & t[33]);
  assign t[24] = (~t[28] & t[34]);
  assign t[25] = (~t[30] & t[35]);
  assign t[26] = (~t[28] & t[36]);
  assign t[27] = (~t[30] & t[37]);
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[6];
  assign t[2] = x[0] ? t[9] : t[8];
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[12];
  assign t[32] = t[42] ^ x[13];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[15];
  assign t[35] = t[45] ^ x[16];
  assign t[36] = t[46] ^ x[17];
  assign t[37] = t[47] ^ x[18];
  assign t[38] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[39] = (x[1]);
  assign t[3] = x[0] ? t[11] : t[10];
  assign t[40] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[41] = (x[7]);
  assign t[42] = (x[2]);
  assign t[43] = (x[8]);
  assign t[44] = (x[3]);
  assign t[45] = (x[9]);
  assign t[46] = (x[4]);
  assign t[47] = (x[10]);
  assign t[4] = (t[12]);
  assign t[5] = (t[13]);
  assign t[6] = (t[14]);
  assign t[7] = (t[15]);
  assign t[8] = (t[16]);
  assign t[9] = (t[17]);
  assign y = (t[0] & ~t[1] & ~t[2] & ~t[3]) | (~t[0] & t[1] & ~t[2] & ~t[3]) | (~t[0] & ~t[1] & t[2] & ~t[3]) | (~t[0] & ~t[1] & ~t[2] & t[3]) | (t[0] & t[1] & t[2] & ~t[3]) | (t[0] & t[1] & ~t[2] & t[3]) | (t[0] & ~t[1] & t[2] & t[3]) | (~t[0] & t[1] & t[2] & t[3]);
endmodule

module R2ind426(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[4]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[10]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind427(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[3]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[9]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind428(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[2]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[8]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2ind429(x, y);
 input [12:0] x;
 output y;

 wire [14:0] t;
  assign t[0] = x[0] ? t[2] : t[1];
  assign t[10] = t[14] ^ x[12];
  assign t[11] = (x[1] & ~x[2] & ~x[3] & ~x[4]) | (~x[1] & x[2] & ~x[3] & ~x[4]) | (~x[1] & ~x[2] & x[3] & ~x[4]) | (~x[1] & ~x[2] & ~x[3] & x[4]) | (x[1] & x[2] & x[3] & ~x[4]) | (x[1] & x[2] & ~x[3] & x[4]) | (x[1] & ~x[2] & x[3] & x[4]) | (~x[1] & x[2] & x[3] & x[4]);
  assign t[12] = (x[1]);
  assign t[13] = (x[7] & ~x[8] & ~x[9] & ~x[10]) | (~x[7] & x[8] & ~x[9] & ~x[10]) | (~x[7] & ~x[8] & x[9] & ~x[10]) | (~x[7] & ~x[8] & ~x[9] & x[10]) | (x[7] & x[8] & x[9] & ~x[10]) | (x[7] & x[8] & ~x[9] & x[10]) | (x[7] & ~x[8] & x[9] & x[10]) | (~x[7] & x[8] & x[9] & x[10]);
  assign t[14] = (x[7]);
  assign t[1] = (t[3]);
  assign t[2] = (t[4]);
  assign t[3] = t[5] ^ x[6];
  assign t[4] = t[6] ^ x[12];
  assign t[5] = (~t[7] & t[8]);
  assign t[6] = (~t[9] & t[10]);
  assign t[7] = t[11] ^ x[5];
  assign t[8] = t[12] ^ x[6];
  assign t[9] = t[13] ^ x[11];
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [787:0] x;
 output [429:0] y;

  R2ind0 R2ind0_inst(.x({x[5], x[4], x[3], x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[5], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[2], x[5], x[0]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[3], x[5], x[0]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[4], x[5], x[0]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[5]));
  R2ind6 R2ind6_inst(.y(y[6]));
  R2ind7 R2ind7_inst(.y(y[7]));
  R2ind8 R2ind8_inst(.y(y[8]));
  R2ind9 R2ind9_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[11], x[10], x[9], x[18]}), .y(y[10]));
  R2ind11 R2ind11_inst(.y(y[11]));
  R2ind12 R2ind12_inst(.y(y[12]));
  R2ind13 R2ind13_inst(.y(y[13]));
  R2ind14 R2ind14_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[11], x[10], x[9], x[18]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[11], x[10], x[9], x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[18]}), .y(y[15]));
  R2ind16 R2ind16_inst(.y(y[16]));
  R2ind17 R2ind17_inst(.y(y[17]));
  R2ind18 R2ind18_inst(.y(y[18]));
  R2ind19 R2ind19_inst(.x({x[11], x[10], x[9], x[14], x[13], x[12], x[17], x[16], x[15], x[8], x[7], x[6], x[18]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[18]}), .y(y[20]));
  R2ind21 R2ind21_inst(.y(y[21]));
  R2ind22 R2ind22_inst(.y(y[22]));
  R2ind23 R2ind23_inst(.y(y[23]));
  R2ind24 R2ind24_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[18]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[18]}), .y(y[25]));
  R2ind26 R2ind26_inst(.y(y[26]));
  R2ind27 R2ind27_inst(.y(y[27]));
  R2ind28 R2ind28_inst(.y(y[28]));
  R2ind29 R2ind29_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[18]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[35], x[34], x[33], x[32], x[31], x[30], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[35], x[34], x[33], x[23], x[22], x[21], x[20], x[19]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[32], x[31], x[30], x[23], x[22], x[21], x[20], x[19]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[29], x[28], x[27], x[23], x[22], x[21], x[20], x[19]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[52], x[51], x[50], x[49], x[48], x[47], x[46], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[52], x[51], x[50], x[40], x[39], x[38], x[37], x[36]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[49], x[48], x[47], x[40], x[39], x[38], x[37], x[36]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[46], x[45], x[44], x[40], x[39], x[38], x[37], x[36]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[69], x[68], x[67], x[66], x[65], x[64], x[63], x[62], x[61], x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[69], x[68], x[67], x[57], x[56], x[55], x[54], x[53]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[66], x[65], x[64], x[57], x[56], x[55], x[54], x[53]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[63], x[62], x[61], x[57], x[56], x[55], x[54], x[53]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[60], x[59], x[58], x[57], x[56], x[55], x[54], x[53]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[86], x[85], x[84], x[83], x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[86], x[85], x[84], x[74], x[73], x[72], x[71], x[70]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[83], x[82], x[81], x[74], x[73], x[72], x[71], x[70]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[80], x[79], x[78], x[74], x[73], x[72], x[71], x[70]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[103], x[102], x[101], x[100], x[99], x[98], x[97], x[96], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[103], x[102], x[101], x[91], x[90], x[89], x[88], x[87]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[100], x[99], x[98], x[91], x[90], x[89], x[88], x[87]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[97], x[96], x[95], x[91], x[90], x[89], x[88], x[87]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[120], x[119], x[118], x[108], x[107], x[106], x[105], x[104]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[117], x[116], x[115], x[108], x[107], x[106], x[105], x[104]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[114], x[113], x[112], x[108], x[107], x[106], x[105], x[104]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[111], x[110], x[109], x[108], x[107], x[106], x[105], x[104]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[137], x[136], x[135], x[134], x[133], x[132], x[131], x[130], x[129], x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[137], x[136], x[135], x[125], x[124], x[123], x[122], x[121]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[134], x[133], x[132], x[125], x[124], x[123], x[122], x[121]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[131], x[130], x[129], x[125], x[124], x[123], x[122], x[121]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[128], x[127], x[126], x[125], x[124], x[123], x[122], x[121]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[154], x[153], x[152], x[151], x[150], x[149], x[148], x[147], x[146], x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[154], x[153], x[152], x[142], x[141], x[140], x[139], x[138]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[151], x[150], x[149], x[142], x[141], x[140], x[139], x[138]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[148], x[147], x[146], x[142], x[141], x[140], x[139], x[138]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[145], x[144], x[143], x[142], x[141], x[140], x[139], x[138]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[171], x[170], x[169], x[168], x[167], x[166], x[165], x[164], x[163], x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[171], x[170], x[169], x[159], x[158], x[157], x[156], x[155]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[168], x[167], x[166], x[159], x[158], x[157], x[156], x[155]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[165], x[164], x[163], x[159], x[158], x[157], x[156], x[155]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[162], x[161], x[160], x[159], x[158], x[157], x[156], x[155]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[188], x[187], x[186], x[176], x[175], x[174], x[173], x[172]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[185], x[184], x[183], x[176], x[175], x[174], x[173], x[172]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[182], x[181], x[180], x[176], x[175], x[174], x[173], x[172]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[205], x[204], x[203], x[193], x[192], x[191], x[190], x[189]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[202], x[201], x[200], x[193], x[192], x[191], x[190], x[189]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[199], x[198], x[197], x[193], x[192], x[191], x[190], x[189]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[222], x[221], x[220], x[210], x[209], x[208], x[207], x[206]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[219], x[218], x[217], x[210], x[209], x[208], x[207], x[206]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[216], x[215], x[214], x[210], x[209], x[208], x[207], x[206]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[239], x[238], x[237], x[227], x[226], x[225], x[224], x[223]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[236], x[235], x[234], x[227], x[226], x[225], x[224], x[223]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[233], x[232], x[231], x[227], x[226], x[225], x[224], x[223]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[256], x[255], x[254], x[244], x[243], x[242], x[241], x[240]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[253], x[252], x[251], x[244], x[243], x[242], x[241], x[240]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[250], x[249], x[248], x[244], x[243], x[242], x[241], x[240]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[273], x[272], x[271], x[261], x[260], x[259], x[258], x[257]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[270], x[269], x[268], x[261], x[260], x[259], x[258], x[257]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[267], x[266], x[265], x[261], x[260], x[259], x[258], x[257]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[282], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[290], x[289], x[288], x[278], x[277], x[276], x[275], x[274]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[287], x[286], x[285], x[278], x[277], x[276], x[275], x[274]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[284], x[283], x[282], x[278], x[277], x[276], x[275], x[274]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[358], x[357], x[356], x[355], x[354], x[35], x[34], x[353], x[352], x[351], x[350], x[349], x[348], x[347], x[346], x[32], x[31], x[345], x[344], x[343], x[342], x[341], x[340], x[339], x[338], x[29], x[28], x[337], x[336], x[335], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[26], x[25], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[18], x[296], x[295], x[294], x[293], x[292], x[291]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[358], x[333], x[332], x[331], x[330], x[329], x[357], x[327], x[326], x[325], x[324], x[323], x[356], x[321], x[320], x[319], x[318], x[317], x[355], x[315], x[314], x[313], x[312], x[311], x[354], x[309], x[308], x[307], x[306], x[305], x[35], x[34], x[353], x[303], x[302], x[301], x[300], x[299], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[352], x[297], x[18], x[351], x[295], x[294], x[293], x[292], x[291]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[350], x[333], x[332], x[331], x[330], x[329], x[349], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[348], x[321], x[320], x[319], x[318], x[317], x[347], x[315], x[314], x[313], x[312], x[311], x[346], x[309], x[308], x[307], x[306], x[305], x[14], x[13], x[12], x[32], x[31], x[345], x[303], x[302], x[301], x[300], x[299], x[344], x[297], x[18], x[343], x[295], x[294], x[293], x[292], x[291]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[342], x[327], x[326], x[325], x[324], x[323], x[341], x[333], x[332], x[331], x[330], x[329], x[340], x[315], x[314], x[313], x[312], x[311], x[339], x[321], x[320], x[319], x[318], x[317], x[338], x[309], x[308], x[307], x[306], x[305], x[29], x[28], x[337], x[303], x[302], x[301], x[300], x[299], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[336], x[297], x[18], x[335], x[295], x[294], x[293], x[292], x[291]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[310], x[309], x[308], x[307], x[306], x[305], x[26], x[25], x[304], x[303], x[302], x[301], x[300], x[299], x[298], x[297], x[18], x[296], x[295], x[294], x[293], x[292], x[291]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[358], x[357], x[407], x[406], x[405], x[52], x[51], x[404], x[403], x[402], x[350], x[349], x[401], x[400], x[399], x[49], x[48], x[398], x[397], x[396], x[342], x[341], x[395], x[394], x[393], x[46], x[45], x[392], x[391], x[390], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[377], x[376], x[375], x[374], x[373], x[372], x[43], x[42], x[371], x[370], x[369], x[368], x[367], x[366], x[365], x[297], x[18], x[364], x[363], x[362], x[361], x[360], x[359]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[358], x[333], x[332], x[331], x[330], x[329], x[357], x[327], x[326], x[325], x[324], x[323], x[407], x[382], x[381], x[380], x[379], x[378], x[406], x[388], x[387], x[386], x[385], x[384], x[405], x[376], x[375], x[374], x[373], x[372], x[52], x[51], x[404], x[370], x[369], x[368], x[367], x[366], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[403], x[297], x[18], x[402], x[363], x[362], x[361], x[360], x[359]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[350], x[333], x[332], x[331], x[330], x[329], x[349], x[327], x[326], x[325], x[324], x[323], x[401], x[382], x[381], x[380], x[379], x[378], x[400], x[388], x[387], x[386], x[385], x[384], x[399], x[376], x[375], x[374], x[373], x[372], x[49], x[48], x[398], x[370], x[369], x[368], x[367], x[366], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[397], x[297], x[18], x[396], x[363], x[362], x[361], x[360], x[359]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[342], x[327], x[326], x[325], x[324], x[323], x[341], x[333], x[332], x[331], x[330], x[329], x[395], x[382], x[381], x[380], x[379], x[378], x[394], x[388], x[387], x[386], x[385], x[384], x[393], x[376], x[375], x[374], x[373], x[372], x[46], x[45], x[392], x[370], x[369], x[368], x[367], x[366], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[391], x[297], x[18], x[390], x[363], x[362], x[361], x[360], x[359]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[377], x[376], x[375], x[374], x[373], x[372], x[43], x[42], x[371], x[370], x[369], x[368], x[367], x[366], x[365], x[297], x[18], x[364], x[363], x[362], x[361], x[360], x[359]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[354], x[405], x[69], x[68], x[357], x[420], x[419], x[346], x[399], x[66], x[65], x[349], x[418], x[417], x[338], x[393], x[63], x[62], x[342], x[416], x[415], x[377], x[376], x[375], x[374], x[373], x[372], x[310], x[309], x[308], x[307], x[306], x[305], x[60], x[59], x[328], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[414], x[297], x[18], x[413], x[412], x[411], x[410], x[409], x[408]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[354], x[309], x[308], x[307], x[306], x[305], x[405], x[376], x[375], x[374], x[373], x[372], x[69], x[68], x[357], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[420], x[297], x[18], x[419], x[412], x[411], x[410], x[409], x[408]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[346], x[309], x[308], x[307], x[306], x[305], x[399], x[376], x[375], x[374], x[373], x[372], x[66], x[65], x[349], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[418], x[297], x[18], x[417], x[412], x[411], x[410], x[409], x[408]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[338], x[309], x[308], x[307], x[306], x[305], x[393], x[376], x[375], x[374], x[373], x[372], x[63], x[62], x[342], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[416], x[297], x[18], x[415], x[412], x[411], x[410], x[409], x[408]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[377], x[376], x[375], x[374], x[373], x[372], x[310], x[309], x[308], x[307], x[306], x[305], x[60], x[59], x[328], x[327], x[326], x[325], x[324], x[323], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[414], x[297], x[18], x[413], x[412], x[411], x[410], x[409], x[408]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[354], x[405], x[460], x[459], x[358], x[86], x[85], x[458], x[457], x[456], x[346], x[399], x[455], x[454], x[350], x[83], x[82], x[453], x[452], x[451], x[338], x[393], x[450], x[449], x[341], x[80], x[79], x[448], x[447], x[446], x[377], x[376], x[375], x[374], x[373], x[372], x[310], x[309], x[308], x[307], x[306], x[305], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[334], x[333], x[332], x[331], x[330], x[329], x[77], x[76], x[433], x[432], x[431], x[430], x[429], x[428], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[427], x[297], x[18], x[426], x[425], x[424], x[423], x[422], x[421]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[354], x[309], x[308], x[307], x[306], x[305], x[405], x[376], x[375], x[374], x[373], x[372], x[460], x[444], x[443], x[442], x[441], x[440], x[459], x[438], x[437], x[436], x[435], x[434], x[358], x[333], x[332], x[331], x[330], x[329], x[86], x[85], x[458], x[432], x[431], x[430], x[429], x[428], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[457], x[297], x[18], x[456], x[425], x[424], x[423], x[422], x[421]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[346], x[309], x[308], x[307], x[306], x[305], x[399], x[376], x[375], x[374], x[373], x[372], x[455], x[444], x[443], x[442], x[441], x[440], x[454], x[438], x[437], x[436], x[435], x[434], x[350], x[333], x[332], x[331], x[330], x[329], x[83], x[82], x[453], x[432], x[431], x[430], x[429], x[428], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[452], x[297], x[18], x[451], x[425], x[424], x[423], x[422], x[421]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[338], x[309], x[308], x[307], x[306], x[305], x[393], x[376], x[375], x[374], x[373], x[372], x[450], x[438], x[437], x[436], x[435], x[434], x[449], x[444], x[443], x[442], x[441], x[440], x[341], x[333], x[332], x[331], x[330], x[329], x[80], x[79], x[448], x[432], x[431], x[430], x[429], x[428], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[447], x[297], x[18], x[446], x[425], x[424], x[423], x[422], x[421]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[377], x[376], x[375], x[374], x[373], x[372], x[310], x[309], x[308], x[307], x[306], x[305], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[334], x[333], x[332], x[331], x[330], x[329], x[77], x[76], x[433], x[432], x[431], x[430], x[429], x[428], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[427], x[297], x[18], x[426], x[425], x[424], x[423], x[422], x[421]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[460], x[459], x[404], x[491], x[490], x[103], x[102], x[406], x[489], x[488], x[455], x[454], x[398], x[487], x[486], x[100], x[99], x[400], x[485], x[484], x[450], x[449], x[483], x[392], x[482], x[97], x[96], x[394], x[481], x[480], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[371], x[370], x[369], x[368], x[367], x[366], x[479], x[478], x[477], x[476], x[475], x[474], x[473], x[472], x[471], x[470], x[469], x[468], x[94], x[93], x[389], x[388], x[387], x[386], x[385], x[384], x[467], x[297], x[18], x[466], x[465], x[464], x[463], x[462], x[461]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[460], x[444], x[443], x[442], x[441], x[440], x[459], x[438], x[437], x[436], x[435], x[434], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[404], x[370], x[369], x[368], x[367], x[366], x[491], x[478], x[477], x[476], x[475], x[474], x[490], x[472], x[471], x[470], x[469], x[468], x[103], x[102], x[406], x[388], x[387], x[386], x[385], x[384], x[489], x[297], x[18], x[488], x[465], x[464], x[463], x[462], x[461]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[455], x[444], x[443], x[442], x[441], x[440], x[454], x[438], x[437], x[436], x[435], x[434], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[398], x[370], x[369], x[368], x[367], x[366], x[487], x[478], x[477], x[476], x[475], x[474], x[486], x[472], x[471], x[470], x[469], x[468], x[100], x[99], x[400], x[388], x[387], x[386], x[385], x[384], x[485], x[297], x[18], x[484], x[465], x[464], x[463], x[462], x[461]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[450], x[438], x[437], x[436], x[435], x[434], x[449], x[444], x[443], x[442], x[441], x[440], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[483], x[478], x[477], x[476], x[475], x[474], x[392], x[370], x[369], x[368], x[367], x[366], x[482], x[472], x[471], x[470], x[469], x[468], x[97], x[96], x[394], x[388], x[387], x[386], x[385], x[384], x[481], x[297], x[18], x[480], x[465], x[464], x[463], x[462], x[461]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[371], x[370], x[369], x[368], x[367], x[366], x[479], x[478], x[477], x[476], x[475], x[474], x[473], x[472], x[471], x[470], x[469], x[468], x[94], x[93], x[389], x[388], x[387], x[386], x[385], x[384], x[467], x[297], x[18], x[466], x[465], x[464], x[463], x[462], x[461]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[460], x[459], x[353], x[513], x[458], x[120], x[119], x[355], x[512], x[511], x[455], x[454], x[345], x[510], x[453], x[117], x[116], x[347], x[509], x[508], x[450], x[449], x[337], x[507], x[448], x[114], x[113], x[340], x[506], x[505], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[504], x[503], x[502], x[501], x[500], x[499], x[304], x[303], x[302], x[301], x[300], x[299], x[433], x[432], x[431], x[430], x[429], x[428], x[111], x[110], x[316], x[315], x[314], x[313], x[312], x[311], x[498], x[297], x[18], x[497], x[496], x[495], x[494], x[493], x[492]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[460], x[444], x[443], x[442], x[441], x[440], x[459], x[438], x[437], x[436], x[435], x[434], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[353], x[303], x[302], x[301], x[300], x[299], x[513], x[503], x[502], x[501], x[500], x[499], x[458], x[432], x[431], x[430], x[429], x[428], x[120], x[119], x[355], x[315], x[314], x[313], x[312], x[311], x[512], x[297], x[18], x[511], x[496], x[495], x[494], x[493], x[492]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[455], x[444], x[443], x[442], x[441], x[440], x[454], x[438], x[437], x[436], x[435], x[434], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[345], x[303], x[302], x[301], x[300], x[299], x[510], x[503], x[502], x[501], x[500], x[499], x[453], x[432], x[431], x[430], x[429], x[428], x[117], x[116], x[347], x[315], x[314], x[313], x[312], x[311], x[509], x[297], x[18], x[508], x[496], x[495], x[494], x[493], x[492]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[450], x[438], x[437], x[436], x[435], x[434], x[449], x[444], x[443], x[442], x[441], x[440], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[337], x[303], x[302], x[301], x[300], x[299], x[507], x[503], x[502], x[501], x[500], x[499], x[448], x[432], x[431], x[430], x[429], x[428], x[114], x[113], x[340], x[315], x[314], x[313], x[312], x[311], x[506], x[297], x[18], x[505], x[496], x[495], x[494], x[493], x[492]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[504], x[503], x[502], x[501], x[500], x[499], x[304], x[303], x[302], x[301], x[300], x[299], x[433], x[432], x[431], x[430], x[429], x[428], x[111], x[110], x[316], x[315], x[314], x[313], x[312], x[311], x[498], x[297], x[18], x[497], x[496], x[495], x[494], x[493], x[492]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[490], x[458], x[459], x[137], x[136], x[460], x[526], x[525], x[486], x[453], x[454], x[134], x[133], x[455], x[524], x[523], x[482], x[448], x[450], x[131], x[130], x[449], x[522], x[521], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[433], x[432], x[431], x[430], x[429], x[428], x[473], x[472], x[471], x[470], x[469], x[468], x[439], x[438], x[437], x[436], x[435], x[434], x[128], x[127], x[445], x[444], x[443], x[442], x[441], x[440], x[520], x[297], x[18], x[519], x[518], x[517], x[516], x[515], x[514]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[490], x[472], x[471], x[470], x[469], x[468], x[458], x[432], x[431], x[430], x[429], x[428], x[459], x[438], x[437], x[436], x[435], x[434], x[137], x[136], x[460], x[444], x[443], x[442], x[441], x[440], x[526], x[297], x[18], x[525], x[518], x[517], x[516], x[515], x[514]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[486], x[472], x[471], x[470], x[469], x[468], x[453], x[432], x[431], x[430], x[429], x[428], x[454], x[438], x[437], x[436], x[435], x[434], x[14], x[13], x[12], x[134], x[133], x[455], x[444], x[443], x[442], x[441], x[440], x[524], x[297], x[18], x[523], x[518], x[517], x[516], x[515], x[514]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[482], x[472], x[471], x[470], x[469], x[468], x[448], x[432], x[431], x[430], x[429], x[428], x[450], x[438], x[437], x[436], x[435], x[434], x[131], x[130], x[449], x[444], x[443], x[442], x[441], x[440], x[522], x[297], x[18], x[521], x[518], x[517], x[516], x[515], x[514]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[433], x[432], x[431], x[430], x[429], x[428], x[473], x[472], x[471], x[470], x[469], x[468], x[439], x[438], x[437], x[436], x[435], x[434], x[128], x[127], x[445], x[444], x[443], x[442], x[441], x[440], x[520], x[297], x[18], x[519], x[518], x[517], x[516], x[515], x[514]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[490], x[458], x[358], x[357], x[460], x[154], x[153], x[354], x[539], x[538], x[486], x[453], x[350], x[349], x[455], x[151], x[150], x[346], x[537], x[536], x[482], x[448], x[342], x[341], x[449], x[148], x[147], x[338], x[535], x[534], x[433], x[432], x[431], x[430], x[429], x[428], x[473], x[472], x[471], x[470], x[469], x[468], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[445], x[444], x[443], x[442], x[441], x[440], x[145], x[144], x[310], x[309], x[308], x[307], x[306], x[305], x[533], x[297], x[18], x[532], x[531], x[530], x[529], x[528], x[527]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[490], x[472], x[471], x[470], x[469], x[468], x[458], x[432], x[431], x[430], x[429], x[428], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[358], x[333], x[332], x[331], x[330], x[329], x[357], x[327], x[326], x[325], x[324], x[323], x[460], x[444], x[443], x[442], x[441], x[440], x[154], x[153], x[354], x[309], x[308], x[307], x[306], x[305], x[539], x[297], x[18], x[538], x[531], x[530], x[529], x[528], x[527]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[486], x[472], x[471], x[470], x[469], x[468], x[453], x[432], x[431], x[430], x[429], x[428], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[350], x[333], x[332], x[331], x[330], x[329], x[349], x[327], x[326], x[325], x[324], x[323], x[455], x[444], x[443], x[442], x[441], x[440], x[151], x[150], x[346], x[309], x[308], x[307], x[306], x[305], x[537], x[297], x[18], x[536], x[531], x[530], x[529], x[528], x[527]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[482], x[472], x[471], x[470], x[469], x[468], x[448], x[432], x[431], x[430], x[429], x[428], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[342], x[327], x[326], x[325], x[324], x[323], x[341], x[333], x[332], x[331], x[330], x[329], x[449], x[444], x[443], x[442], x[441], x[440], x[148], x[147], x[338], x[309], x[308], x[307], x[306], x[305], x[535], x[297], x[18], x[534], x[531], x[530], x[529], x[528], x[527]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[433], x[432], x[431], x[430], x[429], x[428], x[473], x[472], x[471], x[470], x[469], x[468], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[445], x[444], x[443], x[442], x[441], x[440], x[145], x[144], x[310], x[309], x[308], x[307], x[306], x[305], x[533], x[297], x[18], x[532], x[531], x[530], x[529], x[528], x[527]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[404], x[491], x[354], x[405], x[407], x[171], x[170], x[358], x[552], x[551], x[398], x[487], x[346], x[399], x[401], x[168], x[167], x[350], x[550], x[549], x[483], x[392], x[338], x[393], x[395], x[165], x[164], x[341], x[548], x[547], x[371], x[370], x[369], x[368], x[367], x[366], x[479], x[478], x[477], x[476], x[475], x[474], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[377], x[376], x[375], x[374], x[373], x[372], x[310], x[309], x[308], x[307], x[306], x[305], x[383], x[382], x[381], x[380], x[379], x[378], x[162], x[161], x[334], x[333], x[332], x[331], x[330], x[329], x[546], x[297], x[18], x[545], x[544], x[543], x[542], x[541], x[540]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[404], x[370], x[369], x[368], x[367], x[366], x[491], x[478], x[477], x[476], x[475], x[474], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[354], x[309], x[308], x[307], x[306], x[305], x[405], x[376], x[375], x[374], x[373], x[372], x[407], x[382], x[381], x[380], x[379], x[378], x[171], x[170], x[358], x[333], x[332], x[331], x[330], x[329], x[552], x[297], x[18], x[551], x[544], x[543], x[542], x[541], x[540]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[398], x[370], x[369], x[368], x[367], x[366], x[487], x[478], x[477], x[476], x[475], x[474], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[346], x[309], x[308], x[307], x[306], x[305], x[399], x[376], x[375], x[374], x[373], x[372], x[401], x[382], x[381], x[380], x[379], x[378], x[168], x[167], x[350], x[333], x[332], x[331], x[330], x[329], x[550], x[297], x[18], x[549], x[544], x[543], x[542], x[541], x[540]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[483], x[478], x[477], x[476], x[475], x[474], x[392], x[370], x[369], x[368], x[367], x[366], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[338], x[309], x[308], x[307], x[306], x[305], x[393], x[376], x[375], x[374], x[373], x[372], x[395], x[382], x[381], x[380], x[379], x[378], x[165], x[164], x[341], x[333], x[332], x[331], x[330], x[329], x[548], x[297], x[18], x[547], x[544], x[543], x[542], x[541], x[540]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[371], x[370], x[369], x[368], x[367], x[366], x[479], x[478], x[477], x[476], x[475], x[474], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[377], x[376], x[375], x[374], x[373], x[372], x[310], x[309], x[308], x[307], x[306], x[305], x[383], x[382], x[381], x[380], x[379], x[378], x[162], x[161], x[334], x[333], x[332], x[331], x[330], x[329], x[546], x[297], x[18], x[545], x[544], x[543], x[542], x[541], x[540]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[404], x[491], x[460], x[459], x[406], x[188], x[187], x[490], x[565], x[564], x[398], x[487], x[455], x[454], x[400], x[185], x[184], x[486], x[563], x[562], x[483], x[392], x[450], x[449], x[394], x[182], x[181], x[482], x[561], x[560], x[371], x[370], x[369], x[368], x[367], x[366], x[479], x[478], x[477], x[476], x[475], x[474], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[389], x[388], x[387], x[386], x[385], x[384], x[179], x[178], x[473], x[472], x[471], x[470], x[469], x[468], x[559], x[297], x[18], x[558], x[557], x[556], x[555], x[554], x[553]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[404], x[370], x[369], x[368], x[367], x[366], x[491], x[478], x[477], x[476], x[475], x[474], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[460], x[444], x[443], x[442], x[441], x[440], x[459], x[438], x[437], x[436], x[435], x[434], x[406], x[388], x[387], x[386], x[385], x[384], x[188], x[187], x[490], x[472], x[471], x[470], x[469], x[468], x[565], x[297], x[18], x[564], x[557], x[556], x[555], x[554], x[553]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[398], x[370], x[369], x[368], x[367], x[366], x[487], x[478], x[477], x[476], x[475], x[474], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[455], x[444], x[443], x[442], x[441], x[440], x[454], x[438], x[437], x[436], x[435], x[434], x[400], x[388], x[387], x[386], x[385], x[384], x[185], x[184], x[486], x[472], x[471], x[470], x[469], x[468], x[563], x[297], x[18], x[562], x[557], x[556], x[555], x[554], x[553]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[483], x[478], x[477], x[476], x[475], x[474], x[392], x[370], x[369], x[368], x[367], x[366], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[450], x[438], x[437], x[436], x[435], x[434], x[449], x[444], x[443], x[442], x[441], x[440], x[394], x[388], x[387], x[386], x[385], x[384], x[182], x[181], x[482], x[472], x[471], x[470], x[469], x[468], x[561], x[297], x[18], x[560], x[557], x[556], x[555], x[554], x[553]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[371], x[370], x[369], x[368], x[367], x[366], x[479], x[478], x[477], x[476], x[475], x[474], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[445], x[444], x[443], x[442], x[441], x[440], x[439], x[438], x[437], x[436], x[435], x[434], x[389], x[388], x[387], x[386], x[385], x[384], x[179], x[178], x[473], x[472], x[471], x[470], x[469], x[468], x[559], x[297], x[18], x[558], x[557], x[556], x[555], x[554], x[553]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[407], x[406], x[356], x[355], x[491], x[205], x[204], x[513], x[578], x[577], x[401], x[400], x[348], x[347], x[487], x[202], x[201], x[510], x[576], x[575], x[395], x[394], x[340], x[339], x[483], x[199], x[198], x[507], x[574], x[573], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[479], x[478], x[477], x[476], x[475], x[474], x[196], x[195], x[504], x[503], x[502], x[501], x[500], x[499], x[572], x[297], x[18], x[571], x[570], x[569], x[568], x[567], x[566]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[407], x[382], x[381], x[380], x[379], x[378], x[406], x[388], x[387], x[386], x[385], x[384], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[356], x[321], x[320], x[319], x[318], x[317], x[355], x[315], x[314], x[313], x[312], x[311], x[491], x[478], x[477], x[476], x[475], x[474], x[205], x[204], x[513], x[503], x[502], x[501], x[500], x[499], x[578], x[297], x[18], x[577], x[570], x[569], x[568], x[567], x[566]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[401], x[382], x[381], x[380], x[379], x[378], x[400], x[388], x[387], x[386], x[385], x[384], x[348], x[321], x[320], x[319], x[318], x[317], x[347], x[315], x[314], x[313], x[312], x[311], x[487], x[478], x[477], x[476], x[475], x[474], x[202], x[201], x[510], x[503], x[502], x[501], x[500], x[499], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[576], x[297], x[18], x[575], x[570], x[569], x[568], x[567], x[566]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[395], x[382], x[381], x[380], x[379], x[378], x[394], x[388], x[387], x[386], x[385], x[384], x[340], x[315], x[314], x[313], x[312], x[311], x[339], x[321], x[320], x[319], x[318], x[317], x[483], x[478], x[477], x[476], x[475], x[474], x[199], x[198], x[507], x[503], x[502], x[501], x[500], x[499], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[574], x[297], x[18], x[573], x[570], x[569], x[568], x[567], x[566]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[479], x[478], x[477], x[476], x[475], x[474], x[196], x[195], x[504], x[503], x[502], x[501], x[500], x[499], x[572], x[297], x[18], x[571], x[570], x[569], x[568], x[567], x[566]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[407], x[406], x[404], x[222], x[221], x[491], x[591], x[590], x[401], x[400], x[398], x[219], x[218], x[487], x[589], x[588], x[395], x[394], x[392], x[216], x[215], x[483], x[587], x[586], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[371], x[370], x[369], x[368], x[367], x[366], x[213], x[212], x[479], x[478], x[477], x[476], x[475], x[474], x[585], x[297], x[18], x[584], x[583], x[582], x[581], x[580], x[579]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[407], x[382], x[381], x[380], x[379], x[378], x[406], x[388], x[387], x[386], x[385], x[384], x[404], x[370], x[369], x[368], x[367], x[366], x[222], x[221], x[491], x[478], x[477], x[476], x[475], x[474], x[591], x[297], x[18], x[590], x[583], x[582], x[581], x[580], x[579]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[401], x[382], x[381], x[380], x[379], x[378], x[400], x[388], x[387], x[386], x[385], x[384], x[398], x[370], x[369], x[368], x[367], x[366], x[219], x[218], x[487], x[478], x[477], x[476], x[475], x[474], x[589], x[297], x[18], x[588], x[583], x[582], x[581], x[580], x[579]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[395], x[382], x[381], x[380], x[379], x[378], x[394], x[388], x[387], x[386], x[385], x[384], x[392], x[370], x[369], x[368], x[367], x[366], x[216], x[215], x[483], x[478], x[477], x[476], x[475], x[474], x[587], x[297], x[18], x[586], x[583], x[582], x[581], x[580], x[579]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[389], x[388], x[387], x[386], x[385], x[384], x[383], x[382], x[381], x[380], x[379], x[378], x[371], x[370], x[369], x[368], x[367], x[366], x[213], x[212], x[479], x[478], x[477], x[476], x[475], x[474], x[585], x[297], x[18], x[584], x[583], x[582], x[581], x[580], x[579]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[356], x[355], x[490], x[458], x[353], x[239], x[238], x[459], x[604], x[603], x[348], x[347], x[486], x[453], x[345], x[236], x[235], x[454], x[602], x[601], x[340], x[339], x[482], x[448], x[337], x[233], x[232], x[450], x[600], x[599], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[433], x[432], x[431], x[430], x[429], x[428], x[473], x[472], x[471], x[470], x[469], x[468], x[304], x[303], x[302], x[301], x[300], x[299], x[230], x[229], x[439], x[438], x[437], x[436], x[435], x[434], x[598], x[297], x[18], x[597], x[596], x[595], x[594], x[593], x[592]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[356], x[321], x[320], x[319], x[318], x[317], x[355], x[315], x[314], x[313], x[312], x[311], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[490], x[472], x[471], x[470], x[469], x[468], x[458], x[432], x[431], x[430], x[429], x[428], x[353], x[303], x[302], x[301], x[300], x[299], x[239], x[238], x[459], x[438], x[437], x[436], x[435], x[434], x[604], x[297], x[18], x[603], x[596], x[595], x[594], x[593], x[592]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[348], x[321], x[320], x[319], x[318], x[317], x[347], x[315], x[314], x[313], x[312], x[311], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[486], x[472], x[471], x[470], x[469], x[468], x[453], x[432], x[431], x[430], x[429], x[428], x[345], x[303], x[302], x[301], x[300], x[299], x[236], x[235], x[454], x[438], x[437], x[436], x[435], x[434], x[602], x[297], x[18], x[601], x[596], x[595], x[594], x[593], x[592]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[340], x[315], x[314], x[313], x[312], x[311], x[339], x[321], x[320], x[319], x[318], x[317], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[482], x[472], x[471], x[470], x[469], x[468], x[448], x[432], x[431], x[430], x[429], x[428], x[337], x[303], x[302], x[301], x[300], x[299], x[233], x[232], x[450], x[438], x[437], x[436], x[435], x[434], x[600], x[297], x[18], x[599], x[596], x[595], x[594], x[593], x[592]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[433], x[432], x[431], x[430], x[429], x[428], x[473], x[472], x[471], x[470], x[469], x[468], x[304], x[303], x[302], x[301], x[300], x[299], x[230], x[229], x[439], x[438], x[437], x[436], x[435], x[434], x[598], x[297], x[18], x[597], x[596], x[595], x[594], x[593], x[592]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[356], x[355], x[358], x[357], x[513], x[256], x[255], x[405], x[617], x[616], x[348], x[347], x[350], x[349], x[510], x[253], x[252], x[399], x[615], x[614], x[340], x[339], x[342], x[341], x[507], x[250], x[249], x[393], x[613], x[612], x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[504], x[503], x[502], x[501], x[500], x[499], x[247], x[246], x[377], x[376], x[375], x[374], x[373], x[372], x[611], x[297], x[18], x[610], x[609], x[608], x[607], x[606], x[605]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[356], x[321], x[320], x[319], x[318], x[317], x[355], x[315], x[314], x[313], x[312], x[311], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[358], x[333], x[332], x[331], x[330], x[329], x[357], x[327], x[326], x[325], x[324], x[323], x[513], x[503], x[502], x[501], x[500], x[499], x[256], x[255], x[405], x[376], x[375], x[374], x[373], x[372], x[617], x[297], x[18], x[616], x[609], x[608], x[607], x[606], x[605]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[348], x[321], x[320], x[319], x[318], x[317], x[347], x[315], x[314], x[313], x[312], x[311], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[350], x[333], x[332], x[331], x[330], x[329], x[349], x[327], x[326], x[325], x[324], x[323], x[510], x[503], x[502], x[501], x[500], x[499], x[253], x[252], x[399], x[376], x[375], x[374], x[373], x[372], x[615], x[297], x[18], x[614], x[609], x[608], x[607], x[606], x[605]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[340], x[315], x[314], x[313], x[312], x[311], x[339], x[321], x[320], x[319], x[318], x[317], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[342], x[327], x[326], x[325], x[324], x[323], x[341], x[333], x[332], x[331], x[330], x[329], x[507], x[503], x[502], x[501], x[500], x[499], x[250], x[249], x[393], x[376], x[375], x[374], x[373], x[372], x[613], x[297], x[18], x[612], x[609], x[608], x[607], x[606], x[605]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[322], x[321], x[320], x[319], x[318], x[317], x[316], x[315], x[314], x[313], x[312], x[311], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[334], x[333], x[332], x[331], x[330], x[329], x[328], x[327], x[326], x[325], x[324], x[323], x[504], x[503], x[502], x[501], x[500], x[499], x[247], x[246], x[377], x[376], x[375], x[374], x[373], x[372], x[611], x[297], x[18], x[610], x[609], x[608], x[607], x[606], x[605]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[353], x[513], x[404], x[491], x[355], x[273], x[272], x[407], x[630], x[629], x[345], x[510], x[398], x[487], x[347], x[270], x[269], x[401], x[628], x[627], x[337], x[507], x[483], x[392], x[340], x[267], x[266], x[395], x[626], x[625], x[504], x[503], x[502], x[501], x[500], x[499], x[304], x[303], x[302], x[301], x[300], x[299], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[371], x[370], x[369], x[368], x[367], x[366], x[479], x[478], x[477], x[476], x[475], x[474], x[316], x[315], x[314], x[313], x[312], x[311], x[264], x[263], x[383], x[382], x[381], x[380], x[379], x[378], x[624], x[297], x[18], x[623], x[622], x[621], x[620], x[619], x[618]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[353], x[303], x[302], x[301], x[300], x[299], x[513], x[503], x[502], x[501], x[500], x[499], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[404], x[370], x[369], x[368], x[367], x[366], x[491], x[478], x[477], x[476], x[475], x[474], x[355], x[315], x[314], x[313], x[312], x[311], x[273], x[272], x[407], x[382], x[381], x[380], x[379], x[378], x[630], x[297], x[18], x[629], x[622], x[621], x[620], x[619], x[618]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[345], x[303], x[302], x[301], x[300], x[299], x[510], x[503], x[502], x[501], x[500], x[499], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[398], x[370], x[369], x[368], x[367], x[366], x[487], x[478], x[477], x[476], x[475], x[474], x[347], x[315], x[314], x[313], x[312], x[311], x[270], x[269], x[401], x[382], x[381], x[380], x[379], x[378], x[628], x[297], x[18], x[627], x[622], x[621], x[620], x[619], x[618]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[337], x[303], x[302], x[301], x[300], x[299], x[507], x[503], x[502], x[501], x[500], x[499], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[483], x[478], x[477], x[476], x[475], x[474], x[392], x[370], x[369], x[368], x[367], x[366], x[340], x[315], x[314], x[313], x[312], x[311], x[267], x[266], x[395], x[382], x[381], x[380], x[379], x[378], x[626], x[297], x[18], x[625], x[622], x[621], x[620], x[619], x[618]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[504], x[503], x[502], x[501], x[500], x[499], x[304], x[303], x[302], x[301], x[300], x[299], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[371], x[370], x[369], x[368], x[367], x[366], x[479], x[478], x[477], x[476], x[475], x[474], x[316], x[315], x[314], x[313], x[312], x[311], x[264], x[263], x[383], x[382], x[381], x[380], x[379], x[378], x[624], x[297], x[18], x[623], x[622], x[621], x[620], x[619], x[618]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[353], x[513], x[290], x[289], x[356], x[643], x[642], x[345], x[510], x[287], x[286], x[348], x[641], x[640], x[337], x[507], x[284], x[283], x[339], x[639], x[638], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[504], x[503], x[502], x[501], x[500], x[499], x[304], x[303], x[302], x[301], x[300], x[299], x[281], x[280], x[322], x[321], x[320], x[319], x[318], x[317], x[637], x[297], x[18], x[636], x[635], x[634], x[633], x[632], x[631]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[353], x[303], x[302], x[301], x[300], x[299], x[513], x[503], x[502], x[501], x[500], x[499], x[290], x[289], x[356], x[321], x[320], x[319], x[318], x[317], x[643], x[297], x[18], x[642], x[635], x[634], x[633], x[632], x[631]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[345], x[303], x[302], x[301], x[300], x[299], x[510], x[503], x[502], x[501], x[500], x[499], x[287], x[286], x[348], x[321], x[320], x[319], x[318], x[317], x[641], x[297], x[18], x[640], x[635], x[634], x[633], x[632], x[631]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[337], x[303], x[302], x[301], x[300], x[299], x[507], x[503], x[502], x[501], x[500], x[499], x[284], x[283], x[339], x[321], x[320], x[319], x[318], x[317], x[639], x[297], x[18], x[638], x[635], x[634], x[633], x[632], x[631]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[504], x[503], x[502], x[501], x[500], x[499], x[304], x[303], x[302], x[301], x[300], x[299], x[281], x[280], x[322], x[321], x[320], x[319], x[318], x[317], x[637], x[297], x[18], x[636], x[635], x[634], x[633], x[632], x[631]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[532], x[538], x[536], x[534], x[531], x[530], x[529], x[528], x[527]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[536], x[532], x[538], x[534], x[531], x[530], x[529], x[528], x[527]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[536], x[532], x[538], x[534], x[531], x[530], x[529], x[528], x[527]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[538], x[532], x[536], x[531], x[530], x[529], x[528], x[527]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[532], x[538], x[536], x[534], x[531], x[530], x[529], x[528], x[527]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[610], x[616], x[614], x[612], x[609], x[608], x[607], x[606], x[605]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[614], x[610], x[616], x[612], x[609], x[608], x[607], x[606], x[605]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[614], x[610], x[616], x[612], x[609], x[608], x[607], x[606], x[605]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[616], x[610], x[614], x[609], x[608], x[607], x[606], x[605]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[610], x[616], x[614], x[612], x[609], x[608], x[607], x[606], x[605]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[413], x[419], x[417], x[415], x[412], x[411], x[410], x[409], x[408]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[417], x[413], x[419], x[415], x[412], x[411], x[410], x[409], x[408]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[417], x[413], x[419], x[415], x[412], x[411], x[410], x[409], x[408]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[419], x[413], x[417], x[412], x[411], x[410], x[409], x[408]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[413], x[419], x[417], x[415], x[412], x[411], x[410], x[409], x[408]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[545], x[551], x[549], x[547], x[544], x[543], x[542], x[541], x[540]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[549], x[545], x[551], x[547], x[544], x[543], x[542], x[541], x[540]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[549], x[545], x[551], x[547], x[544], x[543], x[542], x[541], x[540]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[551], x[545], x[549], x[544], x[543], x[542], x[541], x[540]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[545], x[551], x[549], x[547], x[544], x[543], x[542], x[541], x[540]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[558], x[564], x[562], x[560], x[557], x[556], x[555], x[554], x[553]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[562], x[558], x[564], x[560], x[557], x[556], x[555], x[554], x[553]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[562], x[558], x[564], x[560], x[557], x[556], x[555], x[554], x[553]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[564], x[558], x[562], x[557], x[556], x[555], x[554], x[553]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[558], x[564], x[562], x[560], x[557], x[556], x[555], x[554], x[553]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[426], x[456], x[451], x[446], x[425], x[424], x[423], x[422], x[421]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[451], x[426], x[456], x[446], x[425], x[424], x[423], x[422], x[421]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[451], x[426], x[456], x[446], x[425], x[424], x[423], x[422], x[421]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[456], x[426], x[451], x[425], x[424], x[423], x[422], x[421]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[426], x[456], x[451], x[446], x[425], x[424], x[423], x[422], x[421]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[597], x[603], x[601], x[599], x[596], x[595], x[594], x[593], x[592]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[601], x[597], x[603], x[599], x[596], x[595], x[594], x[593], x[592]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[601], x[597], x[603], x[599], x[596], x[595], x[594], x[593], x[592]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[603], x[597], x[601], x[596], x[595], x[594], x[593], x[592]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[597], x[603], x[601], x[599], x[596], x[595], x[594], x[593], x[592]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[519], x[525], x[523], x[521], x[518], x[517], x[516], x[515], x[514]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[523], x[519], x[525], x[521], x[518], x[517], x[516], x[515], x[514]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[523], x[519], x[525], x[521], x[518], x[517], x[516], x[515], x[514]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[525], x[519], x[523], x[518], x[517], x[516], x[515], x[514]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[519], x[525], x[523], x[521], x[518], x[517], x[516], x[515], x[514]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[623], x[629], x[627], x[625], x[622], x[621], x[620], x[619], x[618]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[627], x[623], x[629], x[625], x[622], x[621], x[620], x[619], x[618]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[627], x[623], x[629], x[625], x[622], x[621], x[620], x[619], x[618]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[629], x[623], x[627], x[622], x[621], x[620], x[619], x[618]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[623], x[629], x[627], x[625], x[622], x[621], x[620], x[619], x[618]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[466], x[488], x[484], x[480], x[465], x[464], x[463], x[462], x[461]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[484], x[466], x[488], x[480], x[465], x[464], x[463], x[462], x[461]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[484], x[466], x[488], x[480], x[465], x[464], x[463], x[462], x[461]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[488], x[466], x[484], x[465], x[464], x[463], x[462], x[461]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[466], x[488], x[484], x[480], x[465], x[464], x[463], x[462], x[461]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[584], x[590], x[588], x[586], x[583], x[582], x[581], x[580], x[579]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[588], x[584], x[590], x[586], x[583], x[582], x[581], x[580], x[579]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[588], x[584], x[590], x[586], x[583], x[582], x[581], x[580], x[579]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[590], x[584], x[588], x[583], x[582], x[581], x[580], x[579]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[584], x[590], x[588], x[586], x[583], x[582], x[581], x[580], x[579]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[364], x[402], x[396], x[390], x[363], x[362], x[361], x[360], x[359]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[396], x[364], x[402], x[390], x[363], x[362], x[361], x[360], x[359]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[396], x[364], x[402], x[390], x[363], x[362], x[361], x[360], x[359]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[402], x[364], x[396], x[363], x[362], x[361], x[360], x[359]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[364], x[402], x[396], x[390], x[363], x[362], x[361], x[360], x[359]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[296], x[351], x[343], x[335], x[295], x[294], x[293], x[292], x[291]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[343], x[296], x[351], x[335], x[295], x[294], x[293], x[292], x[291]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[343], x[296], x[351], x[335], x[295], x[294], x[293], x[292], x[291]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[351], x[296], x[343], x[295], x[294], x[293], x[292], x[291]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[296], x[351], x[343], x[335], x[295], x[294], x[293], x[292], x[291]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[571], x[577], x[575], x[573], x[570], x[569], x[568], x[567], x[566]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[575], x[571], x[577], x[573], x[570], x[569], x[568], x[567], x[566]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[575], x[571], x[577], x[573], x[570], x[569], x[568], x[567], x[566]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[577], x[571], x[575], x[570], x[569], x[568], x[567], x[566]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[571], x[577], x[575], x[573], x[570], x[569], x[568], x[567], x[566]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[497], x[511], x[508], x[505], x[496], x[495], x[494], x[493], x[492]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[508], x[497], x[511], x[505], x[496], x[495], x[494], x[493], x[492]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[508], x[497], x[511], x[505], x[496], x[495], x[494], x[493], x[492]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[511], x[497], x[508], x[496], x[495], x[494], x[493], x[492]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[497], x[511], x[508], x[505], x[496], x[495], x[494], x[493], x[492]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[636], x[642], x[640], x[638], x[635], x[634], x[633], x[632], x[631]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[640], x[636], x[642], x[638], x[635], x[634], x[633], x[632], x[631]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[640], x[636], x[642], x[638], x[635], x[634], x[633], x[632], x[631]}), .y(y[267]));
  R2ind268 R2ind268_inst(.x({x[642], x[636], x[640], x[635], x[634], x[633], x[632], x[631]}), .y(y[268]));
  R2ind269 R2ind269_inst(.x({x[636], x[642], x[640], x[638], x[635], x[634], x[633], x[632], x[631]}), .y(y[269]));
  R2ind270 R2ind270_inst(.x({x[34], x[35], x[33], x[31], x[32], x[30], x[28], x[29], x[27], x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[25], x[26], x[14], x[13], x[12], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[270]));
  R2ind271 R2ind271_inst(.x({x[34], x[35], x[14], x[13], x[12], x[33], x[23], x[22], x[21], x[20], x[19]}), .y(y[271]));
  R2ind272 R2ind272_inst(.x({x[31], x[32], x[14], x[13], x[12], x[30], x[23], x[22], x[21], x[20], x[19]}), .y(y[272]));
  R2ind273 R2ind273_inst(.x({x[28], x[29], x[14], x[13], x[12], x[27], x[23], x[22], x[21], x[20], x[19]}), .y(y[273]));
  R2ind274 R2ind274_inst(.x({x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[25], x[26], x[14], x[13], x[12], x[24], x[23], x[22], x[21], x[20], x[19]}), .y(y[274]));
  R2ind275 R2ind275_inst(.x({x[52], x[51], x[50], x[48], x[49], x[47], x[45], x[46], x[44], x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[42], x[43], x[14], x[13], x[12], x[41], x[40], x[39], x[38], x[37], x[36]}), .y(y[275]));
  R2ind276 R2ind276_inst(.x({x[14], x[13], x[12], x[52], x[51], x[50], x[40], x[39], x[38], x[37], x[36]}), .y(y[276]));
  R2ind277 R2ind277_inst(.x({x[14], x[13], x[12], x[48], x[49], x[47], x[40], x[39], x[38], x[37], x[36]}), .y(y[277]));
  R2ind278 R2ind278_inst(.x({x[14], x[13], x[12], x[45], x[46], x[44], x[40], x[39], x[38], x[37], x[36]}), .y(y[278]));
  R2ind279 R2ind279_inst(.x({x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[42], x[43], x[14], x[13], x[12], x[41], x[40], x[39], x[38], x[37], x[36]}), .y(y[279]));
  R2ind280 R2ind280_inst(.x({x[68], x[69], x[67], x[65], x[66], x[64], x[63], x[62], x[61], x[297], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[60], x[59], x[14], x[13], x[12], x[58], x[57], x[56], x[55], x[54], x[53]}), .y(y[280]));
  R2ind281 R2ind281_inst(.x({x[68], x[69], x[14], x[13], x[12], x[67], x[57], x[56], x[55], x[54], x[53]}), .y(y[281]));
  R2ind282 R2ind282_inst(.x({x[65], x[66], x[14], x[13], x[12], x[64], x[57], x[56], x[55], x[54], x[53]}), .y(y[282]));
  R2ind283 R2ind283_inst(.x({x[63], x[62], x[14], x[13], x[12], x[61], x[57], x[56], x[55], x[54], x[53]}), .y(y[283]));
  R2ind284 R2ind284_inst(.x({x[297], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[60], x[59], x[14], x[13], x[12], x[58], x[57], x[56], x[55], x[54], x[53]}), .y(y[284]));
  R2ind285 R2ind285_inst(.x({x[85], x[86], x[84], x[82], x[83], x[81], x[79], x[80], x[78], x[297], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[76], x[77], x[75], x[74], x[73], x[72], x[71], x[70]}), .y(y[285]));
  R2ind286 R2ind286_inst(.x({x[85], x[86], x[14], x[13], x[12], x[84], x[74], x[73], x[72], x[71], x[70]}), .y(y[286]));
  R2ind287 R2ind287_inst(.x({x[82], x[83], x[14], x[13], x[12], x[81], x[74], x[73], x[72], x[71], x[70]}), .y(y[287]));
  R2ind288 R2ind288_inst(.x({x[79], x[80], x[14], x[13], x[12], x[78], x[74], x[73], x[72], x[71], x[70]}), .y(y[288]));
  R2ind289 R2ind289_inst(.x({x[297], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[76], x[77], x[75], x[74], x[73], x[72], x[71], x[70]}), .y(y[289]));
  R2ind290 R2ind290_inst(.x({x[102], x[103], x[101], x[99], x[100], x[98], x[96], x[97], x[95], x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[14], x[13], x[12], x[93], x[94], x[92], x[91], x[90], x[89], x[88], x[87]}), .y(y[290]));
  R2ind291 R2ind291_inst(.x({x[14], x[13], x[12], x[102], x[103], x[101], x[91], x[90], x[89], x[88], x[87]}), .y(y[291]));
  R2ind292 R2ind292_inst(.x({x[14], x[13], x[12], x[99], x[100], x[98], x[91], x[90], x[89], x[88], x[87]}), .y(y[292]));
  R2ind293 R2ind293_inst(.x({x[14], x[13], x[12], x[96], x[97], x[95], x[91], x[90], x[89], x[88], x[87]}), .y(y[293]));
  R2ind294 R2ind294_inst(.x({x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[14], x[13], x[12], x[93], x[94], x[92], x[91], x[90], x[89], x[88], x[87]}), .y(y[294]));
  R2ind295 R2ind295_inst(.x({x[119], x[120], x[118], x[116], x[117], x[115], x[113], x[114], x[112], x[11], x[10], x[9], x[17], x[16], x[15], x[297], x[8], x[7], x[6], x[14], x[13], x[12], x[110], x[111], x[109], x[108], x[107], x[106], x[105], x[104]}), .y(y[295]));
  R2ind296 R2ind296_inst(.x({x[14], x[13], x[12], x[119], x[120], x[118], x[108], x[107], x[106], x[105], x[104]}), .y(y[296]));
  R2ind297 R2ind297_inst(.x({x[14], x[13], x[12], x[116], x[117], x[115], x[108], x[107], x[106], x[105], x[104]}), .y(y[297]));
  R2ind298 R2ind298_inst(.x({x[14], x[13], x[12], x[113], x[114], x[112], x[108], x[107], x[106], x[105], x[104]}), .y(y[298]));
  R2ind299 R2ind299_inst(.x({x[11], x[10], x[9], x[17], x[16], x[15], x[297], x[8], x[7], x[6], x[14], x[13], x[12], x[110], x[111], x[109], x[108], x[107], x[106], x[105], x[104]}), .y(y[299]));
  R2ind300 R2ind300_inst(.x({x[136], x[137], x[135], x[133], x[134], x[132], x[130], x[131], x[129], x[297], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[14], x[13], x[12], x[127], x[128], x[126], x[125], x[124], x[123], x[122], x[121]}), .y(y[300]));
  R2ind301 R2ind301_inst(.x({x[14], x[13], x[12], x[136], x[137], x[135], x[125], x[124], x[123], x[122], x[121]}), .y(y[301]));
  R2ind302 R2ind302_inst(.x({x[133], x[134], x[14], x[13], x[12], x[132], x[125], x[124], x[123], x[122], x[121]}), .y(y[302]));
  R2ind303 R2ind303_inst(.x({x[14], x[13], x[12], x[130], x[131], x[129], x[125], x[124], x[123], x[122], x[121]}), .y(y[303]));
  R2ind304 R2ind304_inst(.x({x[297], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[14], x[13], x[12], x[127], x[128], x[126], x[125], x[124], x[123], x[122], x[121]}), .y(y[304]));
  R2ind305 R2ind305_inst(.x({x[153], x[154], x[152], x[150], x[151], x[149], x[147], x[148], x[146], x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[14], x[13], x[12], x[144], x[145], x[143], x[142], x[141], x[140], x[139], x[138]}), .y(y[305]));
  R2ind306 R2ind306_inst(.x({x[14], x[13], x[12], x[153], x[154], x[152], x[142], x[141], x[140], x[139], x[138]}), .y(y[306]));
  R2ind307 R2ind307_inst(.x({x[14], x[13], x[12], x[150], x[151], x[149], x[142], x[141], x[140], x[139], x[138]}), .y(y[307]));
  R2ind308 R2ind308_inst(.x({x[14], x[13], x[12], x[147], x[148], x[146], x[142], x[141], x[140], x[139], x[138]}), .y(y[308]));
  R2ind309 R2ind309_inst(.x({x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[14], x[13], x[12], x[144], x[145], x[143], x[142], x[141], x[140], x[139], x[138]}), .y(y[309]));
  R2ind310 R2ind310_inst(.x({x[170], x[171], x[169], x[167], x[168], x[166], x[164], x[165], x[163], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[161], x[162], x[160], x[159], x[158], x[157], x[156], x[155]}), .y(y[310]));
  R2ind311 R2ind311_inst(.x({x[14], x[13], x[12], x[170], x[171], x[169], x[159], x[158], x[157], x[156], x[155]}), .y(y[311]));
  R2ind312 R2ind312_inst(.x({x[14], x[13], x[12], x[167], x[168], x[166], x[159], x[158], x[157], x[156], x[155]}), .y(y[312]));
  R2ind313 R2ind313_inst(.x({x[14], x[13], x[12], x[164], x[165], x[163], x[159], x[158], x[157], x[156], x[155]}), .y(y[313]));
  R2ind314 R2ind314_inst(.x({x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[11], x[10], x[9], x[14], x[13], x[12], x[161], x[162], x[160], x[159], x[158], x[157], x[156], x[155]}), .y(y[314]));
  R2ind315 R2ind315_inst(.x({x[188], x[187], x[186], x[185], x[184], x[183], x[182], x[181], x[180], x[11], x[10], x[9], x[297], x[8], x[7], x[6], x[17], x[16], x[15], x[14], x[13], x[12], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172]}), .y(y[315]));
  R2ind316 R2ind316_inst(.x({x[14], x[13], x[12], x[188], x[187], x[186], x[176], x[175], x[174], x[173], x[172]}), .y(y[316]));
  R2ind317 R2ind317_inst(.x({x[14], x[13], x[12], x[185], x[184], x[183], x[176], x[175], x[174], x[173], x[172]}), .y(y[317]));
  R2ind318 R2ind318_inst(.x({x[14], x[13], x[12], x[182], x[181], x[180], x[176], x[175], x[174], x[173], x[172]}), .y(y[318]));
  R2ind319 R2ind319_inst(.x({x[11], x[10], x[9], x[297], x[8], x[7], x[6], x[17], x[16], x[15], x[14], x[13], x[12], x[179], x[178], x[177], x[176], x[175], x[174], x[173], x[172]}), .y(y[319]));
  R2ind320 R2ind320_inst(.x({x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[14], x[13], x[12], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189]}), .y(y[320]));
  R2ind321 R2ind321_inst(.x({x[14], x[13], x[12], x[205], x[204], x[203], x[193], x[192], x[191], x[190], x[189]}), .y(y[321]));
  R2ind322 R2ind322_inst(.x({x[14], x[13], x[12], x[202], x[201], x[200], x[193], x[192], x[191], x[190], x[189]}), .y(y[322]));
  R2ind323 R2ind323_inst(.x({x[14], x[13], x[12], x[199], x[198], x[197], x[193], x[192], x[191], x[190], x[189]}), .y(y[323]));
  R2ind324 R2ind324_inst(.x({x[11], x[10], x[9], x[297], x[17], x[16], x[15], x[8], x[7], x[6], x[14], x[13], x[12], x[196], x[195], x[194], x[193], x[192], x[191], x[190], x[189]}), .y(y[324]));
  R2ind325 R2ind325_inst(.x({x[222], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[17], x[16], x[15], x[297], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206]}), .y(y[325]));
  R2ind326 R2ind326_inst(.x({x[14], x[13], x[12], x[222], x[221], x[220], x[210], x[209], x[208], x[207], x[206]}), .y(y[326]));
  R2ind327 R2ind327_inst(.x({x[14], x[13], x[12], x[219], x[218], x[217], x[210], x[209], x[208], x[207], x[206]}), .y(y[327]));
  R2ind328 R2ind328_inst(.x({x[14], x[13], x[12], x[216], x[215], x[214], x[210], x[209], x[208], x[207], x[206]}), .y(y[328]));
  R2ind329 R2ind329_inst(.x({x[17], x[16], x[15], x[297], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206]}), .y(y[329]));
  R2ind330 R2ind330_inst(.x({x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[11], x[10], x[9], x[17], x[16], x[15], x[297], x[8], x[7], x[6], x[14], x[13], x[12], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223]}), .y(y[330]));
  R2ind331 R2ind331_inst(.x({x[14], x[13], x[12], x[239], x[238], x[237], x[227], x[226], x[225], x[224], x[223]}), .y(y[331]));
  R2ind332 R2ind332_inst(.x({x[14], x[13], x[12], x[236], x[235], x[234], x[227], x[226], x[225], x[224], x[223]}), .y(y[332]));
  R2ind333 R2ind333_inst(.x({x[14], x[13], x[12], x[233], x[232], x[231], x[227], x[226], x[225], x[224], x[223]}), .y(y[333]));
  R2ind334 R2ind334_inst(.x({x[11], x[10], x[9], x[17], x[16], x[15], x[297], x[8], x[7], x[6], x[14], x[13], x[12], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223]}), .y(y[334]));
  R2ind335 R2ind335_inst(.x({x[256], x[255], x[254], x[253], x[252], x[251], x[250], x[249], x[248], x[11], x[10], x[9], x[297], x[8], x[7], x[6], x[17], x[16], x[15], x[14], x[13], x[12], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240]}), .y(y[335]));
  R2ind336 R2ind336_inst(.x({x[14], x[13], x[12], x[256], x[255], x[254], x[244], x[243], x[242], x[241], x[240]}), .y(y[336]));
  R2ind337 R2ind337_inst(.x({x[14], x[13], x[12], x[253], x[252], x[251], x[244], x[243], x[242], x[241], x[240]}), .y(y[337]));
  R2ind338 R2ind338_inst(.x({x[14], x[13], x[12], x[250], x[249], x[248], x[244], x[243], x[242], x[241], x[240]}), .y(y[338]));
  R2ind339 R2ind339_inst(.x({x[11], x[10], x[9], x[297], x[8], x[7], x[6], x[17], x[16], x[15], x[14], x[13], x[12], x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240]}), .y(y[339]));
  R2ind340 R2ind340_inst(.x({x[273], x[272], x[271], x[270], x[269], x[268], x[267], x[266], x[265], x[11], x[10], x[9], x[17], x[16], x[15], x[297], x[8], x[7], x[6], x[14], x[13], x[12], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[340]));
  R2ind341 R2ind341_inst(.x({x[14], x[13], x[12], x[273], x[272], x[271], x[261], x[260], x[259], x[258], x[257]}), .y(y[341]));
  R2ind342 R2ind342_inst(.x({x[14], x[13], x[12], x[270], x[269], x[268], x[261], x[260], x[259], x[258], x[257]}), .y(y[342]));
  R2ind343 R2ind343_inst(.x({x[14], x[13], x[12], x[267], x[266], x[265], x[261], x[260], x[259], x[258], x[257]}), .y(y[343]));
  R2ind344 R2ind344_inst(.x({x[11], x[10], x[9], x[17], x[16], x[15], x[297], x[8], x[7], x[6], x[14], x[13], x[12], x[264], x[263], x[262], x[261], x[260], x[259], x[258], x[257]}), .y(y[344]));
  R2ind345 R2ind345_inst(.x({x[290], x[289], x[288], x[287], x[286], x[285], x[284], x[283], x[282], x[11], x[10], x[9], x[17], x[16], x[15], x[297], x[8], x[7], x[6], x[14], x[13], x[12], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274]}), .y(y[345]));
  R2ind346 R2ind346_inst(.x({x[14], x[13], x[12], x[290], x[289], x[288], x[278], x[277], x[276], x[275], x[274]}), .y(y[346]));
  R2ind347 R2ind347_inst(.x({x[14], x[13], x[12], x[287], x[286], x[285], x[278], x[277], x[276], x[275], x[274]}), .y(y[347]));
  R2ind348 R2ind348_inst(.x({x[14], x[13], x[12], x[284], x[283], x[282], x[278], x[277], x[276], x[275], x[274]}), .y(y[348]));
  R2ind349 R2ind349_inst(.x({x[11], x[10], x[9], x[17], x[16], x[15], x[297], x[8], x[7], x[6], x[14], x[13], x[12], x[281], x[280], x[279], x[278], x[277], x[276], x[275], x[274]}), .y(y[349]));
  R2ind350 R2ind350_inst(.x({x[652], x[152], x[651], x[149], x[650], x[146], x[649], x[648], x[647], x[646], x[645], x[644], x[143], x[142], x[141], x[140], x[139], x[138], x[297]}), .y(y[350]));
  R2ind351 R2ind351_inst(.x({x[652], x[648], x[647], x[646], x[645], x[644], x[152], x[142], x[141], x[140], x[139], x[138], x[297]}), .y(y[351]));
  R2ind352 R2ind352_inst(.x({x[651], x[648], x[647], x[646], x[645], x[644], x[149], x[142], x[141], x[140], x[139], x[138], x[297]}), .y(y[352]));
  R2ind353 R2ind353_inst(.x({x[650], x[648], x[647], x[646], x[645], x[644], x[146], x[142], x[141], x[140], x[139], x[138], x[297]}), .y(y[353]));
  R2ind354 R2ind354_inst(.x({x[649], x[648], x[647], x[646], x[645], x[644], x[143], x[142], x[141], x[140], x[139], x[138], x[297]}), .y(y[354]));
  R2ind355 R2ind355_inst(.x({x[661], x[254], x[660], x[251], x[659], x[248], x[658], x[657], x[656], x[655], x[654], x[653], x[245], x[244], x[243], x[242], x[241], x[240], x[297]}), .y(y[355]));
  R2ind356 R2ind356_inst(.x({x[661], x[657], x[656], x[655], x[654], x[653], x[254], x[244], x[243], x[242], x[241], x[240], x[297]}), .y(y[356]));
  R2ind357 R2ind357_inst(.x({x[660], x[657], x[656], x[655], x[654], x[653], x[251], x[244], x[243], x[242], x[241], x[240], x[297]}), .y(y[357]));
  R2ind358 R2ind358_inst(.x({x[659], x[657], x[656], x[655], x[654], x[653], x[248], x[244], x[243], x[242], x[241], x[240], x[297]}), .y(y[358]));
  R2ind359 R2ind359_inst(.x({x[658], x[657], x[656], x[655], x[654], x[653], x[245], x[244], x[243], x[242], x[241], x[240], x[297]}), .y(y[359]));
  R2ind360 R2ind360_inst(.x({x[670], x[67], x[669], x[64], x[668], x[61], x[667], x[666], x[665], x[664], x[663], x[662], x[58], x[57], x[56], x[55], x[54], x[53], x[297]}), .y(y[360]));
  R2ind361 R2ind361_inst(.x({x[670], x[666], x[665], x[664], x[663], x[662], x[67], x[57], x[56], x[55], x[54], x[53], x[297]}), .y(y[361]));
  R2ind362 R2ind362_inst(.x({x[669], x[666], x[665], x[664], x[663], x[662], x[64], x[57], x[56], x[55], x[54], x[53], x[297]}), .y(y[362]));
  R2ind363 R2ind363_inst(.x({x[668], x[666], x[665], x[664], x[663], x[662], x[61], x[57], x[56], x[55], x[54], x[53], x[297]}), .y(y[363]));
  R2ind364 R2ind364_inst(.x({x[667], x[666], x[665], x[664], x[663], x[662], x[58], x[57], x[56], x[55], x[54], x[53], x[297]}), .y(y[364]));
  R2ind365 R2ind365_inst(.x({x[679], x[169], x[678], x[166], x[677], x[163], x[676], x[675], x[674], x[673], x[672], x[671], x[160], x[159], x[158], x[157], x[156], x[155], x[297]}), .y(y[365]));
  R2ind366 R2ind366_inst(.x({x[679], x[675], x[674], x[673], x[672], x[671], x[169], x[159], x[158], x[157], x[156], x[155], x[297]}), .y(y[366]));
  R2ind367 R2ind367_inst(.x({x[678], x[675], x[674], x[673], x[672], x[671], x[166], x[159], x[158], x[157], x[156], x[155], x[297]}), .y(y[367]));
  R2ind368 R2ind368_inst(.x({x[677], x[675], x[674], x[673], x[672], x[671], x[163], x[159], x[158], x[157], x[156], x[155], x[297]}), .y(y[368]));
  R2ind369 R2ind369_inst(.x({x[676], x[675], x[674], x[673], x[672], x[671], x[160], x[159], x[158], x[157], x[156], x[155], x[297]}), .y(y[369]));
  R2ind370 R2ind370_inst(.x({x[688], x[186], x[687], x[183], x[686], x[180], x[685], x[684], x[683], x[682], x[681], x[680], x[177], x[176], x[175], x[174], x[173], x[172], x[297]}), .y(y[370]));
  R2ind371 R2ind371_inst(.x({x[688], x[684], x[683], x[682], x[681], x[680], x[186], x[176], x[175], x[174], x[173], x[172], x[297]}), .y(y[371]));
  R2ind372 R2ind372_inst(.x({x[687], x[684], x[683], x[682], x[681], x[680], x[183], x[176], x[175], x[174], x[173], x[172], x[297]}), .y(y[372]));
  R2ind373 R2ind373_inst(.x({x[686], x[684], x[683], x[682], x[681], x[680], x[180], x[176], x[175], x[174], x[173], x[172], x[297]}), .y(y[373]));
  R2ind374 R2ind374_inst(.x({x[685], x[684], x[683], x[682], x[681], x[680], x[177], x[176], x[175], x[174], x[173], x[172], x[297]}), .y(y[374]));
  R2ind375 R2ind375_inst(.x({x[697], x[84], x[696], x[81], x[695], x[78], x[694], x[693], x[692], x[691], x[690], x[689], x[75], x[74], x[73], x[72], x[71], x[70], x[297]}), .y(y[375]));
  R2ind376 R2ind376_inst(.x({x[697], x[693], x[692], x[691], x[690], x[689], x[84], x[74], x[73], x[72], x[71], x[70], x[297]}), .y(y[376]));
  R2ind377 R2ind377_inst(.x({x[696], x[693], x[692], x[691], x[690], x[689], x[81], x[74], x[73], x[72], x[71], x[70], x[297]}), .y(y[377]));
  R2ind378 R2ind378_inst(.x({x[695], x[693], x[692], x[691], x[690], x[689], x[78], x[74], x[73], x[72], x[71], x[70], x[297]}), .y(y[378]));
  R2ind379 R2ind379_inst(.x({x[694], x[693], x[692], x[691], x[690], x[689], x[75], x[74], x[73], x[72], x[71], x[70], x[297]}), .y(y[379]));
  R2ind380 R2ind380_inst(.x({x[706], x[237], x[705], x[234], x[704], x[231], x[703], x[702], x[701], x[700], x[699], x[698], x[228], x[227], x[226], x[225], x[224], x[223], x[297]}), .y(y[380]));
  R2ind381 R2ind381_inst(.x({x[706], x[702], x[701], x[700], x[699], x[698], x[237], x[227], x[226], x[225], x[224], x[223], x[297]}), .y(y[381]));
  R2ind382 R2ind382_inst(.x({x[705], x[702], x[701], x[700], x[699], x[698], x[234], x[227], x[226], x[225], x[224], x[223], x[297]}), .y(y[382]));
  R2ind383 R2ind383_inst(.x({x[704], x[702], x[701], x[700], x[699], x[698], x[231], x[227], x[226], x[225], x[224], x[223], x[297]}), .y(y[383]));
  R2ind384 R2ind384_inst(.x({x[703], x[702], x[701], x[700], x[699], x[698], x[228], x[227], x[226], x[225], x[224], x[223], x[297]}), .y(y[384]));
  R2ind385 R2ind385_inst(.x({x[715], x[135], x[714], x[132], x[713], x[129], x[712], x[711], x[710], x[709], x[708], x[707], x[126], x[125], x[124], x[123], x[122], x[121], x[297]}), .y(y[385]));
  R2ind386 R2ind386_inst(.x({x[715], x[711], x[710], x[709], x[708], x[707], x[135], x[125], x[124], x[123], x[122], x[121], x[297]}), .y(y[386]));
  R2ind387 R2ind387_inst(.x({x[714], x[711], x[710], x[709], x[708], x[707], x[132], x[125], x[124], x[123], x[122], x[121], x[297]}), .y(y[387]));
  R2ind388 R2ind388_inst(.x({x[713], x[711], x[710], x[709], x[708], x[707], x[129], x[125], x[124], x[123], x[122], x[121], x[297]}), .y(y[388]));
  R2ind389 R2ind389_inst(.x({x[712], x[711], x[710], x[709], x[708], x[707], x[126], x[125], x[124], x[123], x[122], x[121], x[297]}), .y(y[389]));
  R2ind390 R2ind390_inst(.x({x[724], x[271], x[723], x[268], x[722], x[265], x[721], x[720], x[719], x[718], x[717], x[716], x[262], x[261], x[260], x[259], x[258], x[257], x[297]}), .y(y[390]));
  R2ind391 R2ind391_inst(.x({x[724], x[720], x[719], x[718], x[717], x[716], x[271], x[261], x[260], x[259], x[258], x[257], x[297]}), .y(y[391]));
  R2ind392 R2ind392_inst(.x({x[723], x[720], x[719], x[718], x[717], x[716], x[268], x[261], x[260], x[259], x[258], x[257], x[297]}), .y(y[392]));
  R2ind393 R2ind393_inst(.x({x[722], x[720], x[719], x[718], x[717], x[716], x[265], x[261], x[260], x[259], x[258], x[257], x[297]}), .y(y[393]));
  R2ind394 R2ind394_inst(.x({x[721], x[720], x[719], x[718], x[717], x[716], x[262], x[261], x[260], x[259], x[258], x[257], x[297]}), .y(y[394]));
  R2ind395 R2ind395_inst(.x({x[733], x[101], x[732], x[98], x[731], x[95], x[730], x[729], x[728], x[727], x[726], x[725], x[92], x[91], x[90], x[89], x[88], x[87], x[297]}), .y(y[395]));
  R2ind396 R2ind396_inst(.x({x[733], x[729], x[728], x[727], x[726], x[725], x[101], x[91], x[90], x[89], x[88], x[87], x[297]}), .y(y[396]));
  R2ind397 R2ind397_inst(.x({x[732], x[729], x[728], x[727], x[726], x[725], x[98], x[91], x[90], x[89], x[88], x[87], x[297]}), .y(y[397]));
  R2ind398 R2ind398_inst(.x({x[731], x[729], x[728], x[727], x[726], x[725], x[95], x[91], x[90], x[89], x[88], x[87], x[297]}), .y(y[398]));
  R2ind399 R2ind399_inst(.x({x[730], x[729], x[728], x[727], x[726], x[725], x[92], x[91], x[90], x[89], x[88], x[87], x[297]}), .y(y[399]));
  R2ind400 R2ind400_inst(.x({x[742], x[220], x[741], x[217], x[740], x[214], x[739], x[738], x[737], x[736], x[735], x[734], x[211], x[210], x[209], x[208], x[207], x[206], x[297]}), .y(y[400]));
  R2ind401 R2ind401_inst(.x({x[742], x[738], x[737], x[736], x[735], x[734], x[220], x[210], x[209], x[208], x[207], x[206], x[297]}), .y(y[401]));
  R2ind402 R2ind402_inst(.x({x[741], x[738], x[737], x[736], x[735], x[734], x[217], x[210], x[209], x[208], x[207], x[206], x[297]}), .y(y[402]));
  R2ind403 R2ind403_inst(.x({x[740], x[738], x[737], x[736], x[735], x[734], x[214], x[210], x[209], x[208], x[207], x[206], x[297]}), .y(y[403]));
  R2ind404 R2ind404_inst(.x({x[739], x[738], x[737], x[736], x[735], x[734], x[211], x[210], x[209], x[208], x[207], x[206], x[297]}), .y(y[404]));
  R2ind405 R2ind405_inst(.x({x[751], x[50], x[750], x[47], x[749], x[44], x[748], x[747], x[746], x[745], x[744], x[743], x[41], x[40], x[39], x[38], x[37], x[36], x[297]}), .y(y[405]));
  R2ind406 R2ind406_inst(.x({x[751], x[747], x[746], x[745], x[744], x[743], x[50], x[40], x[39], x[38], x[37], x[36], x[297]}), .y(y[406]));
  R2ind407 R2ind407_inst(.x({x[750], x[747], x[746], x[745], x[744], x[743], x[47], x[40], x[39], x[38], x[37], x[36], x[297]}), .y(y[407]));
  R2ind408 R2ind408_inst(.x({x[749], x[747], x[746], x[745], x[744], x[743], x[44], x[40], x[39], x[38], x[37], x[36], x[297]}), .y(y[408]));
  R2ind409 R2ind409_inst(.x({x[748], x[747], x[746], x[745], x[744], x[743], x[41], x[40], x[39], x[38], x[37], x[36], x[297]}), .y(y[409]));
  R2ind410 R2ind410_inst(.x({x[760], x[33], x[759], x[30], x[758], x[27], x[757], x[756], x[755], x[754], x[753], x[752], x[24], x[23], x[22], x[21], x[20], x[19], x[297]}), .y(y[410]));
  R2ind411 R2ind411_inst(.x({x[760], x[756], x[755], x[754], x[753], x[752], x[33], x[23], x[22], x[21], x[20], x[19], x[297]}), .y(y[411]));
  R2ind412 R2ind412_inst(.x({x[759], x[756], x[755], x[754], x[753], x[752], x[30], x[23], x[22], x[21], x[20], x[19], x[297]}), .y(y[412]));
  R2ind413 R2ind413_inst(.x({x[758], x[756], x[755], x[754], x[753], x[752], x[27], x[23], x[22], x[21], x[20], x[19], x[297]}), .y(y[413]));
  R2ind414 R2ind414_inst(.x({x[757], x[756], x[755], x[754], x[753], x[752], x[24], x[23], x[22], x[21], x[20], x[19], x[297]}), .y(y[414]));
  R2ind415 R2ind415_inst(.x({x[769], x[203], x[768], x[200], x[767], x[197], x[766], x[765], x[764], x[763], x[762], x[761], x[194], x[193], x[192], x[191], x[190], x[189], x[297]}), .y(y[415]));
  R2ind416 R2ind416_inst(.x({x[769], x[765], x[764], x[763], x[762], x[761], x[203], x[193], x[192], x[191], x[190], x[189], x[297]}), .y(y[416]));
  R2ind417 R2ind417_inst(.x({x[768], x[765], x[764], x[763], x[762], x[761], x[200], x[193], x[192], x[191], x[190], x[189], x[297]}), .y(y[417]));
  R2ind418 R2ind418_inst(.x({x[767], x[765], x[764], x[763], x[762], x[761], x[197], x[193], x[192], x[191], x[190], x[189], x[297]}), .y(y[418]));
  R2ind419 R2ind419_inst(.x({x[766], x[765], x[764], x[763], x[762], x[761], x[194], x[193], x[192], x[191], x[190], x[189], x[297]}), .y(y[419]));
  R2ind420 R2ind420_inst(.x({x[778], x[118], x[777], x[115], x[776], x[112], x[775], x[774], x[773], x[772], x[771], x[770], x[109], x[108], x[107], x[106], x[105], x[104], x[297]}), .y(y[420]));
  R2ind421 R2ind421_inst(.x({x[778], x[774], x[773], x[772], x[771], x[770], x[118], x[108], x[107], x[106], x[105], x[104], x[297]}), .y(y[421]));
  R2ind422 R2ind422_inst(.x({x[777], x[774], x[773], x[772], x[771], x[770], x[115], x[108], x[107], x[106], x[105], x[104], x[297]}), .y(y[422]));
  R2ind423 R2ind423_inst(.x({x[776], x[774], x[773], x[772], x[771], x[770], x[112], x[108], x[107], x[106], x[105], x[104], x[297]}), .y(y[423]));
  R2ind424 R2ind424_inst(.x({x[775], x[774], x[773], x[772], x[771], x[770], x[109], x[108], x[107], x[106], x[105], x[104], x[297]}), .y(y[424]));
  R2ind425 R2ind425_inst(.x({x[787], x[288], x[786], x[285], x[785], x[282], x[784], x[783], x[782], x[781], x[780], x[779], x[279], x[278], x[277], x[276], x[275], x[274], x[297]}), .y(y[425]));
  R2ind426 R2ind426_inst(.x({x[787], x[783], x[782], x[781], x[780], x[779], x[288], x[278], x[277], x[276], x[275], x[274], x[297]}), .y(y[426]));
  R2ind427 R2ind427_inst(.x({x[786], x[783], x[782], x[781], x[780], x[779], x[285], x[278], x[277], x[276], x[275], x[274], x[297]}), .y(y[427]));
  R2ind428 R2ind428_inst(.x({x[785], x[783], x[782], x[781], x[780], x[779], x[282], x[278], x[277], x[276], x[275], x[274], x[297]}), .y(y[428]));
  R2ind429 R2ind429_inst(.x({x[784], x[783], x[782], x[781], x[780], x[779], x[279], x[278], x[277], x[276], x[275], x[274], x[297]}), .y(y[429]));
endmodule

