/* modified netlist. Source: module sbox in file Designs/AESSbox/lookup/AGEMA/sbox.v */
/* clock gating is added to the circuit, the latency increased 34 time(s)  */

module sbox_GHPC_ClockGating_d1 (SI_s0, clk, SI_s1, Fresh, rst, SO_s0, SO_s1, Synch);
    input [7:0] SI_s0 ;
    input clk ;
    input [7:0] SI_s1 ;
    input rst ;
    input [867:0] Fresh ;
    output [7:0] SO_s0 ;
    output [7:0] SO_s1 ;
    output Synch ;
    wire N169 ;
    wire N277 ;
    wire N379 ;
    wire N470 ;
    wire N563 ;
    wire N639 ;
    wire N723 ;
    wire N789 ;
    wire n1922 ;
    wire n1923 ;
    wire n1924 ;
    wire n1925 ;
    wire n1926 ;
    wire n1927 ;
    wire n1928 ;
    wire n1929 ;
    wire n1930 ;
    wire n1931 ;
    wire n1932 ;
    wire n1933 ;
    wire n1934 ;
    wire n1935 ;
    wire n1936 ;
    wire n1937 ;
    wire n1938 ;
    wire n1939 ;
    wire n1940 ;
    wire n1941 ;
    wire n1942 ;
    wire n1943 ;
    wire n1944 ;
    wire n1945 ;
    wire n1946 ;
    wire n1947 ;
    wire n1948 ;
    wire n1949 ;
    wire n1950 ;
    wire n1951 ;
    wire n1952 ;
    wire n1953 ;
    wire n1954 ;
    wire n1955 ;
    wire n1956 ;
    wire n1957 ;
    wire n1958 ;
    wire n1959 ;
    wire n1960 ;
    wire n1961 ;
    wire n1962 ;
    wire n1963 ;
    wire n1964 ;
    wire n1965 ;
    wire n1966 ;
    wire n1967 ;
    wire n1968 ;
    wire n1969 ;
    wire n1970 ;
    wire n1971 ;
    wire n1972 ;
    wire n1973 ;
    wire n1974 ;
    wire n1975 ;
    wire n1976 ;
    wire n1977 ;
    wire n1978 ;
    wire n1979 ;
    wire n1980 ;
    wire n1981 ;
    wire n1982 ;
    wire n1983 ;
    wire n1984 ;
    wire n1985 ;
    wire n1986 ;
    wire n1987 ;
    wire n1988 ;
    wire n1989 ;
    wire n1990 ;
    wire n1991 ;
    wire n1992 ;
    wire n1993 ;
    wire n1994 ;
    wire n1995 ;
    wire n1996 ;
    wire n1997 ;
    wire n1998 ;
    wire n1999 ;
    wire n2000 ;
    wire n2001 ;
    wire n2002 ;
    wire n2003 ;
    wire n2004 ;
    wire n2005 ;
    wire n2006 ;
    wire n2007 ;
    wire n2008 ;
    wire n2009 ;
    wire n2010 ;
    wire n2011 ;
    wire n2012 ;
    wire n2013 ;
    wire n2014 ;
    wire n2015 ;
    wire n2016 ;
    wire n2017 ;
    wire n2018 ;
    wire n2019 ;
    wire n2020 ;
    wire n2021 ;
    wire n2022 ;
    wire n2023 ;
    wire n2024 ;
    wire n2025 ;
    wire n2026 ;
    wire n2027 ;
    wire n2028 ;
    wire n2029 ;
    wire n2030 ;
    wire n2031 ;
    wire n2032 ;
    wire n2033 ;
    wire n2034 ;
    wire n2035 ;
    wire n2036 ;
    wire n2037 ;
    wire n2038 ;
    wire n2039 ;
    wire n2040 ;
    wire n2041 ;
    wire n2042 ;
    wire n2043 ;
    wire n2044 ;
    wire n2045 ;
    wire n2046 ;
    wire n2047 ;
    wire n2048 ;
    wire n2049 ;
    wire n2050 ;
    wire n2051 ;
    wire n2052 ;
    wire n2053 ;
    wire n2054 ;
    wire n2055 ;
    wire n2056 ;
    wire n2057 ;
    wire n2058 ;
    wire n2059 ;
    wire n2060 ;
    wire n2061 ;
    wire n2062 ;
    wire n2063 ;
    wire n2064 ;
    wire n2065 ;
    wire n2066 ;
    wire n2067 ;
    wire n2068 ;
    wire n2069 ;
    wire n2070 ;
    wire n2071 ;
    wire n2072 ;
    wire n2073 ;
    wire n2074 ;
    wire n2075 ;
    wire n2076 ;
    wire n2077 ;
    wire n2078 ;
    wire n2079 ;
    wire n2080 ;
    wire n2081 ;
    wire n2082 ;
    wire n2083 ;
    wire n2084 ;
    wire n2085 ;
    wire n2086 ;
    wire n2087 ;
    wire n2088 ;
    wire n2089 ;
    wire n2090 ;
    wire n2091 ;
    wire n2092 ;
    wire n2093 ;
    wire n2094 ;
    wire n2095 ;
    wire n2096 ;
    wire n2097 ;
    wire n2098 ;
    wire n2099 ;
    wire n2100 ;
    wire n2101 ;
    wire n2102 ;
    wire n2103 ;
    wire n2104 ;
    wire n2105 ;
    wire n2106 ;
    wire n2107 ;
    wire n2108 ;
    wire n2109 ;
    wire n2110 ;
    wire n2111 ;
    wire n2112 ;
    wire n2113 ;
    wire n2114 ;
    wire n2115 ;
    wire n2116 ;
    wire n2117 ;
    wire n2118 ;
    wire n2119 ;
    wire n2120 ;
    wire n2121 ;
    wire n2122 ;
    wire n2123 ;
    wire n2124 ;
    wire n2125 ;
    wire n2126 ;
    wire n2127 ;
    wire n2128 ;
    wire n2129 ;
    wire n2130 ;
    wire n2131 ;
    wire n2132 ;
    wire n2133 ;
    wire n2134 ;
    wire n2135 ;
    wire n2136 ;
    wire n2137 ;
    wire n2138 ;
    wire n2139 ;
    wire n2140 ;
    wire n2141 ;
    wire n2142 ;
    wire n2143 ;
    wire n2144 ;
    wire n2145 ;
    wire n2146 ;
    wire n2147 ;
    wire n2148 ;
    wire n2149 ;
    wire n2150 ;
    wire n2151 ;
    wire n2152 ;
    wire n2153 ;
    wire n2154 ;
    wire n2155 ;
    wire n2156 ;
    wire n2157 ;
    wire n2158 ;
    wire n2159 ;
    wire n2160 ;
    wire n2161 ;
    wire n2162 ;
    wire n2163 ;
    wire n2164 ;
    wire n2165 ;
    wire n2166 ;
    wire n2167 ;
    wire n2168 ;
    wire n2169 ;
    wire n2170 ;
    wire n2171 ;
    wire n2172 ;
    wire n2173 ;
    wire n2174 ;
    wire n2175 ;
    wire n2176 ;
    wire n2177 ;
    wire n2178 ;
    wire n2179 ;
    wire n2180 ;
    wire n2181 ;
    wire n2182 ;
    wire n2183 ;
    wire n2184 ;
    wire n2185 ;
    wire n2186 ;
    wire n2187 ;
    wire n2188 ;
    wire n2189 ;
    wire n2190 ;
    wire n2191 ;
    wire n2192 ;
    wire n2193 ;
    wire n2194 ;
    wire n2195 ;
    wire n2196 ;
    wire n2197 ;
    wire n2198 ;
    wire n2199 ;
    wire n2200 ;
    wire n2201 ;
    wire n2202 ;
    wire n2203 ;
    wire n2204 ;
    wire n2205 ;
    wire n2206 ;
    wire n2207 ;
    wire n2208 ;
    wire n2209 ;
    wire n2210 ;
    wire n2211 ;
    wire n2212 ;
    wire n2213 ;
    wire n2214 ;
    wire n2215 ;
    wire n2216 ;
    wire n2217 ;
    wire n2218 ;
    wire n2219 ;
    wire n2220 ;
    wire n2221 ;
    wire n2222 ;
    wire n2223 ;
    wire n2224 ;
    wire n2225 ;
    wire n2226 ;
    wire n2227 ;
    wire n2228 ;
    wire n2229 ;
    wire n2230 ;
    wire n2231 ;
    wire n2232 ;
    wire n2233 ;
    wire n2234 ;
    wire n2235 ;
    wire n2236 ;
    wire n2237 ;
    wire n2238 ;
    wire n2239 ;
    wire n2240 ;
    wire n2241 ;
    wire n2242 ;
    wire n2243 ;
    wire n2244 ;
    wire n2245 ;
    wire n2246 ;
    wire n2247 ;
    wire n2248 ;
    wire n2249 ;
    wire n2250 ;
    wire n2251 ;
    wire n2252 ;
    wire n2253 ;
    wire n2254 ;
    wire n2255 ;
    wire n2256 ;
    wire n2257 ;
    wire n2258 ;
    wire n2259 ;
    wire n2260 ;
    wire n2261 ;
    wire n2262 ;
    wire n2263 ;
    wire n2264 ;
    wire n2265 ;
    wire n2266 ;
    wire n2267 ;
    wire n2268 ;
    wire n2269 ;
    wire n2270 ;
    wire n2271 ;
    wire n2272 ;
    wire n2273 ;
    wire n2274 ;
    wire n2275 ;
    wire n2276 ;
    wire n2277 ;
    wire n2278 ;
    wire n2279 ;
    wire n2280 ;
    wire n2281 ;
    wire n2282 ;
    wire n2283 ;
    wire n2284 ;
    wire n2285 ;
    wire n2286 ;
    wire n2287 ;
    wire n2288 ;
    wire n2289 ;
    wire n2290 ;
    wire n2291 ;
    wire n2292 ;
    wire n2293 ;
    wire n2294 ;
    wire n2295 ;
    wire n2296 ;
    wire n2297 ;
    wire n2298 ;
    wire n2299 ;
    wire n2300 ;
    wire n2301 ;
    wire n2302 ;
    wire n2303 ;
    wire n2304 ;
    wire n2305 ;
    wire n2306 ;
    wire n2307 ;
    wire n2308 ;
    wire n2309 ;
    wire n2310 ;
    wire n2311 ;
    wire n2312 ;
    wire n2313 ;
    wire n2314 ;
    wire n2315 ;
    wire n2316 ;
    wire n2317 ;
    wire n2318 ;
    wire n2319 ;
    wire n2320 ;
    wire n2321 ;
    wire n2322 ;
    wire n2323 ;
    wire n2324 ;
    wire n2325 ;
    wire n2326 ;
    wire n2327 ;
    wire n2328 ;
    wire n2329 ;
    wire n2330 ;
    wire n2331 ;
    wire n2332 ;
    wire n2333 ;
    wire n2334 ;
    wire n2335 ;
    wire n2336 ;
    wire n2337 ;
    wire n2338 ;
    wire n2339 ;
    wire n2340 ;
    wire n2341 ;
    wire n2342 ;
    wire n2343 ;
    wire n2344 ;
    wire n2345 ;
    wire n2346 ;
    wire n2347 ;
    wire n2348 ;
    wire n2349 ;
    wire n2350 ;
    wire n2351 ;
    wire n2352 ;
    wire n2353 ;
    wire n2354 ;
    wire n2355 ;
    wire n2356 ;
    wire n2357 ;
    wire n2358 ;
    wire n2359 ;
    wire n2360 ;
    wire n2361 ;
    wire n2362 ;
    wire n2363 ;
    wire n2364 ;
    wire n2365 ;
    wire n2366 ;
    wire n2367 ;
    wire n2368 ;
    wire n2369 ;
    wire n2370 ;
    wire n2371 ;
    wire n2372 ;
    wire n2373 ;
    wire n2374 ;
    wire n2375 ;
    wire n2376 ;
    wire n2377 ;
    wire n2378 ;
    wire n2379 ;
    wire n2380 ;
    wire n2381 ;
    wire n2382 ;
    wire n2383 ;
    wire n2384 ;
    wire n2385 ;
    wire n2386 ;
    wire n2387 ;
    wire n2388 ;
    wire n2389 ;
    wire n2390 ;
    wire n2391 ;
    wire n2392 ;
    wire n2393 ;
    wire n2394 ;
    wire n2395 ;
    wire n2396 ;
    wire n2397 ;
    wire n2398 ;
    wire n2399 ;
    wire n2400 ;
    wire n2401 ;
    wire n2402 ;
    wire n2403 ;
    wire n2404 ;
    wire n2405 ;
    wire n2406 ;
    wire n2407 ;
    wire n2408 ;
    wire n2409 ;
    wire n2410 ;
    wire n2411 ;
    wire n2412 ;
    wire n2413 ;
    wire n2414 ;
    wire n2415 ;
    wire n2416 ;
    wire n2417 ;
    wire n2418 ;
    wire n2419 ;
    wire n2420 ;
    wire n2421 ;
    wire n2422 ;
    wire n2423 ;
    wire n2424 ;
    wire n2425 ;
    wire n2426 ;
    wire n2427 ;
    wire n2428 ;
    wire n2429 ;
    wire n2430 ;
    wire n2431 ;
    wire n2432 ;
    wire n2433 ;
    wire n2434 ;
    wire n2435 ;
    wire n2436 ;
    wire n2437 ;
    wire n2438 ;
    wire n2439 ;
    wire n2440 ;
    wire n2441 ;
    wire n2442 ;
    wire n2443 ;
    wire n2444 ;
    wire n2445 ;
    wire n2446 ;
    wire n2447 ;
    wire n2448 ;
    wire n2449 ;
    wire n2450 ;
    wire n2451 ;
    wire n2452 ;
    wire n2453 ;
    wire n2454 ;
    wire n2455 ;
    wire n2456 ;
    wire n2457 ;
    wire n2458 ;
    wire n2459 ;
    wire n2460 ;
    wire n2461 ;
    wire n2462 ;
    wire n2463 ;
    wire n2464 ;
    wire n2465 ;
    wire n2466 ;
    wire n2467 ;
    wire n2468 ;
    wire n2469 ;
    wire n2470 ;
    wire n2471 ;
    wire n2472 ;
    wire n2473 ;
    wire n2474 ;
    wire n2475 ;
    wire n2476 ;
    wire n2477 ;
    wire n2478 ;
    wire n2479 ;
    wire n2480 ;
    wire n2481 ;
    wire n2482 ;
    wire n2483 ;
    wire n2484 ;
    wire n2485 ;
    wire n2486 ;
    wire n2487 ;
    wire n2488 ;
    wire n2489 ;
    wire n2490 ;
    wire n2491 ;
    wire n2492 ;
    wire n2493 ;
    wire n2494 ;
    wire n2495 ;
    wire n2496 ;
    wire n2497 ;
    wire n2498 ;
    wire n2499 ;
    wire n2500 ;
    wire n2501 ;
    wire n2502 ;
    wire n2503 ;
    wire n2504 ;
    wire n2505 ;
    wire n2506 ;
    wire n2507 ;
    wire n2508 ;
    wire n2509 ;
    wire n2510 ;
    wire n2511 ;
    wire n2512 ;
    wire n2513 ;
    wire n2514 ;
    wire n2515 ;
    wire n2516 ;
    wire n2517 ;
    wire n2518 ;
    wire n2519 ;
    wire n2520 ;
    wire n2521 ;
    wire n2522 ;
    wire n2523 ;
    wire n2524 ;
    wire n2525 ;
    wire n2526 ;
    wire n2527 ;
    wire n2528 ;
    wire n2529 ;
    wire n2530 ;
    wire n2531 ;
    wire n2532 ;
    wire n2533 ;
    wire n2534 ;
    wire n2535 ;
    wire n2536 ;
    wire n2537 ;
    wire n2538 ;
    wire n2539 ;
    wire n2540 ;
    wire n2541 ;
    wire n2542 ;
    wire n2543 ;
    wire n2544 ;
    wire n2545 ;
    wire n2546 ;
    wire n2547 ;
    wire n2548 ;
    wire n2549 ;
    wire n2550 ;
    wire n2551 ;
    wire n2552 ;
    wire n2553 ;
    wire n2554 ;
    wire n2555 ;
    wire n2556 ;
    wire n2557 ;
    wire n2558 ;
    wire n2559 ;
    wire n2560 ;
    wire n2561 ;
    wire n2562 ;
    wire n2563 ;
    wire n2564 ;
    wire n2565 ;
    wire n2566 ;
    wire n2567 ;
    wire n2568 ;
    wire n2569 ;
    wire n2570 ;
    wire n2571 ;
    wire n2572 ;
    wire n2573 ;
    wire n2574 ;
    wire n2575 ;
    wire n2576 ;
    wire n2577 ;
    wire n2578 ;
    wire n2579 ;
    wire n2580 ;
    wire n2581 ;
    wire n2582 ;
    wire n2583 ;
    wire n2584 ;
    wire n2585 ;
    wire n2586 ;
    wire n2587 ;
    wire n2588 ;
    wire n2589 ;
    wire n2590 ;
    wire n2591 ;
    wire n2592 ;
    wire n2593 ;
    wire n2594 ;
    wire n2595 ;
    wire n2596 ;
    wire n2597 ;
    wire n2598 ;
    wire n2599 ;
    wire n2600 ;
    wire n2601 ;
    wire n2602 ;
    wire n2603 ;
    wire n2604 ;
    wire n2605 ;
    wire n2606 ;
    wire n2607 ;
    wire n2608 ;
    wire n2609 ;
    wire n2610 ;
    wire n2611 ;
    wire n2612 ;
    wire n2613 ;
    wire n2614 ;
    wire n2615 ;
    wire n2616 ;
    wire n2617 ;
    wire n2618 ;
    wire n2619 ;
    wire n2620 ;
    wire n2621 ;
    wire n2622 ;
    wire n2623 ;
    wire n2624 ;
    wire n2625 ;
    wire n2626 ;
    wire n2627 ;
    wire n2628 ;
    wire n2629 ;
    wire n2630 ;
    wire n2631 ;
    wire n2632 ;
    wire n2633 ;
    wire n2634 ;
    wire n2635 ;
    wire n2636 ;
    wire n2637 ;
    wire n2638 ;
    wire n2639 ;
    wire n2640 ;
    wire n2641 ;
    wire n2642 ;
    wire n2643 ;
    wire n2644 ;
    wire n2645 ;
    wire n2646 ;
    wire n2647 ;
    wire n2648 ;
    wire n2649 ;
    wire n2650 ;
    wire n2651 ;
    wire n2652 ;
    wire n2653 ;
    wire n2654 ;
    wire n2655 ;
    wire n2656 ;
    wire n2657 ;
    wire n2658 ;
    wire n2659 ;
    wire n2660 ;
    wire n2661 ;
    wire n2662 ;
    wire n2663 ;
    wire n2664 ;
    wire n2665 ;
    wire n2666 ;
    wire n2667 ;
    wire n2668 ;
    wire n2669 ;
    wire n2670 ;
    wire n2671 ;
    wire n2672 ;
    wire n2673 ;
    wire n2674 ;
    wire n2675 ;
    wire n2676 ;
    wire n2677 ;
    wire n2678 ;
    wire n2679 ;
    wire n2680 ;
    wire n2681 ;
    wire n2682 ;
    wire n2683 ;
    wire n2684 ;
    wire n2685 ;
    wire n2686 ;
    wire n2687 ;
    wire n2688 ;
    wire n2689 ;
    wire n2690 ;
    wire n2691 ;
    wire n2692 ;
    wire n2693 ;
    wire n2694 ;
    wire n2695 ;
    wire n2696 ;
    wire n2697 ;
    wire n2698 ;
    wire n2699 ;
    wire n2700 ;
    wire n2701 ;
    wire n2702 ;
    wire n2703 ;
    wire n2704 ;
    wire n2705 ;
    wire n2706 ;
    wire n2707 ;
    wire n2708 ;
    wire n2709 ;
    wire n2710 ;
    wire n2711 ;
    wire n2712 ;
    wire n2713 ;
    wire n2714 ;
    wire n2715 ;
    wire n2716 ;
    wire n2717 ;
    wire n2718 ;
    wire n2719 ;
    wire n2720 ;
    wire n2721 ;
    wire n2722 ;
    wire n2723 ;
    wire n2724 ;
    wire n2725 ;
    wire n2726 ;
    wire n2727 ;
    wire n2728 ;
    wire n2729 ;
    wire n2730 ;
    wire n2731 ;
    wire n2732 ;
    wire n2733 ;
    wire n2734 ;
    wire n2735 ;
    wire n2736 ;
    wire n2737 ;
    wire n2738 ;
    wire n2739 ;
    wire n2740 ;
    wire n2741 ;
    wire n2742 ;
    wire n2743 ;
    wire n2744 ;
    wire n2745 ;
    wire n2746 ;
    wire n2747 ;
    wire n2748 ;
    wire n2749 ;
    wire n2750 ;
    wire n2751 ;
    wire n2752 ;
    wire n2753 ;
    wire n2754 ;
    wire n2755 ;
    wire n2756 ;
    wire n2757 ;
    wire n2758 ;
    wire n2759 ;
    wire n2760 ;
    wire n2761 ;
    wire n2762 ;
    wire n2763 ;
    wire n2764 ;
    wire n2765 ;
    wire n2766 ;
    wire n2767 ;
    wire n2768 ;
    wire n2769 ;
    wire n2770 ;
    wire n2771 ;
    wire n2772 ;
    wire n2773 ;
    wire n2774 ;
    wire n2775 ;
    wire n2776 ;
    wire n2777 ;
    wire n2778 ;
    wire n2779 ;
    wire n2780 ;
    wire n2781 ;
    wire n2782 ;
    wire n2783 ;
    wire n2784 ;
    wire n2785 ;
    wire n2786 ;
    wire n2787 ;
    wire n2788 ;
    wire n2789 ;
    wire n2790 ;
    wire n2791 ;
    wire n2792 ;
    wire n2793 ;
    wire n2794 ;
    wire n2795 ;
    wire n2796 ;
    wire n2797 ;
    wire n2798 ;
    wire n2799 ;
    wire n2800 ;
    wire n2801 ;
    wire n2802 ;
    wire n2803 ;
    wire n2804 ;
    wire n2805 ;
    wire n2806 ;
    wire n2807 ;
    wire n2808 ;
    wire n2809 ;
    wire n2810 ;
    wire n2811 ;
    wire n2812 ;
    wire n2813 ;
    wire n2814 ;
    wire n2815 ;
    wire n2816 ;
    wire n2817 ;
    wire n2818 ;
    wire n2819 ;
    wire n2820 ;
    wire n2821 ;
    wire n2822 ;
    wire n2823 ;
    wire n2824 ;
    wire n2825 ;
    wire n2826 ;
    wire n2827 ;
    wire n2828 ;
    wire n2829 ;
    wire n2830 ;
    wire n2831 ;
    wire n2832 ;
    wire new_AGEMA_signal_943 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_947 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_951 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_955 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_958 ;
    wire new_AGEMA_signal_959 ;
    wire new_AGEMA_signal_960 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_962 ;
    wire new_AGEMA_signal_963 ;
    wire new_AGEMA_signal_964 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_966 ;
    wire new_AGEMA_signal_967 ;
    wire new_AGEMA_signal_968 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_970 ;
    wire new_AGEMA_signal_971 ;
    wire new_AGEMA_signal_972 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_974 ;
    wire new_AGEMA_signal_975 ;
    wire new_AGEMA_signal_976 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_978 ;
    wire new_AGEMA_signal_979 ;
    wire new_AGEMA_signal_980 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_982 ;
    wire new_AGEMA_signal_983 ;
    wire new_AGEMA_signal_984 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_986 ;
    wire new_AGEMA_signal_987 ;
    wire new_AGEMA_signal_988 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_990 ;
    wire new_AGEMA_signal_991 ;
    wire new_AGEMA_signal_992 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_994 ;
    wire new_AGEMA_signal_995 ;
    wire new_AGEMA_signal_996 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_998 ;
    wire new_AGEMA_signal_999 ;
    wire new_AGEMA_signal_1000 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1002 ;
    wire new_AGEMA_signal_1003 ;
    wire new_AGEMA_signal_1004 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1006 ;
    wire new_AGEMA_signal_1007 ;
    wire new_AGEMA_signal_1008 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1010 ;
    wire new_AGEMA_signal_1011 ;
    wire new_AGEMA_signal_1012 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1014 ;
    wire new_AGEMA_signal_1015 ;
    wire new_AGEMA_signal_1016 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1018 ;
    wire new_AGEMA_signal_1019 ;
    wire new_AGEMA_signal_1020 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1022 ;
    wire new_AGEMA_signal_1023 ;
    wire new_AGEMA_signal_1024 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1026 ;
    wire new_AGEMA_signal_1027 ;
    wire new_AGEMA_signal_1028 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1030 ;
    wire new_AGEMA_signal_1031 ;
    wire new_AGEMA_signal_1032 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1034 ;
    wire new_AGEMA_signal_1035 ;
    wire new_AGEMA_signal_1036 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1038 ;
    wire new_AGEMA_signal_1039 ;
    wire new_AGEMA_signal_1040 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1042 ;
    wire new_AGEMA_signal_1043 ;
    wire new_AGEMA_signal_1044 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1046 ;
    wire new_AGEMA_signal_1047 ;
    wire new_AGEMA_signal_1048 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1050 ;
    wire new_AGEMA_signal_1051 ;
    wire new_AGEMA_signal_1052 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1054 ;
    wire new_AGEMA_signal_1055 ;
    wire new_AGEMA_signal_1056 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1058 ;
    wire new_AGEMA_signal_1059 ;
    wire new_AGEMA_signal_1060 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1062 ;
    wire new_AGEMA_signal_1063 ;
    wire new_AGEMA_signal_1064 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1066 ;
    wire new_AGEMA_signal_1067 ;
    wire new_AGEMA_signal_1068 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1070 ;
    wire new_AGEMA_signal_1071 ;
    wire new_AGEMA_signal_1072 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1074 ;
    wire new_AGEMA_signal_1075 ;
    wire new_AGEMA_signal_1076 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1078 ;
    wire new_AGEMA_signal_1079 ;
    wire new_AGEMA_signal_1080 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1082 ;
    wire new_AGEMA_signal_1083 ;
    wire new_AGEMA_signal_1084 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1086 ;
    wire new_AGEMA_signal_1087 ;
    wire new_AGEMA_signal_1088 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1090 ;
    wire new_AGEMA_signal_1091 ;
    wire new_AGEMA_signal_1092 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1094 ;
    wire new_AGEMA_signal_1095 ;
    wire new_AGEMA_signal_1096 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1098 ;
    wire new_AGEMA_signal_1099 ;
    wire new_AGEMA_signal_1100 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1102 ;
    wire new_AGEMA_signal_1103 ;
    wire new_AGEMA_signal_1104 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1106 ;
    wire new_AGEMA_signal_1107 ;
    wire new_AGEMA_signal_1108 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1110 ;
    wire new_AGEMA_signal_1111 ;
    wire new_AGEMA_signal_1112 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1114 ;
    wire new_AGEMA_signal_1115 ;
    wire new_AGEMA_signal_1116 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1264 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1266 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1268 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1270 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1272 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1274 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1276 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1278 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1280 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1282 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1284 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1286 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1288 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1290 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1292 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1294 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1344 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1346 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1348 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1350 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1352 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1354 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1356 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1358 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1360 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1362 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1364 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1366 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1368 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1370 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1372 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1374 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1376 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1378 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1380 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1382 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1384 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1386 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1388 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1390 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1392 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1394 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1396 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1398 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1400 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1402 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1404 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1406 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1408 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1410 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1412 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1414 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1416 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1418 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1420 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1422 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1424 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1426 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1428 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1430 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1432 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1434 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1436 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1438 ;
    wire new_AGEMA_signal_1439 ;
    wire new_AGEMA_signal_1440 ;
    wire new_AGEMA_signal_1441 ;
    wire new_AGEMA_signal_1442 ;
    wire new_AGEMA_signal_1443 ;
    wire new_AGEMA_signal_1444 ;
    wire new_AGEMA_signal_1445 ;
    wire new_AGEMA_signal_1446 ;
    wire new_AGEMA_signal_1447 ;
    wire new_AGEMA_signal_1448 ;
    wire new_AGEMA_signal_1449 ;
    wire new_AGEMA_signal_1450 ;
    wire new_AGEMA_signal_1451 ;
    wire new_AGEMA_signal_1452 ;
    wire new_AGEMA_signal_1453 ;
    wire new_AGEMA_signal_1454 ;
    wire new_AGEMA_signal_1455 ;
    wire new_AGEMA_signal_1456 ;
    wire new_AGEMA_signal_1457 ;
    wire new_AGEMA_signal_1458 ;
    wire new_AGEMA_signal_1459 ;
    wire new_AGEMA_signal_1460 ;
    wire new_AGEMA_signal_1461 ;
    wire new_AGEMA_signal_1462 ;
    wire new_AGEMA_signal_1463 ;
    wire new_AGEMA_signal_1464 ;
    wire new_AGEMA_signal_1465 ;
    wire new_AGEMA_signal_1466 ;
    wire new_AGEMA_signal_1467 ;
    wire new_AGEMA_signal_1468 ;
    wire new_AGEMA_signal_1469 ;
    wire new_AGEMA_signal_1470 ;
    wire new_AGEMA_signal_1471 ;
    wire new_AGEMA_signal_1472 ;
    wire new_AGEMA_signal_1473 ;
    wire new_AGEMA_signal_1474 ;
    wire new_AGEMA_signal_1475 ;
    wire new_AGEMA_signal_1476 ;
    wire new_AGEMA_signal_1477 ;
    wire new_AGEMA_signal_1478 ;
    wire new_AGEMA_signal_1479 ;
    wire new_AGEMA_signal_1480 ;
    wire new_AGEMA_signal_1481 ;
    wire new_AGEMA_signal_1482 ;
    wire new_AGEMA_signal_1483 ;
    wire new_AGEMA_signal_1484 ;
    wire new_AGEMA_signal_1485 ;
    wire new_AGEMA_signal_1486 ;
    wire new_AGEMA_signal_1487 ;
    wire new_AGEMA_signal_1488 ;
    wire new_AGEMA_signal_1489 ;
    wire new_AGEMA_signal_1490 ;
    wire new_AGEMA_signal_1491 ;
    wire new_AGEMA_signal_1492 ;
    wire new_AGEMA_signal_1493 ;
    wire new_AGEMA_signal_1494 ;
    wire new_AGEMA_signal_1495 ;
    wire new_AGEMA_signal_1496 ;
    wire new_AGEMA_signal_1497 ;
    wire new_AGEMA_signal_1498 ;
    wire new_AGEMA_signal_1499 ;
    wire new_AGEMA_signal_1500 ;
    wire new_AGEMA_signal_1501 ;
    wire new_AGEMA_signal_1502 ;
    wire new_AGEMA_signal_1503 ;
    wire new_AGEMA_signal_1504 ;
    wire new_AGEMA_signal_1505 ;
    wire new_AGEMA_signal_1506 ;
    wire new_AGEMA_signal_1507 ;
    wire new_AGEMA_signal_1508 ;
    wire new_AGEMA_signal_1509 ;
    wire new_AGEMA_signal_1510 ;
    wire new_AGEMA_signal_1511 ;
    wire new_AGEMA_signal_1512 ;
    wire new_AGEMA_signal_1513 ;
    wire new_AGEMA_signal_1514 ;
    wire new_AGEMA_signal_1515 ;
    wire new_AGEMA_signal_1516 ;
    wire new_AGEMA_signal_1517 ;
    wire new_AGEMA_signal_1518 ;
    wire new_AGEMA_signal_1519 ;
    wire new_AGEMA_signal_1520 ;
    wire new_AGEMA_signal_1521 ;
    wire new_AGEMA_signal_1522 ;
    wire new_AGEMA_signal_1523 ;
    wire new_AGEMA_signal_1524 ;
    wire new_AGEMA_signal_1525 ;
    wire new_AGEMA_signal_1526 ;
    wire new_AGEMA_signal_1527 ;
    wire new_AGEMA_signal_1528 ;
    wire new_AGEMA_signal_1529 ;
    wire new_AGEMA_signal_1530 ;
    wire new_AGEMA_signal_1531 ;
    wire new_AGEMA_signal_1532 ;
    wire new_AGEMA_signal_1533 ;
    wire new_AGEMA_signal_1534 ;
    wire new_AGEMA_signal_1535 ;
    wire new_AGEMA_signal_1536 ;
    wire new_AGEMA_signal_1537 ;
    wire new_AGEMA_signal_1538 ;
    wire new_AGEMA_signal_1539 ;
    wire new_AGEMA_signal_1540 ;
    wire new_AGEMA_signal_1541 ;
    wire new_AGEMA_signal_1542 ;
    wire new_AGEMA_signal_1543 ;
    wire new_AGEMA_signal_1544 ;
    wire new_AGEMA_signal_1545 ;
    wire new_AGEMA_signal_1546 ;
    wire new_AGEMA_signal_1547 ;
    wire new_AGEMA_signal_1548 ;
    wire new_AGEMA_signal_1549 ;
    wire new_AGEMA_signal_1550 ;
    wire new_AGEMA_signal_1551 ;
    wire new_AGEMA_signal_1552 ;
    wire new_AGEMA_signal_1553 ;
    wire new_AGEMA_signal_1554 ;
    wire new_AGEMA_signal_1555 ;
    wire new_AGEMA_signal_1556 ;
    wire new_AGEMA_signal_1557 ;
    wire new_AGEMA_signal_1558 ;
    wire new_AGEMA_signal_1559 ;
    wire new_AGEMA_signal_1560 ;
    wire new_AGEMA_signal_1561 ;
    wire new_AGEMA_signal_1562 ;
    wire new_AGEMA_signal_1563 ;
    wire new_AGEMA_signal_1564 ;
    wire new_AGEMA_signal_1565 ;
    wire new_AGEMA_signal_1566 ;
    wire new_AGEMA_signal_1567 ;
    wire new_AGEMA_signal_1568 ;
    wire new_AGEMA_signal_1569 ;
    wire new_AGEMA_signal_1570 ;
    wire new_AGEMA_signal_1571 ;
    wire new_AGEMA_signal_1572 ;
    wire new_AGEMA_signal_1573 ;
    wire new_AGEMA_signal_1574 ;
    wire new_AGEMA_signal_1575 ;
    wire new_AGEMA_signal_1576 ;
    wire new_AGEMA_signal_1577 ;
    wire new_AGEMA_signal_1578 ;
    wire new_AGEMA_signal_1579 ;
    wire new_AGEMA_signal_1580 ;
    wire new_AGEMA_signal_1581 ;
    wire new_AGEMA_signal_1582 ;
    wire new_AGEMA_signal_1583 ;
    wire new_AGEMA_signal_1584 ;
    wire new_AGEMA_signal_1585 ;
    wire new_AGEMA_signal_1586 ;
    wire new_AGEMA_signal_1587 ;
    wire new_AGEMA_signal_1588 ;
    wire new_AGEMA_signal_1589 ;
    wire new_AGEMA_signal_1590 ;
    wire new_AGEMA_signal_1591 ;
    wire new_AGEMA_signal_1592 ;
    wire new_AGEMA_signal_1593 ;
    wire new_AGEMA_signal_1594 ;
    wire new_AGEMA_signal_1595 ;
    wire new_AGEMA_signal_1596 ;
    wire new_AGEMA_signal_1597 ;
    wire new_AGEMA_signal_1598 ;
    wire new_AGEMA_signal_1599 ;
    wire new_AGEMA_signal_1600 ;
    wire new_AGEMA_signal_1601 ;
    wire new_AGEMA_signal_1602 ;
    wire new_AGEMA_signal_1603 ;
    wire new_AGEMA_signal_1604 ;
    wire new_AGEMA_signal_1605 ;
    wire new_AGEMA_signal_1606 ;
    wire new_AGEMA_signal_1607 ;
    wire new_AGEMA_signal_1608 ;
    wire new_AGEMA_signal_1609 ;
    wire new_AGEMA_signal_1610 ;
    wire new_AGEMA_signal_1611 ;
    wire new_AGEMA_signal_1612 ;
    wire new_AGEMA_signal_1613 ;
    wire new_AGEMA_signal_1614 ;
    wire new_AGEMA_signal_1615 ;
    wire new_AGEMA_signal_1616 ;
    wire new_AGEMA_signal_1617 ;
    wire new_AGEMA_signal_1618 ;
    wire new_AGEMA_signal_1619 ;
    wire new_AGEMA_signal_1620 ;
    wire new_AGEMA_signal_1621 ;
    wire new_AGEMA_signal_1622 ;
    wire new_AGEMA_signal_1623 ;
    wire new_AGEMA_signal_1624 ;
    wire new_AGEMA_signal_1625 ;
    wire new_AGEMA_signal_1626 ;
    wire new_AGEMA_signal_1627 ;
    wire new_AGEMA_signal_1628 ;
    wire new_AGEMA_signal_1629 ;
    wire new_AGEMA_signal_1630 ;
    wire new_AGEMA_signal_1631 ;
    wire new_AGEMA_signal_1632 ;
    wire new_AGEMA_signal_1633 ;
    wire new_AGEMA_signal_1634 ;
    wire new_AGEMA_signal_1635 ;
    wire new_AGEMA_signal_1636 ;
    wire new_AGEMA_signal_1637 ;
    wire new_AGEMA_signal_1638 ;
    wire new_AGEMA_signal_1639 ;
    wire new_AGEMA_signal_1640 ;
    wire new_AGEMA_signal_1641 ;
    wire new_AGEMA_signal_1642 ;
    wire new_AGEMA_signal_1643 ;
    wire new_AGEMA_signal_1644 ;
    wire new_AGEMA_signal_1645 ;
    wire new_AGEMA_signal_1646 ;
    wire new_AGEMA_signal_1647 ;
    wire new_AGEMA_signal_1648 ;
    wire new_AGEMA_signal_1649 ;
    wire new_AGEMA_signal_1650 ;
    wire new_AGEMA_signal_1651 ;
    wire new_AGEMA_signal_1652 ;
    wire new_AGEMA_signal_1653 ;
    wire new_AGEMA_signal_1654 ;
    wire new_AGEMA_signal_1655 ;
    wire new_AGEMA_signal_1656 ;
    wire new_AGEMA_signal_1657 ;
    wire new_AGEMA_signal_1658 ;
    wire new_AGEMA_signal_1659 ;
    wire new_AGEMA_signal_1660 ;
    wire new_AGEMA_signal_1661 ;
    wire new_AGEMA_signal_1662 ;
    wire new_AGEMA_signal_1663 ;
    wire new_AGEMA_signal_1664 ;
    wire new_AGEMA_signal_1665 ;
    wire new_AGEMA_signal_1666 ;
    wire new_AGEMA_signal_1667 ;
    wire new_AGEMA_signal_1668 ;
    wire new_AGEMA_signal_1669 ;
    wire new_AGEMA_signal_1670 ;
    wire new_AGEMA_signal_1671 ;
    wire new_AGEMA_signal_1672 ;
    wire new_AGEMA_signal_1673 ;
    wire new_AGEMA_signal_1674 ;
    wire new_AGEMA_signal_1675 ;
    wire new_AGEMA_signal_1676 ;
    wire new_AGEMA_signal_1677 ;
    wire new_AGEMA_signal_1678 ;
    wire new_AGEMA_signal_1679 ;
    wire new_AGEMA_signal_1680 ;
    wire new_AGEMA_signal_1681 ;
    wire new_AGEMA_signal_1682 ;
    wire new_AGEMA_signal_1683 ;
    wire new_AGEMA_signal_1684 ;
    wire new_AGEMA_signal_1685 ;
    wire new_AGEMA_signal_1686 ;
    wire new_AGEMA_signal_1687 ;
    wire new_AGEMA_signal_1688 ;
    wire new_AGEMA_signal_1689 ;
    wire new_AGEMA_signal_1690 ;
    wire new_AGEMA_signal_1691 ;
    wire new_AGEMA_signal_1692 ;
    wire new_AGEMA_signal_1693 ;
    wire new_AGEMA_signal_1694 ;
    wire new_AGEMA_signal_1695 ;
    wire new_AGEMA_signal_1696 ;
    wire new_AGEMA_signal_1697 ;
    wire new_AGEMA_signal_1698 ;
    wire new_AGEMA_signal_1699 ;
    wire new_AGEMA_signal_1700 ;
    wire new_AGEMA_signal_1701 ;
    wire new_AGEMA_signal_1702 ;
    wire new_AGEMA_signal_1703 ;
    wire new_AGEMA_signal_1704 ;
    wire new_AGEMA_signal_1705 ;
    wire new_AGEMA_signal_1706 ;
    wire new_AGEMA_signal_1707 ;
    wire new_AGEMA_signal_1708 ;
    wire new_AGEMA_signal_1709 ;
    wire new_AGEMA_signal_1710 ;
    wire new_AGEMA_signal_1711 ;
    wire new_AGEMA_signal_1712 ;
    wire new_AGEMA_signal_1713 ;
    wire new_AGEMA_signal_1714 ;
    wire new_AGEMA_signal_1715 ;
    wire new_AGEMA_signal_1716 ;
    wire new_AGEMA_signal_1717 ;
    wire new_AGEMA_signal_1718 ;
    wire new_AGEMA_signal_1719 ;
    wire new_AGEMA_signal_1720 ;
    wire new_AGEMA_signal_1721 ;
    wire new_AGEMA_signal_1722 ;
    wire new_AGEMA_signal_1723 ;
    wire new_AGEMA_signal_1724 ;
    wire new_AGEMA_signal_1725 ;
    wire new_AGEMA_signal_1726 ;
    wire new_AGEMA_signal_1727 ;
    wire new_AGEMA_signal_1728 ;
    wire new_AGEMA_signal_1729 ;
    wire new_AGEMA_signal_1730 ;
    wire new_AGEMA_signal_1731 ;
    wire new_AGEMA_signal_1732 ;
    wire new_AGEMA_signal_1733 ;
    wire new_AGEMA_signal_1734 ;
    wire new_AGEMA_signal_1735 ;
    wire new_AGEMA_signal_1736 ;
    wire new_AGEMA_signal_1737 ;
    wire new_AGEMA_signal_1738 ;
    wire new_AGEMA_signal_1739 ;
    wire new_AGEMA_signal_1740 ;
    wire new_AGEMA_signal_1741 ;
    wire new_AGEMA_signal_1742 ;
    wire new_AGEMA_signal_1743 ;
    wire new_AGEMA_signal_1744 ;
    wire new_AGEMA_signal_1745 ;
    wire new_AGEMA_signal_1746 ;
    wire new_AGEMA_signal_1747 ;
    wire new_AGEMA_signal_1748 ;
    wire new_AGEMA_signal_1749 ;
    wire new_AGEMA_signal_1750 ;
    wire new_AGEMA_signal_1751 ;
    wire new_AGEMA_signal_1752 ;
    wire new_AGEMA_signal_1753 ;
    wire new_AGEMA_signal_1754 ;
    wire new_AGEMA_signal_1755 ;
    wire new_AGEMA_signal_1756 ;
    wire new_AGEMA_signal_1757 ;
    wire new_AGEMA_signal_1758 ;
    wire new_AGEMA_signal_1759 ;
    wire new_AGEMA_signal_1760 ;
    wire new_AGEMA_signal_1761 ;
    wire new_AGEMA_signal_1762 ;
    wire new_AGEMA_signal_1763 ;
    wire new_AGEMA_signal_1764 ;
    wire new_AGEMA_signal_1765 ;
    wire new_AGEMA_signal_1766 ;
    wire new_AGEMA_signal_1767 ;
    wire new_AGEMA_signal_1768 ;
    wire new_AGEMA_signal_1769 ;
    wire new_AGEMA_signal_1770 ;
    wire new_AGEMA_signal_1771 ;
    wire new_AGEMA_signal_1772 ;
    wire new_AGEMA_signal_1773 ;
    wire new_AGEMA_signal_1774 ;
    wire new_AGEMA_signal_1775 ;
    wire new_AGEMA_signal_1776 ;
    wire new_AGEMA_signal_1777 ;
    wire new_AGEMA_signal_1778 ;
    wire new_AGEMA_signal_1779 ;
    wire new_AGEMA_signal_1780 ;
    wire new_AGEMA_signal_1781 ;
    wire new_AGEMA_signal_1782 ;
    wire new_AGEMA_signal_1783 ;
    wire new_AGEMA_signal_1784 ;
    wire new_AGEMA_signal_1785 ;
    wire new_AGEMA_signal_1786 ;
    wire new_AGEMA_signal_1787 ;
    wire new_AGEMA_signal_1788 ;
    wire new_AGEMA_signal_1789 ;
    wire new_AGEMA_signal_1790 ;
    wire new_AGEMA_signal_1791 ;
    wire new_AGEMA_signal_1792 ;
    wire new_AGEMA_signal_1793 ;
    wire new_AGEMA_signal_1794 ;
    wire new_AGEMA_signal_1795 ;
    wire new_AGEMA_signal_1796 ;
    wire new_AGEMA_signal_1797 ;
    wire new_AGEMA_signal_1798 ;
    wire new_AGEMA_signal_1799 ;
    wire new_AGEMA_signal_1800 ;
    wire new_AGEMA_signal_1801 ;
    wire new_AGEMA_signal_1802 ;
    wire new_AGEMA_signal_1803 ;
    wire new_AGEMA_signal_1804 ;
    wire new_AGEMA_signal_1805 ;
    wire new_AGEMA_signal_1806 ;
    wire new_AGEMA_signal_1807 ;
    wire new_AGEMA_signal_1808 ;
    wire new_AGEMA_signal_1809 ;
    wire new_AGEMA_signal_1810 ;
    wire new_AGEMA_signal_1811 ;
    wire new_AGEMA_signal_1812 ;
    wire new_AGEMA_signal_1813 ;
    wire new_AGEMA_signal_1814 ;
    wire new_AGEMA_signal_1815 ;
    wire new_AGEMA_signal_1816 ;
    wire new_AGEMA_signal_1817 ;
    wire new_AGEMA_signal_1818 ;
    wire new_AGEMA_signal_1819 ;
    wire new_AGEMA_signal_1820 ;
    wire new_AGEMA_signal_1821 ;
    wire new_AGEMA_signal_1822 ;
    wire new_AGEMA_signal_1823 ;
    wire new_AGEMA_signal_1824 ;
    wire new_AGEMA_signal_1825 ;
    wire new_AGEMA_signal_1826 ;
    wire new_AGEMA_signal_1827 ;
    wire new_AGEMA_signal_1828 ;
    wire new_AGEMA_signal_1829 ;
    wire new_AGEMA_signal_1830 ;
    wire new_AGEMA_signal_1831 ;
    wire new_AGEMA_signal_1832 ;
    wire new_AGEMA_signal_1833 ;
    wire new_AGEMA_signal_1834 ;
    wire new_AGEMA_signal_1835 ;
    wire new_AGEMA_signal_1836 ;
    wire new_AGEMA_signal_1837 ;
    wire new_AGEMA_signal_1838 ;
    wire new_AGEMA_signal_1839 ;
    wire new_AGEMA_signal_1840 ;
    wire new_AGEMA_signal_1841 ;
    wire new_AGEMA_signal_1842 ;
    wire new_AGEMA_signal_1843 ;
    wire new_AGEMA_signal_1844 ;
    wire new_AGEMA_signal_1845 ;
    wire new_AGEMA_signal_1846 ;
    wire new_AGEMA_signal_1847 ;
    wire new_AGEMA_signal_1848 ;
    wire new_AGEMA_signal_1849 ;
    wire new_AGEMA_signal_1850 ;
    wire new_AGEMA_signal_1851 ;
    wire new_AGEMA_signal_1852 ;
    wire new_AGEMA_signal_1853 ;
    wire new_AGEMA_signal_1854 ;
    wire new_AGEMA_signal_1855 ;
    wire new_AGEMA_signal_1856 ;
    wire new_AGEMA_signal_1857 ;
    wire new_AGEMA_signal_1858 ;
    wire new_AGEMA_signal_1859 ;
    wire new_AGEMA_signal_1860 ;
    wire new_AGEMA_signal_1861 ;
    wire new_AGEMA_signal_1862 ;
    wire new_AGEMA_signal_1863 ;
    wire new_AGEMA_signal_1864 ;
    wire new_AGEMA_signal_1865 ;
    wire new_AGEMA_signal_1866 ;
    wire new_AGEMA_signal_1867 ;
    wire new_AGEMA_signal_1868 ;
    wire clk_gated ;

    /* cells in depth 0 */
    not_masked #(.low_latency(0), .pipeline(0)) U1938 ( .a ({SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_943, n2796}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1939 ( .a ({SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_945, n2810}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1940 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_947, n2462}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1941 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_949, n2760}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1942 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_951, n2791}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1944 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_953, n2813}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1945 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_955, n2630}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1946 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_957, n2765}) ) ;
    ClockGatingController #(35) ClockGatingInst ( .clk ( clk ), .rst ( rst ), .GatedClk ( clk_gated ), .Synch ( Synch ) ) ;

    /* cells in depth 1 */

    /* cells in depth 2 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1937 ( .a ({new_AGEMA_signal_943, n2796}), .b ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ( Fresh[0] ), .c ({new_AGEMA_signal_970, n2719}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1943 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_1023, n2672}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1947 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[1] ), .c ({new_AGEMA_signal_958, n2635}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1948 ( .a ({new_AGEMA_signal_947, n2462}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ( Fresh[2] ), .c ({new_AGEMA_signal_971, n2641}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1949 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[3] ), .c ({new_AGEMA_signal_959, n2790}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1950 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ( Fresh[4] ), .c ({new_AGEMA_signal_960, n2519}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1951 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_972, n2750}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1952 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[5] ), .c ({new_AGEMA_signal_973, n2615}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1953 ( .a ({new_AGEMA_signal_973, n2615}), .b ({new_AGEMA_signal_1024, n2640}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1955 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[6] ), .c ({new_AGEMA_signal_974, n2699}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1956 ( .a ({new_AGEMA_signal_974, n2699}), .b ({new_AGEMA_signal_1025, n2737}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1957 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[7] ), .c ({new_AGEMA_signal_975, n2816}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1958 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_1026, n2767}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1961 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[8] ), .c ({new_AGEMA_signal_976, n2780}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1962 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1027, n2789}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1963 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_945, n2810}), .clk ( clk ), .r ( Fresh[9] ), .c ({new_AGEMA_signal_977, n2317}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1965 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[10] ), .c ({new_AGEMA_signal_978, n2694}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1966 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1028, n2769}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1969 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[11] ), .c ({new_AGEMA_signal_979, n2073}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1970 ( .a ({new_AGEMA_signal_979, n2073}), .b ({new_AGEMA_signal_1029, n2707}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1971 ( .a ({SI_s1[7], SI_s0[7]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[12] ), .c ({new_AGEMA_signal_961, n2315}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1972 ( .a ({SI_s1[0], SI_s0[0]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[13] ), .c ({new_AGEMA_signal_962, n2682}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1973 ( .a ({new_AGEMA_signal_962, n2682}), .b ({new_AGEMA_signal_980, n2713}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1975 ( .a ({new_AGEMA_signal_953, n2813}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[14] ), .c ({new_AGEMA_signal_981, n2723}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1976 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1031, n2688}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1978 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ( Fresh[15] ), .c ({new_AGEMA_signal_982, n2725}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1979 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1032, n2541}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1984 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[16] ), .c ({new_AGEMA_signal_983, n2815}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1985 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_1033, n2086}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1987 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[17] ), .c ({new_AGEMA_signal_984, n2600}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1990 ( .a ({new_AGEMA_signal_947, n2462}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[18] ), .c ({new_AGEMA_signal_985, n2538}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1991 ( .a ({new_AGEMA_signal_985, n2538}), .b ({new_AGEMA_signal_1035, n2786}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1995 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[19] ), .c ({new_AGEMA_signal_963, n2595}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1996 ( .a ({new_AGEMA_signal_963, n2595}), .b ({new_AGEMA_signal_986, n2742}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1999 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[20] ), .c ({new_AGEMA_signal_987, n2753}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2000 ( .a ({new_AGEMA_signal_987, n2753}), .b ({new_AGEMA_signal_1037, n2577}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2004 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[21] ), .c ({new_AGEMA_signal_988, n2400}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2008 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[22] ), .c ({new_AGEMA_signal_989, n2785}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2009 ( .a ({new_AGEMA_signal_989, n2785}), .b ({new_AGEMA_signal_1039, n2792}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2013 ( .a ({new_AGEMA_signal_953, n2813}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[23] ), .c ({new_AGEMA_signal_990, n2609}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2014 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_1040, n2724}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2017 ( .a ({new_AGEMA_signal_949, n2760}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[24] ), .c ({new_AGEMA_signal_991, n2661}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2018 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1041, n2174}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2020 ( .a ({SI_s1[2], SI_s0[2]}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[25] ), .c ({new_AGEMA_signal_964, n2708}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2021 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_992, n2493}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2025 ( .a ({new_AGEMA_signal_943, n2796}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[26] ), .c ({new_AGEMA_signal_993, n2587}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2028 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1044, n2570}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2029 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[27] ), .c ({new_AGEMA_signal_965, n2559}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2035 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[28] ), .c ({new_AGEMA_signal_994, n2643}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2036 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1045, n2442}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2038 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_995, n2739}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2044 ( .a ({new_AGEMA_signal_947, n2462}), .b ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .r ( Fresh[29] ), .c ({new_AGEMA_signal_996, n2437}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2045 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[4], SI_s0[4]}), .clk ( clk ), .r ( Fresh[30] ), .c ({new_AGEMA_signal_966, n2261}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2046 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_997, n2778}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2052 ( .a ({SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[31] ), .c ({new_AGEMA_signal_998, n2452}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2055 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_1050, n2766}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2068 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[32] ), .c ({new_AGEMA_signal_1000, n2772}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2070 ( .a ({new_AGEMA_signal_951, n2791}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[33] ), .c ({new_AGEMA_signal_1001, n2824}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2071 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1053, n2612}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2074 ( .a ({new_AGEMA_signal_988, n2400}), .b ({new_AGEMA_signal_1054, n2313}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2089 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[34] ), .c ({new_AGEMA_signal_1002, n2395}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2090 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1058, n2818}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2094 ( .a ({SI_s1[6], SI_s0[6]}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[35] ), .c ({new_AGEMA_signal_967, n2779}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2096 ( .a ({new_AGEMA_signal_955, n2630}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[36] ), .c ({new_AGEMA_signal_1003, n2624}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2097 ( .a ({SI_s1[4], SI_s0[4]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[37] ), .c ({new_AGEMA_signal_968, n2242}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2100 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[38] ), .c ({new_AGEMA_signal_1004, n2356}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2119 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_1063, n2823}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2122 ( .a ({new_AGEMA_signal_949, n2760}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[39] ), .c ({new_AGEMA_signal_1005, n2611}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2131 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1065, n2828}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2133 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[40] ), .c ({new_AGEMA_signal_1006, n2616}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2134 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1066, n2679}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2138 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[41] ), .c ({new_AGEMA_signal_1007, n2563}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2139 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1067, n2809}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2150 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_1068, n2709}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2163 ( .a ({new_AGEMA_signal_943, n2796}), .b ({new_AGEMA_signal_945, n2810}), .clk ( clk ), .r ( Fresh[42] ), .c ({new_AGEMA_signal_1008, n2401}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2211 ( .a ({new_AGEMA_signal_957, n2765}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[43] ), .c ({new_AGEMA_signal_1010, n2061}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2232 ( .a ({new_AGEMA_signal_943, n2796}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[44] ), .c ({new_AGEMA_signal_1011, n2721}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2276 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_957, n2765}), .clk ( clk ), .r ( Fresh[45] ), .c ({new_AGEMA_signal_1012, n2298}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2278 ( .a ({new_AGEMA_signal_1008, n2401}), .b ({new_AGEMA_signal_1080, n2118}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2307 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[46] ), .c ({new_AGEMA_signal_1013, n2346}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2341 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[47] ), .c ({new_AGEMA_signal_1015, n2430}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2383 ( .a ({SI_s1[5], SI_s0[5]}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[48] ), .c ({new_AGEMA_signal_969, n2712}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2402 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[49] ), .c ({new_AGEMA_signal_1017, n2777}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2615 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_947, n2462}), .clk ( clk ), .r ( Fresh[50] ), .c ({new_AGEMA_signal_1019, n2463}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2627 ( .a ({new_AGEMA_signal_945, n2810}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[51] ), .c ({new_AGEMA_signal_1020, n2474}) ) ;

    /* cells in depth 3 */

    /* cells in depth 4 */
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1954 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ( Fresh[52] ), .c ({new_AGEMA_signal_1127, n2575}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1959 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[53] ), .c ({new_AGEMA_signal_1128, n1962}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1964 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ( Fresh[54] ), .c ({new_AGEMA_signal_1129, n1922}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1974 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[55] ), .c ({new_AGEMA_signal_1030, n2755}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1977 ( .a ({new_AGEMA_signal_977, n2317}), .b ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .r ( Fresh[56] ), .c ({new_AGEMA_signal_1130, n1926}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1980 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1032, n2541}), .clk ( clk ), .r ( Fresh[57] ), .c ({new_AGEMA_signal_1131, n1925}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1986 ( .a ({new_AGEMA_signal_1033, n2086}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ( Fresh[58] ), .c ({new_AGEMA_signal_1132, n2151}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1988 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ( Fresh[59] ), .c ({new_AGEMA_signal_1034, n2631}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U1989 ( .a ({new_AGEMA_signal_1034, n2631}), .b ({new_AGEMA_signal_1133, n2734}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1992 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ( Fresh[60] ), .c ({new_AGEMA_signal_1134, n2763}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1997 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[61] ), .c ({new_AGEMA_signal_1036, n1930}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2005 ( .a ({new_AGEMA_signal_988, n2400}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ( Fresh[62] ), .c ({new_AGEMA_signal_1038, n2492}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2006 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_1135, n2732}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2010 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ( Fresh[63] ), .c ({new_AGEMA_signal_1136, n1937}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2022 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_992, n2493}), .clk ( clk ), .r ( Fresh[64] ), .c ({new_AGEMA_signal_1042, n1942}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(0)) U2026 ( .a ({new_AGEMA_signal_993, n2587}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ( Fresh[65] ), .c ({new_AGEMA_signal_1043, n2676}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2030 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ( Fresh[66] ), .c ({new_AGEMA_signal_1139, n1944}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2037 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[67] ), .c ({new_AGEMA_signal_1140, n1950}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2039 ( .a ({SI_s1[7], SI_s0[7]}), .b ({new_AGEMA_signal_995, n2739}), .clk ( clk ), .r ( Fresh[68] ), .c ({new_AGEMA_signal_1046, n1949}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2042 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ( Fresh[69] ), .c ({new_AGEMA_signal_1047, n2677}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2043 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_1141, n2662}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2047 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ( Fresh[70] ), .c ({new_AGEMA_signal_1048, n2627}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2053 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_998, n2452}), .clk ( clk ), .r ( Fresh[71] ), .c ({new_AGEMA_signal_1049, n1957}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2056 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ( Fresh[72] ), .c ({new_AGEMA_signal_1142, n2088}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2062 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ( Fresh[73] ), .c ({new_AGEMA_signal_999, n1964}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2063 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[74] ), .c ({new_AGEMA_signal_1051, n2736}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2069 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[75] ), .c ({new_AGEMA_signal_1052, n2673}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2072 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ( Fresh[76] ), .c ({new_AGEMA_signal_1144, n2761}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2073 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1323, n2720}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2075 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ( Fresh[77] ), .c ({new_AGEMA_signal_1145, n2412}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2076 ( .a ({new_AGEMA_signal_1145, n2412}), .b ({new_AGEMA_signal_1324, n2417}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2079 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_966, n2261}), .clk ( clk ), .r ( Fresh[78] ), .c ({new_AGEMA_signal_1055, n2571}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2080 ( .a ({new_AGEMA_signal_1055, n2571}), .b ({new_AGEMA_signal_1146, n2505}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2081 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .r ( Fresh[79] ), .c ({new_AGEMA_signal_1056, n2651}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2083 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[80] ), .c ({new_AGEMA_signal_1147, n2359}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2086 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ( Fresh[81] ), .c ({new_AGEMA_signal_1057, n2101}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2087 ( .a ({new_AGEMA_signal_1057, n2101}), .b ({new_AGEMA_signal_1148, n2625}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2091 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[82] ), .c ({new_AGEMA_signal_1059, n2190}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2095 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ( Fresh[83] ), .c ({new_AGEMA_signal_1060, n1976}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2098 ( .a ({new_AGEMA_signal_1023, n2672}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ( Fresh[84] ), .c ({new_AGEMA_signal_1150, n2535}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2101 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1004, n2356}), .clk ( clk ), .r ( Fresh[85] ), .c ({new_AGEMA_signal_1151, n1973}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2105 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ( Fresh[86] ), .c ({new_AGEMA_signal_1061, n2690}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2111 ( .a ({new_AGEMA_signal_992, n2493}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[87] ), .c ({new_AGEMA_signal_1062, n2817}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2113 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ( Fresh[88] ), .c ({new_AGEMA_signal_1153, n2741}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2118 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ( Fresh[89] ), .c ({new_AGEMA_signal_1154, n1992}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2120 ( .a ({new_AGEMA_signal_1063, n2823}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[90] ), .c ({new_AGEMA_signal_1155, n1991}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2123 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .r ( Fresh[91] ), .c ({new_AGEMA_signal_1064, n1993}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2125 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ( Fresh[92] ), .c ({new_AGEMA_signal_1156, n1995}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2132 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ( Fresh[93] ), .c ({new_AGEMA_signal_1157, n2241}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2135 ( .a ({SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_1066, n2679}), .clk ( clk ), .r ( Fresh[94] ), .c ({new_AGEMA_signal_1158, n2003}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2140 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .r ( Fresh[95] ), .c ({new_AGEMA_signal_1159, n2008}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2141 ( .a ({new_AGEMA_signal_1066, n2679}), .b ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .r ( Fresh[96] ), .c ({new_AGEMA_signal_1160, n2572}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2143 ( .a ({new_AGEMA_signal_1067, n2809}), .b ({new_AGEMA_signal_1004, n2356}), .clk ( clk ), .r ( Fresh[97] ), .c ({new_AGEMA_signal_1161, n2004}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2147 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[98] ), .c ({new_AGEMA_signal_1162, n2009}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2151 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[99] ), .c ({new_AGEMA_signal_1163, n2533}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2157 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[100] ), .c ({new_AGEMA_signal_1069, n2026}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2158 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_992, n2493}), .clk ( clk ), .r ( Fresh[101] ), .c ({new_AGEMA_signal_1164, n2022}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2159 ( .a ({new_AGEMA_signal_947, n2462}), .b ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .r ( Fresh[102] ), .c ({new_AGEMA_signal_1070, n2227}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2167 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[103] ), .c ({new_AGEMA_signal_1009, n2027}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2171 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ( Fresh[104] ), .c ({new_AGEMA_signal_1167, n2214}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2173 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[105] ), .c ({new_AGEMA_signal_1168, n2290}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2174 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[106] ), .c ({new_AGEMA_signal_1169, n2376}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2178 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_988, n2400}), .clk ( clk ), .r ( Fresh[107] ), .c ({new_AGEMA_signal_1072, n2034}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2182 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ( Fresh[108] ), .c ({new_AGEMA_signal_1073, n2171}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2183 ( .a ({new_AGEMA_signal_1065, n2828}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[109] ), .c ({new_AGEMA_signal_1170, n2039}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2188 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[110] ), .c ({new_AGEMA_signal_1172, n2042}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2191 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ( Fresh[111] ), .c ({new_AGEMA_signal_1173, n2754}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2192 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_959, n2790}), .clk ( clk ), .r ( Fresh[112] ), .c ({new_AGEMA_signal_1174, n2044}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2198 ( .a ({new_AGEMA_signal_1054, n2313}), .b ({new_AGEMA_signal_971, n2641}), .clk ( clk ), .r ( Fresh[113] ), .c ({new_AGEMA_signal_1175, n2654}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2202 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1037, n2577}), .clk ( clk ), .r ( Fresh[114] ), .c ({new_AGEMA_signal_1176, n2055}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2205 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[115] ), .c ({new_AGEMA_signal_1177, n2057}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2208 ( .a ({new_AGEMA_signal_1066, n2679}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[116] ), .c ({new_AGEMA_signal_1178, n2407}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2212 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1010, n2061}), .clk ( clk ), .r ( Fresh[117] ), .c ({new_AGEMA_signal_1179, n2062}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2216 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ( Fresh[118] ), .c ({new_AGEMA_signal_1180, n2731}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2220 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1181, n2068}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2224 ( .a ({new_AGEMA_signal_1005, n2611}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ( Fresh[119] ), .c ({new_AGEMA_signal_1074, n2642}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2225 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ( Fresh[120] ), .c ({new_AGEMA_signal_1182, n2252}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2228 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ( Fresh[121] ), .c ({new_AGEMA_signal_1075, n2075}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(0)) U2233 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .r ( Fresh[122] ), .c ({new_AGEMA_signal_1076, n2081}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2234 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[123] ), .c ({new_AGEMA_signal_1183, n2080}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2237 ( .a ({new_AGEMA_signal_984, n2600}), .b ({new_AGEMA_signal_970, n2719}), .clk ( clk ), .r ( Fresh[124] ), .c ({new_AGEMA_signal_1077, n2498}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2238 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_1184, n2773}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2239 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ( Fresh[125] ), .c ({new_AGEMA_signal_1185, n2083}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2244 ( .a ({SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_1033, n2086}), .clk ( clk ), .r ( Fresh[126] ), .c ({new_AGEMA_signal_1186, n2562}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2247 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .r ( Fresh[127] ), .c ({new_AGEMA_signal_1078, n2087}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2251 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1041, n2174}), .clk ( clk ), .r ( Fresh[128] ), .c ({new_AGEMA_signal_1187, n2156}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2260 ( .a ({new_AGEMA_signal_1028, n2769}), .b ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .r ( Fresh[129] ), .c ({new_AGEMA_signal_1188, n2100}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2277 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_1012, n2298}), .clk ( clk ), .r ( Fresh[130] ), .c ({new_AGEMA_signal_1079, n2544}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2279 ( .a ({new_AGEMA_signal_1004, n2356}), .b ({new_AGEMA_signal_1080, n2118}), .clk ( clk ), .r ( Fresh[131] ), .c ({new_AGEMA_signal_1191, n2121}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2284 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ( Fresh[132] ), .c ({new_AGEMA_signal_1193, n2122}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2286 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ( Fresh[133] ), .c ({new_AGEMA_signal_1194, n2811}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2294 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[134] ), .c ({new_AGEMA_signal_1081, n2647}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2297 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ( Fresh[135] ), .c ({new_AGEMA_signal_1082, n2132}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2304 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[136] ), .c ({new_AGEMA_signal_1199, n2220}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2305 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[137] ), .c ({new_AGEMA_signal_1200, n2138}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2312 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[138] ), .c ({new_AGEMA_signal_1201, n2555}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2322 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .r ( Fresh[139] ), .c ({new_AGEMA_signal_1202, n2429}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2328 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[140] ), .c ({new_AGEMA_signal_1083, n2162}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2337 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ( Fresh[141] ), .c ({new_AGEMA_signal_1014, n2545}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2340 ( .a ({new_AGEMA_signal_965, n2559}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[142] ), .c ({new_AGEMA_signal_1085, n2178}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2342 ( .a ({new_AGEMA_signal_1015, n2430}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[143] ), .c ({new_AGEMA_signal_1204, n2176}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2343 ( .a ({new_AGEMA_signal_1041, n2174}), .b ({SI_s1[5], SI_s0[5]}), .clk ( clk ), .r ( Fresh[144] ), .c ({new_AGEMA_signal_1205, n2175}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2348 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .r ( Fresh[145] ), .c ({new_AGEMA_signal_1016, n2182}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2353 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_1015, n2430}), .clk ( clk ), .r ( Fresh[146] ), .c ({new_AGEMA_signal_1206, n2188}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2355 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ( Fresh[147] ), .c ({new_AGEMA_signal_1207, n2189}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2357 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[148] ), .c ({new_AGEMA_signal_1208, n2446}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2362 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_965, n2559}), .clk ( clk ), .r ( Fresh[149] ), .c ({new_AGEMA_signal_1087, n2576}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2363 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_957, n2765}), .clk ( clk ), .r ( Fresh[150] ), .c ({new_AGEMA_signal_1088, n2748}) ) ;
    not_masked #(.low_latency(0), .pipeline(0)) U2368 ( .a ({new_AGEMA_signal_1175, n2654}), .b ({new_AGEMA_signal_1375, n2674}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2378 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ( Fresh[151] ), .c ({new_AGEMA_signal_1089, n2213}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2380 ( .a ({new_AGEMA_signal_975, n2816}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[152] ), .c ({new_AGEMA_signal_1090, n2215}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2384 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[153] ), .c ({new_AGEMA_signal_1211, n2218}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2386 ( .a ({new_AGEMA_signal_1012, n2298}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[154] ), .c ({new_AGEMA_signal_1212, n2219}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2405 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[155] ), .c ({new_AGEMA_signal_1217, n2240}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2407 ( .a ({new_AGEMA_signal_1068, n2709}), .b ({new_AGEMA_signal_968, n2242}), .clk ( clk ), .r ( Fresh[156] ), .c ({new_AGEMA_signal_1218, n2561}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2408 ( .a ({SI_s1[5], SI_s0[5]}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ( Fresh[157] ), .c ({new_AGEMA_signal_1219, n2243}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2411 ( .a ({new_AGEMA_signal_973, n2615}), .b ({new_AGEMA_signal_1045, n2442}), .clk ( clk ), .r ( Fresh[158] ), .c ({new_AGEMA_signal_1220, n2245}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2422 ( .a ({new_AGEMA_signal_1023, n2672}), .b ({new_AGEMA_signal_1015, n2430}), .clk ( clk ), .r ( Fresh[159] ), .c ({new_AGEMA_signal_1221, n2540}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2423 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ( Fresh[160] ), .c ({new_AGEMA_signal_1222, n2259}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2426 ( .a ({new_AGEMA_signal_966, n2261}), .b ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .r ( Fresh[161] ), .c ({new_AGEMA_signal_1091, n2262}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2431 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ( Fresh[162] ), .c ({new_AGEMA_signal_1092, n2266}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2432 ( .a ({new_AGEMA_signal_1000, n2772}), .b ({new_AGEMA_signal_943, n2796}), .clk ( clk ), .r ( Fresh[163] ), .c ({new_AGEMA_signal_1093, n2645}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2436 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .r ( Fresh[164] ), .c ({new_AGEMA_signal_1094, n2268}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2443 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_1035, n2786}), .clk ( clk ), .r ( Fresh[165] ), .c ({new_AGEMA_signal_1225, n2278}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2448 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[166] ), .c ({new_AGEMA_signal_1095, n2383}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2455 ( .a ({new_AGEMA_signal_997, n2778}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ( Fresh[167] ), .c ({new_AGEMA_signal_1228, n2774}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2458 ( .a ({new_AGEMA_signal_1063, n2823}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ( Fresh[168] ), .c ({new_AGEMA_signal_1229, n2287}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2470 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[169] ), .c ({new_AGEMA_signal_1231, n2438}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2471 ( .a ({new_AGEMA_signal_1012, n2298}), .b ({new_AGEMA_signal_961, n2315}), .clk ( clk ), .r ( Fresh[170] ), .c ({new_AGEMA_signal_1096, n2299}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2481 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_1054, n2313}), .clk ( clk ), .r ( Fresh[171] ), .c ({new_AGEMA_signal_1232, n2371}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2484 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ( Fresh[172] ), .c ({new_AGEMA_signal_1018, n2316}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2486 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_977, n2317}), .clk ( clk ), .r ( Fresh[173] ), .c ({new_AGEMA_signal_1098, n2318}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2492 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[174] ), .c ({new_AGEMA_signal_1235, n2325}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2494 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[175] ), .c ({new_AGEMA_signal_1236, n2328}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2495 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .r ( Fresh[176] ), .c ({new_AGEMA_signal_1099, n2327}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2505 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_978, n2694}), .clk ( clk ), .r ( Fresh[177] ), .c ({new_AGEMA_signal_1237, n2343}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2510 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[178] ), .c ({new_AGEMA_signal_1239, n2344}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) U2512 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_1013, n2346}), .clk ( clk ), .r ( Fresh[179] ), .c ({new_AGEMA_signal_1100, n2348}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2513 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ( Fresh[180] ), .c ({new_AGEMA_signal_1101, n2347}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2520 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .r ( Fresh[181] ), .c ({new_AGEMA_signal_1102, n2363}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2521 ( .a ({new_AGEMA_signal_1067, n2809}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[182] ), .c ({new_AGEMA_signal_1243, n2353}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2524 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[183] ), .c ({new_AGEMA_signal_1244, n2355}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2530 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[184] ), .c ({new_AGEMA_signal_1245, n2364}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2543 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .r ( Fresh[185] ), .c ({new_AGEMA_signal_1103, n2415}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2558 ( .a ({new_AGEMA_signal_1002, n2395}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ( Fresh[186] ), .c ({new_AGEMA_signal_1104, n2700}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2563 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_988, n2400}), .clk ( clk ), .r ( Fresh[187] ), .c ({new_AGEMA_signal_1105, n2594}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2564 ( .a ({new_AGEMA_signal_1008, n2401}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[188] ), .c ({new_AGEMA_signal_1106, n2402}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2585 ( .a ({new_AGEMA_signal_969, n2712}), .b ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .r ( Fresh[189] ), .c ({new_AGEMA_signal_1255, n2428}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2588 ( .a ({new_AGEMA_signal_1015, n2430}), .b ({new_AGEMA_signal_1044, n2570}), .clk ( clk ), .r ( Fresh[190] ), .c ({new_AGEMA_signal_1256, n2431}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2594 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ( Fresh[191] ), .c ({new_AGEMA_signal_1107, n2483}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2599 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[192] ), .c ({new_AGEMA_signal_1258, n2443}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2606 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[193] ), .c ({new_AGEMA_signal_1259, n2693}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2608 ( .a ({new_AGEMA_signal_998, n2452}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[194] ), .c ({new_AGEMA_signal_1108, n2453}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2616 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1019, n2463}), .clk ( clk ), .r ( Fresh[195] ), .c ({new_AGEMA_signal_1109, n2464}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2620 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[196] ), .c ({new_AGEMA_signal_1110, n2468}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2624 ( .a ({new_AGEMA_signal_997, n2778}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[197] ), .c ({new_AGEMA_signal_1111, n2473}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2625 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ( Fresh[198] ), .c ({new_AGEMA_signal_1112, n2472}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2628 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1020, n2474}), .clk ( clk ), .r ( Fresh[199] ), .c ({new_AGEMA_signal_1113, n2475}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2632 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_1065, n2828}), .clk ( clk ), .r ( Fresh[200] ), .c ({new_AGEMA_signal_1263, n2480}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2638 ( .a ({new_AGEMA_signal_1037, n2577}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ( Fresh[201] ), .c ({new_AGEMA_signal_1264, n2487}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2641 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .r ( Fresh[202] ), .c ({new_AGEMA_signal_1114, n2488}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2665 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_960, n2519}), .clk ( clk ), .r ( Fresh[203] ), .c ({new_AGEMA_signal_1270, n2520}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2667 ( .a ({new_AGEMA_signal_980, n2713}), .b ({new_AGEMA_signal_993, n2587}), .clk ( clk ), .r ( Fresh[204] ), .c ({new_AGEMA_signal_1115, n2521}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2674 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_963, n2595}), .clk ( clk ), .r ( Fresh[205] ), .c ({new_AGEMA_signal_1271, n2531}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2689 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ( Fresh[206] ), .c ({new_AGEMA_signal_1273, n2553}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2691 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1039, n2792}), .clk ( clk ), .r ( Fresh[207] ), .c ({new_AGEMA_signal_1274, n2554}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) U2695 ( .a ({new_AGEMA_signal_965, n2559}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[208] ), .c ({new_AGEMA_signal_1116, n2560}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2698 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_1007, n2563}), .clk ( clk ), .r ( Fresh[209] ), .c ({new_AGEMA_signal_1275, n2564}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2714 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_978, n2694}), .clk ( clk ), .r ( Fresh[210] ), .c ({new_AGEMA_signal_1278, n2586}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2720 ( .a ({new_AGEMA_signal_963, n2595}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[211] ), .c ({new_AGEMA_signal_1117, n2597}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2721 ( .a ({new_AGEMA_signal_1024, n2640}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ( Fresh[212] ), .c ({new_AGEMA_signal_1280, n2596}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2723 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_976, n2780}), .clk ( clk ), .r ( Fresh[213] ), .c ({new_AGEMA_signal_1281, n2598}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2725 ( .a ({new_AGEMA_signal_958, n2635}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[214] ), .c ({new_AGEMA_signal_1021, n2599}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2732 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1058, n2818}), .clk ( clk ), .r ( Fresh[215] ), .c ({new_AGEMA_signal_1283, n2610}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2734 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .r ( Fresh[216] ), .c ({new_AGEMA_signal_1284, n2614}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2735 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ( Fresh[217] ), .c ({new_AGEMA_signal_1285, n2613}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2737 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ( Fresh[218] ), .c ({new_AGEMA_signal_1119, n2617}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2742 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_972, n2750}), .clk ( clk ), .r ( Fresh[219] ), .c ({new_AGEMA_signal_1120, n2629}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2751 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1024, n2640}), .clk ( clk ), .r ( Fresh[220] ), .c ({new_AGEMA_signal_1287, n2784}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2757 ( .a ({new_AGEMA_signal_989, n2785}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ( Fresh[221] ), .c ({new_AGEMA_signal_1121, n2650}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2775 ( .a ({new_AGEMA_signal_949, n2760}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[222] ), .c ({new_AGEMA_signal_1022, n2683}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2789 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1029, n2707}), .clk ( clk ), .r ( Fresh[223] ), .c ({new_AGEMA_signal_1294, n2711}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2790 ( .a ({new_AGEMA_signal_1068, n2709}), .b ({new_AGEMA_signal_964, n2708}), .clk ( clk ), .r ( Fresh[224] ), .c ({new_AGEMA_signal_1295, n2710}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2792 ( .a ({new_AGEMA_signal_980, n2713}), .b ({new_AGEMA_signal_969, n2712}), .clk ( clk ), .r ( Fresh[225] ), .c ({new_AGEMA_signal_1122, n2714}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2797 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1011, n2721}), .clk ( clk ), .r ( Fresh[226] ), .c ({new_AGEMA_signal_1123, n2722}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2799 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1040, n2724}), .clk ( clk ), .r ( Fresh[227] ), .c ({new_AGEMA_signal_1297, n2726}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2806 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .r ( Fresh[228] ), .c ({new_AGEMA_signal_1298, n2738}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2822 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1050, n2766}), .clk ( clk ), .r ( Fresh[229] ), .c ({new_AGEMA_signal_1301, n2768}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2828 ( .a ({new_AGEMA_signal_997, n2778}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ( Fresh[230] ), .c ({new_AGEMA_signal_1124, n2782}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2829 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ( Fresh[231] ), .c ({new_AGEMA_signal_1125, n2781}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2832 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_989, n2785}), .clk ( clk ), .r ( Fresh[232] ), .c ({new_AGEMA_signal_1303, n2787}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2834 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ( Fresh[233] ), .c ({new_AGEMA_signal_1304, n2794}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2835 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[234] ), .c ({new_AGEMA_signal_1305, n2793}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2844 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .r ( Fresh[235] ), .c ({new_AGEMA_signal_1306, n2812}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2847 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_983, n2815}), .clk ( clk ), .r ( Fresh[236] ), .c ({new_AGEMA_signal_1126, n2820}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2851 ( .a ({new_AGEMA_signal_1001, n2824}), .b ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .r ( Fresh[237] ), .c ({new_AGEMA_signal_1308, n2825}) ) ;

    /* cells in depth 5 */

    /* cells in depth 6 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1960 ( .a ({new_AGEMA_signal_1127, n2575}), .b ({new_AGEMA_signal_1128, n1962}), .clk ( clk ), .r ( Fresh[238] ), .c ({new_AGEMA_signal_1309, n1924}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1967 ( .a ({new_AGEMA_signal_1129, n1922}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[239] ), .c ({new_AGEMA_signal_1310, n1923}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1981 ( .a ({new_AGEMA_signal_1130, n1926}), .b ({new_AGEMA_signal_1131, n1925}), .clk ( clk ), .r ( Fresh[240] ), .c ({new_AGEMA_signal_1311, n1927}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1993 ( .a ({new_AGEMA_signal_1133, n2734}), .b ({new_AGEMA_signal_1134, n2763}), .clk ( clk ), .r ( Fresh[241] ), .c ({new_AGEMA_signal_1312, n1929}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2007 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ( Fresh[242] ), .c ({new_AGEMA_signal_1313, n2665}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2011 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_1136, n1937}), .clk ( clk ), .r ( Fresh[243] ), .c ({new_AGEMA_signal_1314, n1938}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2019 ( .a ({new_AGEMA_signal_1041, n2174}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ( Fresh[244] ), .c ({new_AGEMA_signal_1315, n2235}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2023 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_1042, n1942}), .clk ( clk ), .r ( Fresh[245] ), .c ({new_AGEMA_signal_1137, n1943}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2027 ( .a ({new_AGEMA_signal_1043, n2676}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[246] ), .c ({new_AGEMA_signal_1138, n1946}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2031 ( .a ({new_AGEMA_signal_1044, n2570}), .b ({new_AGEMA_signal_1139, n1944}), .clk ( clk ), .r ( Fresh[247] ), .c ({new_AGEMA_signal_1316, n1945}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2034 ( .a ({new_AGEMA_signal_1039, n2792}), .b ({new_AGEMA_signal_1133, n2734}), .clk ( clk ), .r ( Fresh[248] ), .c ({new_AGEMA_signal_1317, n1956}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2040 ( .a ({new_AGEMA_signal_1140, n1950}), .b ({new_AGEMA_signal_1046, n1949}), .clk ( clk ), .r ( Fresh[249] ), .c ({new_AGEMA_signal_1318, n1951}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2048 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .r ( Fresh[250] ), .c ({new_AGEMA_signal_1319, n1952}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2057 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1142, n2088}), .clk ( clk ), .r ( Fresh[251] ), .c ({new_AGEMA_signal_1320, n2687}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(0)) U2061 ( .a ({new_AGEMA_signal_1128, n1962}), .b ({new_AGEMA_signal_993, n2587}), .clk ( clk ), .r ( Fresh[252] ), .c ({new_AGEMA_signal_1321, n1966}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2064 ( .a ({new_AGEMA_signal_1051, n2736}), .b ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .r ( Fresh[253] ), .c ({new_AGEMA_signal_1143, n1963}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2077 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .r ( Fresh[254] ), .c ({new_AGEMA_signal_1480, n1968}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2082 ( .a ({new_AGEMA_signal_1146, n2505}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[255] ), .c ({new_AGEMA_signal_1325, n2684}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2088 ( .a ({new_AGEMA_signal_964, n2708}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ( Fresh[256] ), .c ({new_AGEMA_signal_1326, n1972}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2092 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_1059, n2190}), .clk ( clk ), .r ( Fresh[257] ), .c ({new_AGEMA_signal_1149, n1971}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2099 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1150, n2535}), .clk ( clk ), .r ( Fresh[258] ), .c ({new_AGEMA_signal_1327, n1974}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2106 ( .a ({new_AGEMA_signal_1135, n2732}), .b ({new_AGEMA_signal_958, n2635}), .clk ( clk ), .r ( Fresh[259] ), .c ({new_AGEMA_signal_1328, n1979}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2112 ( .a ({new_AGEMA_signal_1035, n2786}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[260] ), .c ({new_AGEMA_signal_1152, n1985}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2121 ( .a ({new_AGEMA_signal_1154, n1992}), .b ({new_AGEMA_signal_1155, n1991}), .clk ( clk ), .r ( Fresh[261] ), .c ({new_AGEMA_signal_1330, n1994}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2126 ( .a ({new_AGEMA_signal_988, n2400}), .b ({new_AGEMA_signal_1156, n1995}), .clk ( clk ), .r ( Fresh[262] ), .c ({new_AGEMA_signal_1331, n1996}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2136 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_1158, n2003}), .clk ( clk ), .r ( Fresh[263] ), .c ({new_AGEMA_signal_1332, n2137}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2142 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_1160, n2572}), .clk ( clk ), .r ( Fresh[264] ), .c ({new_AGEMA_signal_1333, n2006}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2144 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1161, n2004}), .clk ( clk ), .r ( Fresh[265] ), .c ({new_AGEMA_signal_1334, n2005}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2152 ( .a ({new_AGEMA_signal_1068, n2709}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[266] ), .c ({new_AGEMA_signal_1335, n2013}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2160 ( .a ({new_AGEMA_signal_987, n2753}), .b ({new_AGEMA_signal_1070, n2227}), .clk ( clk ), .r ( Fresh[267] ), .c ({new_AGEMA_signal_1165, n2020}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2164 ( .a ({new_AGEMA_signal_1062, n2817}), .b ({new_AGEMA_signal_1008, n2401}), .clk ( clk ), .r ( Fresh[268] ), .c ({new_AGEMA_signal_1166, n2023}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2168 ( .a ({new_AGEMA_signal_1009, n2027}), .b ({new_AGEMA_signal_957, n2765}), .clk ( clk ), .r ( Fresh[269] ), .c ({new_AGEMA_signal_1071, n2028}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2172 ( .a ({new_AGEMA_signal_1167, n2214}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[270] ), .c ({new_AGEMA_signal_1337, n2033}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2175 ( .a ({new_AGEMA_signal_1169, n2376}), .b ({new_AGEMA_signal_973, n2615}), .clk ( clk ), .r ( Fresh[271] ), .c ({new_AGEMA_signal_1338, n2031}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2184 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_1170, n2039}), .clk ( clk ), .r ( Fresh[272] ), .c ({new_AGEMA_signal_1339, n2040}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2187 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[273] ), .c ({new_AGEMA_signal_1171, n2050}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2193 ( .a ({new_AGEMA_signal_1007, n2563}), .b ({new_AGEMA_signal_1174, n2044}), .clk ( clk ), .r ( Fresh[274] ), .c ({new_AGEMA_signal_1340, n2045}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2199 ( .a ({new_AGEMA_signal_1175, n2654}), .b ({new_AGEMA_signal_958, n2635}), .clk ( clk ), .r ( Fresh[275] ), .c ({new_AGEMA_signal_1341, n2051}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2203 ( .a ({new_AGEMA_signal_1053, n2612}), .b ({new_AGEMA_signal_1176, n2055}), .clk ( clk ), .r ( Fresh[276] ), .c ({new_AGEMA_signal_1342, n2056}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2209 ( .a ({new_AGEMA_signal_1178, n2407}), .b ({new_AGEMA_signal_1001, n2824}), .clk ( clk ), .r ( Fresh[277] ), .c ({new_AGEMA_signal_1343, n2060}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2215 ( .a ({new_AGEMA_signal_975, n2816}), .b ({new_AGEMA_signal_1175, n2654}), .clk ( clk ), .r ( Fresh[278] ), .c ({new_AGEMA_signal_1344, n2066}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2217 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ( Fresh[279] ), .c ({new_AGEMA_signal_1345, n2065}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2221 ( .a ({new_AGEMA_signal_1181, n2068}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[280] ), .c ({new_AGEMA_signal_1346, n2069}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2226 ( .a ({new_AGEMA_signal_979, n2073}), .b ({new_AGEMA_signal_1182, n2252}), .clk ( clk ), .r ( Fresh[281] ), .c ({new_AGEMA_signal_1347, n2074}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2235 ( .a ({new_AGEMA_signal_1076, n2081}), .b ({new_AGEMA_signal_1183, n2080}), .clk ( clk ), .r ( Fresh[282] ), .c ({new_AGEMA_signal_1348, n2082}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2240 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1185, n2083}), .clk ( clk ), .r ( Fresh[283] ), .c ({new_AGEMA_signal_1349, n2084}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2242 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[284] ), .c ({new_AGEMA_signal_1350, n2085}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2245 ( .a ({new_AGEMA_signal_960, n2519}), .b ({new_AGEMA_signal_1186, n2562}), .clk ( clk ), .r ( Fresh[285] ), .c ({new_AGEMA_signal_1351, n2131}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2248 ( .a ({new_AGEMA_signal_1142, n2088}), .b ({new_AGEMA_signal_1078, n2087}), .clk ( clk ), .r ( Fresh[286] ), .c ({new_AGEMA_signal_1352, n2089}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2252 ( .a ({new_AGEMA_signal_955, n2630}), .b ({new_AGEMA_signal_1187, n2156}), .clk ( clk ), .r ( Fresh[287] ), .c ({new_AGEMA_signal_1353, n2330}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2254 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1132, n2151}), .clk ( clk ), .r ( Fresh[288] ), .c ({new_AGEMA_signal_1354, n2092}) ) ;
    or_GHPC #(.low_latency(0), .pipeline(0)) U2256 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1147, n2359}), .clk ( clk ), .r ( Fresh[289] ), .c ({new_AGEMA_signal_1355, n2094}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2261 ( .a ({new_AGEMA_signal_1057, n2101}), .b ({new_AGEMA_signal_1188, n2100}), .clk ( clk ), .r ( Fresh[290] ), .c ({new_AGEMA_signal_1356, n2160}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2265 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[291] ), .c ({new_AGEMA_signal_1189, n2504}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2271 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[292] ), .c ({new_AGEMA_signal_1504, n2114}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2273 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_981, n2723}), .clk ( clk ), .r ( Fresh[293] ), .c ({new_AGEMA_signal_1190, n2115}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2280 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ( Fresh[294] ), .c ({new_AGEMA_signal_1358, n2291}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2281 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ( Fresh[295] ), .c ({new_AGEMA_signal_1192, n2119}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2291 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ( Fresh[296] ), .c ({new_AGEMA_signal_1195, n2130}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2292 ( .a ({new_AGEMA_signal_1062, n2817}), .b ({new_AGEMA_signal_1034, n2631}), .clk ( clk ), .r ( Fresh[297] ), .c ({new_AGEMA_signal_1196, n2129}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2295 ( .a ({new_AGEMA_signal_1081, n2647}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[298] ), .c ({new_AGEMA_signal_1197, n2150}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2298 ( .a ({new_AGEMA_signal_1038, n2492}), .b ({new_AGEMA_signal_1082, n2132}), .clk ( clk ), .r ( Fresh[299] ), .c ({new_AGEMA_signal_1198, n2133}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2302 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[300] ), .c ({new_AGEMA_signal_1361, n2136}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2306 ( .a ({new_AGEMA_signal_1160, n2572}), .b ({new_AGEMA_signal_1200, n2138}), .clk ( clk ), .r ( Fresh[301] ), .c ({new_AGEMA_signal_1362, n2139}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2313 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_1201, n2555}), .clk ( clk ), .r ( Fresh[302] ), .c ({new_AGEMA_signal_1363, n2144}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2318 ( .a ({new_AGEMA_signal_1132, n2151}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[303] ), .c ({new_AGEMA_signal_1364, n2152}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2321 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_1187, n2156}), .clk ( clk ), .r ( Fresh[304] ), .c ({new_AGEMA_signal_1365, n2170}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2323 ( .a ({new_AGEMA_signal_1202, n2429}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ( Fresh[305] ), .c ({new_AGEMA_signal_1366, n2157}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2329 ( .a ({new_AGEMA_signal_977, n2317}), .b ({new_AGEMA_signal_1083, n2162}), .clk ( clk ), .r ( Fresh[306] ), .c ({new_AGEMA_signal_1203, n2163}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2335 ( .a ({new_AGEMA_signal_1073, n2171}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ( Fresh[307] ), .c ({new_AGEMA_signal_1368, n2172}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2338 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_1014, n2545}), .clk ( clk ), .r ( Fresh[308] ), .c ({new_AGEMA_signal_1084, n2186}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2339 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1168, n2290}), .clk ( clk ), .r ( Fresh[309] ), .c ({new_AGEMA_signal_1369, n2181}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2344 ( .a ({new_AGEMA_signal_1204, n2176}), .b ({new_AGEMA_signal_1205, n2175}), .clk ( clk ), .r ( Fresh[310] ), .c ({new_AGEMA_signal_1370, n2177}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2349 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1016, n2182}), .clk ( clk ), .r ( Fresh[311] ), .c ({new_AGEMA_signal_1086, n2183}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2354 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1206, n2188}), .clk ( clk ), .r ( Fresh[312] ), .c ({new_AGEMA_signal_1371, n2195}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2356 ( .a ({new_AGEMA_signal_1059, n2190}), .b ({new_AGEMA_signal_1207, n2189}), .clk ( clk ), .r ( Fresh[313] ), .c ({new_AGEMA_signal_1372, n2193}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2358 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_1208, n2446}), .clk ( clk ), .r ( Fresh[314] ), .c ({new_AGEMA_signal_1373, n2191}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2364 ( .a ({new_AGEMA_signal_1087, n2576}), .b ({new_AGEMA_signal_1088, n2748}), .clk ( clk ), .r ( Fresh[315] ), .c ({new_AGEMA_signal_1209, n2196}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2367 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1146, n2505}), .clk ( clk ), .r ( Fresh[316] ), .c ({new_AGEMA_signal_1374, n2201}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2369 ( .a ({new_AGEMA_signal_1375, n2674}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[317] ), .c ({new_AGEMA_signal_1515, n2200}) ) ;
    mux2_GHPC #(.low_latency(0), .pipeline(0)) U2371 ( .s ({new_AGEMA_signal_953, n2813}), .b ({new_AGEMA_signal_1133, n2734}), .a ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .r ( Fresh[318] ), .c ({new_AGEMA_signal_1516, n2202}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2379 ( .a ({new_AGEMA_signal_1167, n2214}), .b ({new_AGEMA_signal_1089, n2213}), .clk ( clk ), .r ( Fresh[319] ), .c ({new_AGEMA_signal_1376, n2217}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2381 ( .a ({new_AGEMA_signal_1024, n2640}), .b ({new_AGEMA_signal_1090, n2215}), .clk ( clk ), .r ( Fresh[320] ), .c ({new_AGEMA_signal_1210, n2216}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2385 ( .a ({new_AGEMA_signal_1211, n2218}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[321] ), .c ({new_AGEMA_signal_1377, n2222}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2387 ( .a ({new_AGEMA_signal_1199, n2220}), .b ({new_AGEMA_signal_1212, n2219}), .clk ( clk ), .r ( Fresh[322] ), .c ({new_AGEMA_signal_1378, n2221}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2391 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[323] ), .c ({new_AGEMA_signal_1213, n2226}) ) ;
    mux2_GHPC #(.low_latency(0), .pipeline(0)) U2393 ( .s ({new_AGEMA_signal_953, n2813}), .b ({new_AGEMA_signal_1056, n2651}), .a ({new_AGEMA_signal_1070, n2227}), .clk ( clk ), .r ( Fresh[324] ), .c ({new_AGEMA_signal_1214, n2228}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2397 ( .a ({new_AGEMA_signal_987, n2753}), .b ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[325] ), .c ({new_AGEMA_signal_1215, n2237}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2398 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[326] ), .c ({new_AGEMA_signal_1520, n2233}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2403 ( .a ({new_AGEMA_signal_1017, n2777}), .b ({new_AGEMA_signal_1034, n2631}), .clk ( clk ), .r ( Fresh[327] ), .c ({new_AGEMA_signal_1216, n2238}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2406 ( .a ({new_AGEMA_signal_1157, n2241}), .b ({new_AGEMA_signal_1217, n2240}), .clk ( clk ), .r ( Fresh[328] ), .c ({new_AGEMA_signal_1380, n2248}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2409 ( .a ({new_AGEMA_signal_1218, n2561}), .b ({new_AGEMA_signal_1219, n2243}), .clk ( clk ), .r ( Fresh[329] ), .c ({new_AGEMA_signal_1381, n2244}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2414 ( .a ({new_AGEMA_signal_1169, n2376}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[330] ), .c ({new_AGEMA_signal_1382, n2249}) ) ;
    mux2_GHPC #(.low_latency(0), .pipeline(0)) U2417 ( .s ({new_AGEMA_signal_953, n2813}), .b ({new_AGEMA_signal_1182, n2252}), .a ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[331] ), .c ({new_AGEMA_signal_1383, n2253}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2424 ( .a ({new_AGEMA_signal_1163, n2533}), .b ({new_AGEMA_signal_1222, n2259}), .clk ( clk ), .r ( Fresh[332] ), .c ({new_AGEMA_signal_1384, n2260}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2429 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ( Fresh[333] ), .c ({new_AGEMA_signal_1524, n2273}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2430 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1323, n2720}), .clk ( clk ), .r ( Fresh[334] ), .c ({new_AGEMA_signal_1525, n2752}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2433 ( .a ({new_AGEMA_signal_1093, n2645}), .b ({new_AGEMA_signal_951, n2791}), .clk ( clk ), .r ( Fresh[335] ), .c ({new_AGEMA_signal_1223, n2265}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2437 ( .a ({new_AGEMA_signal_947, n2462}), .b ({new_AGEMA_signal_1094, n2268}), .clk ( clk ), .r ( Fresh[336] ), .c ({new_AGEMA_signal_1224, n2269}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2444 ( .a ({new_AGEMA_signal_982, n2725}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[337] ), .c ({new_AGEMA_signal_1226, n2277}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2449 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1095, n2383}), .clk ( clk ), .r ( Fresh[338] ), .c ({new_AGEMA_signal_1227, n2282}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2452 ( .a ({new_AGEMA_signal_1051, n2736}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[339] ), .c ({new_AGEMA_signal_1389, n2284}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2456 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[340] ), .c ({new_AGEMA_signal_1390, n2459}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2459 ( .a ({SI_s1[6], SI_s0[6]}), .b ({new_AGEMA_signal_1229, n2287}), .clk ( clk ), .r ( Fresh[341] ), .c ({new_AGEMA_signal_1391, n2288}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2462 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_1144, n2761}), .clk ( clk ), .r ( Fresh[342] ), .c ({new_AGEMA_signal_1392, n2458}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2464 ( .a ({new_AGEMA_signal_977, n2317}), .b ({new_AGEMA_signal_1168, n2290}), .clk ( clk ), .r ( Fresh[343] ), .c ({new_AGEMA_signal_1393, n2293}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2467 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1074, n2642}), .clk ( clk ), .r ( Fresh[344] ), .c ({new_AGEMA_signal_1230, n2294}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2472 ( .a ({new_AGEMA_signal_1231, n2438}), .b ({new_AGEMA_signal_1096, n2299}), .clk ( clk ), .r ( Fresh[345] ), .c ({new_AGEMA_signal_1394, n2300}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2480 ( .a ({new_AGEMA_signal_1133, n2734}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[346] ), .c ({new_AGEMA_signal_1395, n2323}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) U2482 ( .a ({new_AGEMA_signal_1055, n2571}), .b ({new_AGEMA_signal_1232, n2371}), .clk ( clk ), .r ( Fresh[347] ), .c ({new_AGEMA_signal_1396, n2314}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2485 ( .a ({new_AGEMA_signal_1018, n2316}), .b ({new_AGEMA_signal_962, n2682}), .clk ( clk ), .r ( Fresh[348] ), .c ({new_AGEMA_signal_1097, n2319}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2491 ( .a ({new_AGEMA_signal_1074, n2642}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ( Fresh[349] ), .c ({new_AGEMA_signal_1234, n2326}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2496 ( .a ({new_AGEMA_signal_1236, n2328}), .b ({new_AGEMA_signal_1099, n2327}), .clk ( clk ), .r ( Fresh[350] ), .c ({new_AGEMA_signal_1398, n2329}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2501 ( .a ({new_AGEMA_signal_1324, n2417}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ( Fresh[351] ), .c ({new_AGEMA_signal_1537, n2335}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2506 ( .a ({new_AGEMA_signal_1068, n2709}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ( Fresh[352] ), .c ({new_AGEMA_signal_1399, n2341}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2507 ( .a ({new_AGEMA_signal_945, n2810}), .b ({new_AGEMA_signal_1051, n2736}), .clk ( clk ), .r ( Fresh[353] ), .c ({new_AGEMA_signal_1238, n2340}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2514 ( .a ({new_AGEMA_signal_1100, n2348}), .b ({new_AGEMA_signal_1101, n2347}), .clk ( clk ), .r ( Fresh[354] ), .c ({new_AGEMA_signal_1240, n2349}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2517 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_1061, n2690}), .clk ( clk ), .r ( Fresh[355] ), .c ({new_AGEMA_signal_1241, n2375}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2518 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_1051, n2736}), .clk ( clk ), .r ( Fresh[356] ), .c ({new_AGEMA_signal_1242, n2352}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2522 ( .a ({new_AGEMA_signal_1243, n2353}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[357] ), .c ({new_AGEMA_signal_1401, n2354}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2525 ( .a ({new_AGEMA_signal_1004, n2356}), .b ({new_AGEMA_signal_1244, n2355}), .clk ( clk ), .r ( Fresh[358] ), .c ({new_AGEMA_signal_1402, n2357}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2527 ( .a ({new_AGEMA_signal_1147, n2359}), .b ({new_AGEMA_signal_997, n2778}), .clk ( clk ), .r ( Fresh[359] ), .c ({new_AGEMA_signal_1403, n2360}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2534 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ( Fresh[360] ), .c ({new_AGEMA_signal_1540, n2369}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2536 ( .a ({new_AGEMA_signal_1232, n2371}), .b ({new_AGEMA_signal_980, n2713}), .clk ( clk ), .r ( Fresh[361] ), .c ({new_AGEMA_signal_1404, n2372}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2539 ( .a ({new_AGEMA_signal_1087, n2576}), .b ({new_AGEMA_signal_1169, n2376}), .clk ( clk ), .r ( Fresh[362] ), .c ({new_AGEMA_signal_1405, n2377}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2544 ( .a ({new_AGEMA_signal_990, n2609}), .b ({new_AGEMA_signal_1103, n2415}), .clk ( clk ), .r ( Fresh[363] ), .c ({new_AGEMA_signal_1246, n2467}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2545 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_1095, n2383}), .clk ( clk ), .r ( Fresh[364] ), .c ({new_AGEMA_signal_1247, n2385}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2546 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[365] ), .c ({new_AGEMA_signal_1248, n2384}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2548 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1202, n2429}), .clk ( clk ), .r ( Fresh[366] ), .c ({new_AGEMA_signal_1407, n2386}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2552 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1081, n2647}), .clk ( clk ), .r ( Fresh[367] ), .c ({new_AGEMA_signal_1249, n2394}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2553 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[368] ), .c ({new_AGEMA_signal_1250, n2391}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2554 ( .a ({new_AGEMA_signal_1146, n2505}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[369] ), .c ({new_AGEMA_signal_1408, n2390}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2559 ( .a ({new_AGEMA_signal_1006, n2616}), .b ({new_AGEMA_signal_1104, n2700}), .clk ( clk ), .r ( Fresh[370] ), .c ({new_AGEMA_signal_1251, n2396}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2562 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1231, n2438}), .clk ( clk ), .r ( Fresh[371] ), .c ({new_AGEMA_signal_1409, n2406}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2565 ( .a ({new_AGEMA_signal_1105, n2594}), .b ({new_AGEMA_signal_1106, n2402}), .clk ( clk ), .r ( Fresh[372] ), .c ({new_AGEMA_signal_1252, n2403}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2569 ( .a ({new_AGEMA_signal_1178, n2407}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[373] ), .c ({new_AGEMA_signal_1411, n2408}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2573 ( .a ({new_AGEMA_signal_1145, n2412}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ( Fresh[374] ), .c ({new_AGEMA_signal_1412, n2574}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2574 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({new_AGEMA_signal_1007, n2563}), .clk ( clk ), .r ( Fresh[375] ), .c ({new_AGEMA_signal_1253, n2413}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2577 ( .a ({new_AGEMA_signal_1103, n2415}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[376] ), .c ({new_AGEMA_signal_1254, n2416}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2586 ( .a ({new_AGEMA_signal_1255, n2428}), .b ({new_AGEMA_signal_971, n2641}), .clk ( clk ), .r ( Fresh[377] ), .c ({new_AGEMA_signal_1414, n2433}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2587 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_1202, n2429}), .clk ( clk ), .r ( Fresh[378] ), .c ({new_AGEMA_signal_1415, n2689}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2591 ( .a ({new_AGEMA_signal_1081, n2647}), .b ({new_AGEMA_signal_1038, n2492}), .clk ( clk ), .r ( Fresh[379] ), .c ({new_AGEMA_signal_1257, n2434}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2595 ( .a ({new_AGEMA_signal_1231, n2438}), .b ({new_AGEMA_signal_1107, n2483}), .clk ( clk ), .r ( Fresh[380] ), .c ({new_AGEMA_signal_1417, n2439}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2598 ( .a ({new_AGEMA_signal_1050, n2766}), .b ({new_AGEMA_signal_1221, n2540}), .clk ( clk ), .r ( Fresh[381] ), .c ({new_AGEMA_signal_1418, n2445}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2600 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1258, n2443}), .clk ( clk ), .r ( Fresh[382] ), .c ({new_AGEMA_signal_1419, n2444}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2602 ( .a ({new_AGEMA_signal_959, n2790}), .b ({new_AGEMA_signal_1208, n2446}), .clk ( clk ), .r ( Fresh[383] ), .c ({new_AGEMA_signal_1420, n2447}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2607 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1259, n2693}), .clk ( clk ), .r ( Fresh[384] ), .c ({new_AGEMA_signal_1421, n2454}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2617 ( .a ({new_AGEMA_signal_951, n2791}), .b ({new_AGEMA_signal_1109, n2464}), .clk ( clk ), .r ( Fresh[385] ), .c ({new_AGEMA_signal_1260, n2465}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2622 ( .a ({new_AGEMA_signal_953, n2813}), .b ({new_AGEMA_signal_1087, n2576}), .clk ( clk ), .r ( Fresh[386] ), .c ({new_AGEMA_signal_1261, n2470}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2626 ( .a ({new_AGEMA_signal_1111, n2473}), .b ({new_AGEMA_signal_1112, n2472}), .clk ( clk ), .r ( Fresh[387] ), .c ({new_AGEMA_signal_1262, n2476}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2633 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1263, n2480}), .clk ( clk ), .r ( Fresh[388] ), .c ({new_AGEMA_signal_1424, n2481}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2639 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[389] ), .c ({new_AGEMA_signal_1265, n2486}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2642 ( .a ({new_AGEMA_signal_991, n2661}), .b ({new_AGEMA_signal_1114, n2488}), .clk ( clk ), .r ( Fresh[390] ), .c ({new_AGEMA_signal_1266, n2489}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2645 ( .a ({new_AGEMA_signal_992, n2493}), .b ({new_AGEMA_signal_1038, n2492}), .clk ( clk ), .r ( Fresh[391] ), .c ({new_AGEMA_signal_1267, n2497}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2646 ( .a ({new_AGEMA_signal_1037, n2577}), .b ({new_AGEMA_signal_1104, n2700}), .clk ( clk ), .r ( Fresh[392] ), .c ({new_AGEMA_signal_1268, n2495}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2647 ( .a ({new_AGEMA_signal_976, n2780}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ( Fresh[393] ), .c ({new_AGEMA_signal_1426, n2494}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2650 ( .a ({new_AGEMA_signal_1077, n2498}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[394] ), .c ({new_AGEMA_signal_1269, n2499}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2653 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ( Fresh[395] ), .c ({new_AGEMA_signal_1557, n2503}) ) ;
    mux2_GHPC #(.low_latency(0), .pipeline(0)) U2655 ( .s ({new_AGEMA_signal_953, n2813}), .b ({new_AGEMA_signal_1146, n2505}), .a ({new_AGEMA_signal_1056, n2651}), .clk ( clk ), .r ( Fresh[396] ), .c ({new_AGEMA_signal_1427, n2506}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2662 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({SI_s1[1], SI_s0[1]}), .clk ( clk ), .r ( Fresh[397] ), .c ({new_AGEMA_signal_1428, n2518}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2663 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[398] ), .c ({new_AGEMA_signal_1558, n2517}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2666 ( .a ({new_AGEMA_signal_1270, n2520}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[399] ), .c ({new_AGEMA_signal_1429, n2523}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2668 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({new_AGEMA_signal_1115, n2521}), .clk ( clk ), .r ( Fresh[400] ), .c ({new_AGEMA_signal_1430, n2522}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2675 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_1271, n2531}), .clk ( clk ), .r ( Fresh[401] ), .c ({new_AGEMA_signal_1431, n2532}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2677 ( .a ({new_AGEMA_signal_1028, n2769}), .b ({new_AGEMA_signal_1163, n2533}), .clk ( clk ), .r ( Fresh[402] ), .c ({new_AGEMA_signal_1432, n2534}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2681 ( .a ({new_AGEMA_signal_1032, n2541}), .b ({new_AGEMA_signal_1221, n2540}), .clk ( clk ), .r ( Fresh[403] ), .c ({new_AGEMA_signal_1433, n2542}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2683 ( .a ({new_AGEMA_signal_1014, n2545}), .b ({new_AGEMA_signal_1079, n2544}), .clk ( clk ), .r ( Fresh[404] ), .c ({new_AGEMA_signal_1272, n2546}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2687 ( .a ({new_AGEMA_signal_1052, n2673}), .b ({new_AGEMA_signal_1135, n2732}), .clk ( clk ), .r ( Fresh[405] ), .c ({new_AGEMA_signal_1435, n2551}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2690 ( .a ({new_AGEMA_signal_1273, n2553}), .b ({new_AGEMA_signal_1066, n2679}), .clk ( clk ), .r ( Fresh[406] ), .c ({new_AGEMA_signal_1436, n2558}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2692 ( .a ({new_AGEMA_signal_1201, n2555}), .b ({new_AGEMA_signal_1274, n2554}), .clk ( clk ), .r ( Fresh[407] ), .c ({new_AGEMA_signal_1437, n2556}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2696 ( .a ({new_AGEMA_signal_1218, n2561}), .b ({new_AGEMA_signal_1116, n2560}), .clk ( clk ), .r ( Fresh[408] ), .c ({new_AGEMA_signal_1438, n2566}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2697 ( .a ({new_AGEMA_signal_974, n2699}), .b ({new_AGEMA_signal_1186, n2562}), .clk ( clk ), .r ( Fresh[409] ), .c ({new_AGEMA_signal_1439, n2715}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2703 ( .a ({new_AGEMA_signal_1160, n2572}), .b ({new_AGEMA_signal_1055, n2571}), .clk ( clk ), .r ( Fresh[410] ), .c ({new_AGEMA_signal_1440, n2573}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2705 ( .a ({new_AGEMA_signal_1026, n2767}), .b ({new_AGEMA_signal_1173, n2754}), .clk ( clk ), .r ( Fresh[411] ), .c ({new_AGEMA_signal_1441, n2585}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2706 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .r ( Fresh[412] ), .c ({new_AGEMA_signal_1276, n2581}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2707 ( .a ({new_AGEMA_signal_1127, n2575}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[413] ), .c ({new_AGEMA_signal_1442, n2579}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2708 ( .a ({new_AGEMA_signal_1037, n2577}), .b ({new_AGEMA_signal_1087, n2576}), .clk ( clk ), .r ( Fresh[414] ), .c ({new_AGEMA_signal_1277, n2578}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2711 ( .a ({new_AGEMA_signal_1148, n2625}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[415] ), .c ({new_AGEMA_signal_1443, n2582}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2715 ( .a ({new_AGEMA_signal_993, n2587}), .b ({new_AGEMA_signal_1278, n2586}), .clk ( clk ), .r ( Fresh[416] ), .c ({new_AGEMA_signal_1444, n2588}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2719 ( .a ({new_AGEMA_signal_1105, n2594}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[417] ), .c ({new_AGEMA_signal_1279, n2607}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2722 ( .a ({new_AGEMA_signal_1117, n2597}), .b ({new_AGEMA_signal_1280, n2596}), .clk ( clk ), .r ( Fresh[418] ), .c ({new_AGEMA_signal_1445, n2605}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2724 ( .a ({new_AGEMA_signal_1281, n2598}), .b ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .r ( Fresh[419] ), .c ({new_AGEMA_signal_1446, n2603}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2726 ( .a ({new_AGEMA_signal_1021, n2599}), .b ({new_AGEMA_signal_1017, n2777}), .clk ( clk ), .r ( Fresh[420] ), .c ({new_AGEMA_signal_1118, n2601}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2733 ( .a ({new_AGEMA_signal_1283, n2610}), .b ({new_AGEMA_signal_990, n2609}), .clk ( clk ), .r ( Fresh[421] ), .c ({new_AGEMA_signal_1447, n2620}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2736 ( .a ({new_AGEMA_signal_1284, n2614}), .b ({new_AGEMA_signal_1285, n2613}), .clk ( clk ), .r ( Fresh[422] ), .c ({new_AGEMA_signal_1448, n2618}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2743 ( .a ({new_AGEMA_signal_953, n2813}), .b ({new_AGEMA_signal_1148, n2625}), .clk ( clk ), .r ( Fresh[423] ), .c ({new_AGEMA_signal_1449, n2626}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2746 ( .a ({new_AGEMA_signal_1034, n2631}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[424] ), .c ({new_AGEMA_signal_1286, n2632}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2752 ( .a ({new_AGEMA_signal_1287, n2784}), .b ({new_AGEMA_signal_1074, n2642}), .clk ( clk ), .r ( Fresh[425] ), .c ({new_AGEMA_signal_1450, n2644}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2754 ( .a ({SI_s1[4], SI_s0[4]}), .b ({new_AGEMA_signal_1093, n2645}), .clk ( clk ), .r ( Fresh[426] ), .c ({new_AGEMA_signal_1288, n2646}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2758 ( .a ({new_AGEMA_signal_1056, n2651}), .b ({new_AGEMA_signal_1121, n2650}), .clk ( clk ), .r ( Fresh[427] ), .c ({new_AGEMA_signal_1289, n2653}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2760 ( .a ({new_AGEMA_signal_1017, n2777}), .b ({new_AGEMA_signal_1175, n2654}), .clk ( clk ), .r ( Fresh[428] ), .c ({new_AGEMA_signal_1452, n2655}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2764 ( .a ({new_AGEMA_signal_1141, n2662}), .b ({new_AGEMA_signal_991, n2661}), .clk ( clk ), .r ( Fresh[429] ), .c ({new_AGEMA_signal_1453, n2663}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2770 ( .a ({new_AGEMA_signal_1052, n2673}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[430] ), .c ({new_AGEMA_signal_1290, n2675}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2772 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_1043, n2676}), .clk ( clk ), .r ( Fresh[431] ), .c ({new_AGEMA_signal_1291, n2678}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2780 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1027, n2789}), .clk ( clk ), .r ( Fresh[432] ), .c ({new_AGEMA_signal_1292, n2691}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2782 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1259, n2693}), .clk ( clk ), .r ( Fresh[433] ), .c ({new_AGEMA_signal_1455, n2695}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2785 ( .a ({new_AGEMA_signal_1104, n2700}), .b ({new_AGEMA_signal_974, n2699}), .clk ( clk ), .r ( Fresh[434] ), .c ({new_AGEMA_signal_1293, n2701}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2791 ( .a ({new_AGEMA_signal_1294, n2711}), .b ({new_AGEMA_signal_1295, n2710}), .clk ( clk ), .r ( Fresh[435] ), .c ({new_AGEMA_signal_1456, n2717}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2796 ( .a ({new_AGEMA_signal_1323, n2720}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[436] ), .c ({new_AGEMA_signal_1576, n2729}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2798 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1123, n2722}), .clk ( clk ), .r ( Fresh[437] ), .c ({new_AGEMA_signal_1296, n2727}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2803 ( .a ({new_AGEMA_signal_1135, n2732}), .b ({new_AGEMA_signal_1180, n2731}), .clk ( clk ), .r ( Fresh[438] ), .c ({new_AGEMA_signal_1458, n2733}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2807 ( .a ({new_AGEMA_signal_995, n2739}), .b ({new_AGEMA_signal_1298, n2738}), .clk ( clk ), .r ( Fresh[439] ), .c ({new_AGEMA_signal_1459, n2740}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2812 ( .a ({new_AGEMA_signal_1088, n2748}), .b ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[440] ), .c ({new_AGEMA_signal_1299, n2749}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2815 ( .a ({new_AGEMA_signal_1173, n2754}), .b ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .r ( Fresh[441] ), .c ({new_AGEMA_signal_1461, n2757}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2816 ( .a ({new_AGEMA_signal_1030, n2755}), .b ({new_AGEMA_signal_1000, n2772}), .clk ( clk ), .r ( Fresh[442] ), .c ({new_AGEMA_signal_1300, n2756}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2819 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_949, n2760}), .clk ( clk ), .r ( Fresh[443] ), .c ({new_AGEMA_signal_1462, n2762}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2823 ( .a ({new_AGEMA_signal_1028, n2769}), .b ({new_AGEMA_signal_1301, n2768}), .clk ( clk ), .r ( Fresh[444] ), .c ({new_AGEMA_signal_1463, n2770}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2825 ( .a ({new_AGEMA_signal_1184, n2773}), .b ({new_AGEMA_signal_1000, n2772}), .clk ( clk ), .r ( Fresh[445] ), .c ({new_AGEMA_signal_1464, n2776}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2826 ( .a ({new_AGEMA_signal_1228, n2774}), .b ({SI_s1[3], SI_s0[3]}), .clk ( clk ), .r ( Fresh[446] ), .c ({new_AGEMA_signal_1465, n2775}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2830 ( .a ({new_AGEMA_signal_1124, n2782}), .b ({new_AGEMA_signal_1125, n2781}), .clk ( clk ), .r ( Fresh[447] ), .c ({new_AGEMA_signal_1302, n2783}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2836 ( .a ({new_AGEMA_signal_1304, n2794}), .b ({new_AGEMA_signal_1305, n2793}), .clk ( clk ), .r ( Fresh[448] ), .c ({new_AGEMA_signal_1467, n2795}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2845 ( .a ({new_AGEMA_signal_1306, n2812}), .b ({new_AGEMA_signal_1194, n2811}), .clk ( clk ), .r ( Fresh[449] ), .c ({new_AGEMA_signal_1468, n2814}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2848 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_1062, n2817}), .clk ( clk ), .r ( Fresh[450] ), .c ({new_AGEMA_signal_1307, n2819}) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1968 ( .a ({new_AGEMA_signal_1309, n1924}), .b ({new_AGEMA_signal_1310, n1923}), .clk ( clk ), .r ( Fresh[451] ), .c ({new_AGEMA_signal_1470, n1936}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1982 ( .a ({new_AGEMA_signal_1030, n2755}), .b ({new_AGEMA_signal_1311, n1927}), .clk ( clk ), .r ( Fresh[452] ), .c ({new_AGEMA_signal_1471, n1928}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U1994 ( .a ({new_AGEMA_signal_1132, n2151}), .b ({new_AGEMA_signal_1312, n1929}), .clk ( clk ), .r ( Fresh[453] ), .c ({new_AGEMA_signal_1472, n1931}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2012 ( .a ({new_AGEMA_signal_1313, n2665}), .b ({new_AGEMA_signal_1314, n1938}), .clk ( clk ), .r ( Fresh[454] ), .c ({new_AGEMA_signal_1473, n1939}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2024 ( .a ({new_AGEMA_signal_1315, n2235}), .b ({new_AGEMA_signal_1137, n1943}), .clk ( clk ), .r ( Fresh[455] ), .c ({new_AGEMA_signal_1474, n1948}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2032 ( .a ({new_AGEMA_signal_1138, n1946}), .b ({new_AGEMA_signal_1316, n1945}), .clk ( clk ), .r ( Fresh[456] ), .c ({new_AGEMA_signal_1475, n1947}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2041 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_1318, n1951}), .clk ( clk ), .r ( Fresh[457] ), .c ({new_AGEMA_signal_1476, n1954}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2049 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1319, n1952}), .clk ( clk ), .r ( Fresh[458] ), .c ({new_AGEMA_signal_1477, n1953}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2058 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1320, n2687}), .clk ( clk ), .r ( Fresh[459] ), .c ({new_AGEMA_signal_1478, n2658}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2065 ( .a ({new_AGEMA_signal_999, n1964}), .b ({new_AGEMA_signal_1143, n1963}), .clk ( clk ), .r ( Fresh[460] ), .c ({new_AGEMA_signal_1322, n1965}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2078 ( .a ({new_AGEMA_signal_1052, n2673}), .b ({new_AGEMA_signal_1480, n1968}), .clk ( clk ), .r ( Fresh[461] ), .c ({new_AGEMA_signal_1591, n1970}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2084 ( .a ({new_AGEMA_signal_1325, n2684}), .b ({new_AGEMA_signal_1147, n2359}), .clk ( clk ), .r ( Fresh[462] ), .c ({new_AGEMA_signal_1481, n1969}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2093 ( .a ({new_AGEMA_signal_1326, n1972}), .b ({new_AGEMA_signal_1149, n1971}), .clk ( clk ), .r ( Fresh[463] ), .c ({new_AGEMA_signal_1482, n1978}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2102 ( .a ({new_AGEMA_signal_1327, n1974}), .b ({new_AGEMA_signal_1151, n1973}), .clk ( clk ), .r ( Fresh[464] ), .c ({new_AGEMA_signal_1483, n1975}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2107 ( .a ({new_AGEMA_signal_1061, n2690}), .b ({new_AGEMA_signal_1328, n1979}), .clk ( clk ), .r ( Fresh[465] ), .c ({new_AGEMA_signal_1484, n1980}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2114 ( .a ({new_AGEMA_signal_1152, n1985}), .b ({new_AGEMA_signal_1153, n2741}), .clk ( clk ), .r ( Fresh[466] ), .c ({new_AGEMA_signal_1329, n1986}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2124 ( .a ({new_AGEMA_signal_1330, n1994}), .b ({new_AGEMA_signal_1064, n1993}), .clk ( clk ), .r ( Fresh[467] ), .c ({new_AGEMA_signal_1486, n1997}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2137 ( .a ({new_AGEMA_signal_1157, n2241}), .b ({new_AGEMA_signal_1332, n2137}), .clk ( clk ), .r ( Fresh[468] ), .c ({new_AGEMA_signal_1487, n2012}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2145 ( .a ({new_AGEMA_signal_1333, n2006}), .b ({new_AGEMA_signal_1334, n2005}), .clk ( clk ), .r ( Fresh[469] ), .c ({new_AGEMA_signal_1488, n2007}) ) ;
    mux2_GHPC #(.low_latency(0), .pipeline(0)) U2161 ( .s ({new_AGEMA_signal_953, n2813}), .b ({new_AGEMA_signal_1165, n2020}), .a ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ( Fresh[470] ), .c ({new_AGEMA_signal_1336, n2021}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2176 ( .a ({new_AGEMA_signal_1168, n2290}), .b ({new_AGEMA_signal_1338, n2031}), .clk ( clk ), .r ( Fresh[471] ), .c ({new_AGEMA_signal_1490, n2032}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2185 ( .a ({new_AGEMA_signal_1073, n2171}), .b ({new_AGEMA_signal_1339, n2040}), .clk ( clk ), .r ( Fresh[472] ), .c ({new_AGEMA_signal_1491, n2041}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2189 ( .a ({new_AGEMA_signal_1313, n2665}), .b ({new_AGEMA_signal_1172, n2042}), .clk ( clk ), .r ( Fresh[473] ), .c ({new_AGEMA_signal_1492, n2043}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2194 ( .a ({new_AGEMA_signal_1173, n2754}), .b ({new_AGEMA_signal_1340, n2045}), .clk ( clk ), .r ( Fresh[474] ), .c ({new_AGEMA_signal_1493, n2046}) ) ;
    mux2_GHPC #(.low_latency(0), .pipeline(0)) U2204 ( .s ({new_AGEMA_signal_953, n2813}), .b ({new_AGEMA_signal_1342, n2056}), .a ({new_AGEMA_signal_1028, n2769}), .clk ( clk ), .r ( Fresh[475] ), .c ({new_AGEMA_signal_1494, n2058}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2210 ( .a ({new_AGEMA_signal_1150, n2535}), .b ({new_AGEMA_signal_1343, n2060}), .clk ( clk ), .r ( Fresh[476] ), .c ({new_AGEMA_signal_1495, n2063}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2218 ( .a ({new_AGEMA_signal_1344, n2066}), .b ({new_AGEMA_signal_1345, n2065}), .clk ( clk ), .r ( Fresh[477] ), .c ({new_AGEMA_signal_1496, n2652}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2227 ( .a ({new_AGEMA_signal_1074, n2642}), .b ({new_AGEMA_signal_1347, n2074}), .clk ( clk ), .r ( Fresh[478] ), .c ({new_AGEMA_signal_1497, n2076}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2236 ( .a ({new_AGEMA_signal_1011, n2721}), .b ({new_AGEMA_signal_1348, n2082}), .clk ( clk ), .r ( Fresh[479] ), .c ({new_AGEMA_signal_1498, n2105}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2241 ( .a ({new_AGEMA_signal_1184, n2773}), .b ({new_AGEMA_signal_1349, n2084}), .clk ( clk ), .r ( Fresh[480] ), .c ({new_AGEMA_signal_1499, n2099}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2243 ( .a ({new_AGEMA_signal_1350, n2085}), .b ({new_AGEMA_signal_1048, n2627}), .clk ( clk ), .r ( Fresh[481] ), .c ({new_AGEMA_signal_1500, n2091}) ) ;
    and_GHPC #(.low_latency(0), .pipeline(0)) U2246 ( .a ({new_AGEMA_signal_987, n2753}), .b ({new_AGEMA_signal_1351, n2131}), .clk ( clk ), .r ( Fresh[482] ), .c ({new_AGEMA_signal_1501, n2090}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2253 ( .a ({new_AGEMA_signal_1034, n2631}), .b ({new_AGEMA_signal_1353, n2330}), .clk ( clk ), .r ( Fresh[483] ), .c ({new_AGEMA_signal_1502, n2093}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2262 ( .a ({new_AGEMA_signal_1169, n2376}), .b ({new_AGEMA_signal_1356, n2160}), .clk ( clk ), .r ( Fresh[484] ), .c ({new_AGEMA_signal_1503, n2102}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2266 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_1063, n2823}), .clk ( clk ), .r ( Fresh[485] ), .c ({new_AGEMA_signal_1357, n2106}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2272 ( .a ({new_AGEMA_signal_980, n2713}), .b ({new_AGEMA_signal_1504, n2114}), .clk ( clk ), .r ( Fresh[486] ), .c ({new_AGEMA_signal_1606, n2116}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2282 ( .a ({new_AGEMA_signal_1358, n2291}), .b ({new_AGEMA_signal_1192, n2119}), .clk ( clk ), .r ( Fresh[487] ), .c ({new_AGEMA_signal_1505, n2120}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2293 ( .a ({new_AGEMA_signal_1195, n2130}), .b ({new_AGEMA_signal_1196, n2129}), .clk ( clk ), .r ( Fresh[488] ), .c ({new_AGEMA_signal_1359, n2155}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2296 ( .a ({new_AGEMA_signal_994, n2643}), .b ({new_AGEMA_signal_1351, n2131}), .clk ( clk ), .r ( Fresh[489] ), .c ({new_AGEMA_signal_1506, n2543}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2299 ( .a ({new_AGEMA_signal_1198, n2133}), .b ({new_AGEMA_signal_975, n2816}), .clk ( clk ), .r ( Fresh[490] ), .c ({new_AGEMA_signal_1360, n2134}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2303 ( .a ({new_AGEMA_signal_1332, n2137}), .b ({new_AGEMA_signal_1361, n2136}), .clk ( clk ), .r ( Fresh[491] ), .c ({new_AGEMA_signal_1508, n2143}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2308 ( .a ({new_AGEMA_signal_1362, n2139}), .b ({new_AGEMA_signal_1013, n2346}), .clk ( clk ), .r ( Fresh[492] ), .c ({new_AGEMA_signal_1509, n2140}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2324 ( .a ({new_AGEMA_signal_1366, n2157}), .b ({new_AGEMA_signal_1066, n2679}), .clk ( clk ), .r ( Fresh[493] ), .c ({new_AGEMA_signal_1510, n2159}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2326 ( .a ({new_AGEMA_signal_1356, n2160}), .b ({new_AGEMA_signal_1077, n2498}), .clk ( clk ), .r ( Fresh[494] ), .c ({new_AGEMA_signal_1511, n2161}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2330 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_1203, n2163}), .clk ( clk ), .r ( Fresh[495] ), .c ({new_AGEMA_signal_1367, n2164}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2345 ( .a ({new_AGEMA_signal_1085, n2178}), .b ({new_AGEMA_signal_1370, n2177}), .clk ( clk ), .r ( Fresh[496] ), .c ({new_AGEMA_signal_1513, n2179}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2359 ( .a ({new_AGEMA_signal_961, n2315}), .b ({new_AGEMA_signal_1373, n2191}), .clk ( clk ), .r ( Fresh[497] ), .c ({new_AGEMA_signal_1514, n2192}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2370 ( .a ({new_AGEMA_signal_1374, n2201}), .b ({new_AGEMA_signal_1515, n2200}), .clk ( clk ), .r ( Fresh[498] ), .c ({new_AGEMA_signal_1613, n2203}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2382 ( .a ({new_AGEMA_signal_1376, n2217}), .b ({new_AGEMA_signal_1210, n2216}), .clk ( clk ), .r ( Fresh[499] ), .c ({new_AGEMA_signal_1517, n2224}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2388 ( .a ({new_AGEMA_signal_1377, n2222}), .b ({new_AGEMA_signal_1378, n2221}), .clk ( clk ), .r ( Fresh[500] ), .c ({new_AGEMA_signal_1518, n2223}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2392 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_1213, n2226}), .clk ( clk ), .r ( Fresh[501] ), .c ({new_AGEMA_signal_1379, n2229}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2399 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1520, n2233}), .clk ( clk ), .r ( Fresh[502] ), .c ({new_AGEMA_signal_1616, n2234}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2410 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1381, n2244}), .clk ( clk ), .r ( Fresh[503] ), .c ({new_AGEMA_signal_1521, n2246}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2418 ( .a ({new_AGEMA_signal_1146, n2505}), .b ({new_AGEMA_signal_1383, n2253}), .clk ( clk ), .r ( Fresh[504] ), .c ({new_AGEMA_signal_1522, n2254}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2425 ( .a ({new_AGEMA_signal_1221, n2540}), .b ({new_AGEMA_signal_1384, n2260}), .clk ( clk ), .r ( Fresh[505] ), .c ({new_AGEMA_signal_1523, n2263}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2434 ( .a ({new_AGEMA_signal_1092, n2266}), .b ({new_AGEMA_signal_1223, n2265}), .clk ( clk ), .r ( Fresh[506] ), .c ({new_AGEMA_signal_1385, n2267}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2438 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1224, n2269}), .clk ( clk ), .r ( Fresh[507] ), .c ({new_AGEMA_signal_1386, n2270}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2445 ( .a ({new_AGEMA_signal_1225, n2278}), .b ({new_AGEMA_signal_1226, n2277}), .clk ( clk ), .r ( Fresh[508] ), .c ({new_AGEMA_signal_1387, n2279}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2450 ( .a ({new_AGEMA_signal_967, n2779}), .b ({new_AGEMA_signal_1227, n2282}), .clk ( clk ), .r ( Fresh[509] ), .c ({new_AGEMA_signal_1388, n2283}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2453 ( .a ({new_AGEMA_signal_1184, n2773}), .b ({new_AGEMA_signal_1389, n2284}), .clk ( clk ), .r ( Fresh[510] ), .c ({new_AGEMA_signal_1528, n2285}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2457 ( .a ({new_AGEMA_signal_1045, n2442}), .b ({new_AGEMA_signal_1390, n2459}), .clk ( clk ), .r ( Fresh[511] ), .c ({new_AGEMA_signal_1529, n2686}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2460 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1391, n2288}), .clk ( clk ), .r ( Fresh[512] ), .c ({new_AGEMA_signal_1530, n2289}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2463 ( .a ({new_AGEMA_signal_1392, n2458}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[513] ), .c ({new_AGEMA_signal_1531, n2297}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2465 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_1358, n2291}), .clk ( clk ), .r ( Fresh[514] ), .c ({new_AGEMA_signal_1532, n2292}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2473 ( .a ({new_AGEMA_signal_981, n2723}), .b ({new_AGEMA_signal_1394, n2300}), .clk ( clk ), .r ( Fresh[515] ), .c ({new_AGEMA_signal_1533, n2301}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2483 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_1396, n2314}), .clk ( clk ), .r ( Fresh[516] ), .c ({new_AGEMA_signal_1534, n2321}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2487 ( .a ({new_AGEMA_signal_1097, n2319}), .b ({new_AGEMA_signal_1098, n2318}), .clk ( clk ), .r ( Fresh[517] ), .c ({new_AGEMA_signal_1233, n2320}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2493 ( .a ({new_AGEMA_signal_1234, n2326}), .b ({new_AGEMA_signal_1235, n2325}), .clk ( clk ), .r ( Fresh[518] ), .c ({new_AGEMA_signal_1397, n2334}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2497 ( .a ({new_AGEMA_signal_1398, n2329}), .b ({new_AGEMA_signal_967, n2779}), .clk ( clk ), .r ( Fresh[519] ), .c ({new_AGEMA_signal_1535, n2332}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2498 ( .a ({new_AGEMA_signal_1047, n2677}), .b ({new_AGEMA_signal_1353, n2330}), .clk ( clk ), .r ( Fresh[520] ), .c ({new_AGEMA_signal_1536, n2331}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2502 ( .a ({new_AGEMA_signal_1037, n2577}), .b ({new_AGEMA_signal_1537, n2335}), .clk ( clk ), .r ( Fresh[521] ), .c ({new_AGEMA_signal_1626, n2336}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2508 ( .a ({new_AGEMA_signal_1399, n2341}), .b ({new_AGEMA_signal_1238, n2340}), .clk ( clk ), .r ( Fresh[522] ), .c ({new_AGEMA_signal_1538, n2342}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2519 ( .a ({new_AGEMA_signal_1242, n2352}), .b ({new_AGEMA_signal_1005, n2611}), .clk ( clk ), .r ( Fresh[523] ), .c ({new_AGEMA_signal_1400, n2367}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2523 ( .a ({new_AGEMA_signal_1401, n2354}), .b ({new_AGEMA_signal_1053, n2612}), .clk ( clk ), .r ( Fresh[524] ), .c ({new_AGEMA_signal_1539, n2358}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2547 ( .a ({new_AGEMA_signal_1247, n2385}), .b ({new_AGEMA_signal_1248, n2384}), .clk ( clk ), .r ( Fresh[525] ), .c ({new_AGEMA_signal_1406, n2387}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2555 ( .a ({new_AGEMA_signal_1250, n2391}), .b ({new_AGEMA_signal_1408, n2390}), .clk ( clk ), .r ( Fresh[526] ), .c ({new_AGEMA_signal_1542, n2392}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2566 ( .a ({new_AGEMA_signal_1252, n2403}), .b ({SI_s1[6], SI_s0[6]}), .clk ( clk ), .r ( Fresh[527] ), .c ({new_AGEMA_signal_1410, n2404}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2570 ( .a ({new_AGEMA_signal_1150, n2535}), .b ({new_AGEMA_signal_1411, n2408}), .clk ( clk ), .r ( Fresh[528] ), .c ({new_AGEMA_signal_1544, n2409}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2575 ( .a ({new_AGEMA_signal_1412, n2574}), .b ({new_AGEMA_signal_1253, n2413}), .clk ( clk ), .r ( Fresh[529] ), .c ({new_AGEMA_signal_1545, n2414}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2578 ( .a ({new_AGEMA_signal_1148, n2625}), .b ({new_AGEMA_signal_1254, n2416}), .clk ( clk ), .r ( Fresh[530] ), .c ({new_AGEMA_signal_1413, n2418}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2589 ( .a ({new_AGEMA_signal_1415, n2689}), .b ({new_AGEMA_signal_1256, n2431}), .clk ( clk ), .r ( Fresh[531] ), .c ({new_AGEMA_signal_1547, n2432}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2592 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_1257, n2434}), .clk ( clk ), .r ( Fresh[532] ), .c ({new_AGEMA_signal_1416, n2435}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2601 ( .a ({new_AGEMA_signal_1418, n2445}), .b ({new_AGEMA_signal_1419, n2444}), .clk ( clk ), .r ( Fresh[533] ), .c ({new_AGEMA_signal_1548, n2449}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2603 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_1420, n2447}), .clk ( clk ), .r ( Fresh[534] ), .c ({new_AGEMA_signal_1549, n2448}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2609 ( .a ({new_AGEMA_signal_1421, n2454}), .b ({new_AGEMA_signal_1108, n2453}), .clk ( clk ), .r ( Fresh[535] ), .c ({new_AGEMA_signal_1550, n2455}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2612 ( .a ({new_AGEMA_signal_1320, n2687}), .b ({new_AGEMA_signal_1392, n2458}), .clk ( clk ), .r ( Fresh[536] ), .c ({new_AGEMA_signal_1551, n2460}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2618 ( .a ({new_AGEMA_signal_1003, n2624}), .b ({new_AGEMA_signal_1260, n2465}), .clk ( clk ), .r ( Fresh[537] ), .c ({new_AGEMA_signal_1422, n2466}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2629 ( .a ({new_AGEMA_signal_1262, n2476}), .b ({new_AGEMA_signal_1113, n2475}), .clk ( clk ), .r ( Fresh[538] ), .c ({new_AGEMA_signal_1423, n2477}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2634 ( .a ({new_AGEMA_signal_1028, n2769}), .b ({new_AGEMA_signal_1424, n2481}), .clk ( clk ), .r ( Fresh[539] ), .c ({new_AGEMA_signal_1554, n2482}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2640 ( .a ({new_AGEMA_signal_1264, n2487}), .b ({new_AGEMA_signal_1265, n2486}), .clk ( clk ), .r ( Fresh[540] ), .c ({new_AGEMA_signal_1425, n2490}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2648 ( .a ({new_AGEMA_signal_1268, n2495}), .b ({new_AGEMA_signal_1426, n2494}), .clk ( clk ), .r ( Fresh[541] ), .c ({new_AGEMA_signal_1556, n2496}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2654 ( .a ({new_AGEMA_signal_1189, n2504}), .b ({new_AGEMA_signal_1557, n2503}), .clk ( clk ), .r ( Fresh[542] ), .c ({new_AGEMA_signal_1643, n2507}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2664 ( .a ({new_AGEMA_signal_1428, n2518}), .b ({new_AGEMA_signal_1558, n2517}), .clk ( clk ), .r ( Fresh[543] ), .c ({new_AGEMA_signal_1644, n2525}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2669 ( .a ({new_AGEMA_signal_1429, n2523}), .b ({new_AGEMA_signal_1430, n2522}), .clk ( clk ), .r ( Fresh[544] ), .c ({new_AGEMA_signal_1559, n2524}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2676 ( .a ({new_AGEMA_signal_1431, n2532}), .b ({SI_s1[7], SI_s0[7]}), .clk ( clk ), .r ( Fresh[545] ), .c ({new_AGEMA_signal_1560, n2537}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2678 ( .a ({new_AGEMA_signal_1150, n2535}), .b ({new_AGEMA_signal_1432, n2534}), .clk ( clk ), .r ( Fresh[546] ), .c ({new_AGEMA_signal_1561, n2536}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2684 ( .a ({new_AGEMA_signal_1040, n2724}), .b ({new_AGEMA_signal_1272, n2546}), .clk ( clk ), .r ( Fresh[547] ), .c ({new_AGEMA_signal_1434, n2547}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2693 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1437, n2556}), .clk ( clk ), .r ( Fresh[548] ), .c ({new_AGEMA_signal_1562, n2557}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2699 ( .a ({new_AGEMA_signal_1439, n2715}), .b ({new_AGEMA_signal_1275, n2564}), .clk ( clk ), .r ( Fresh[549] ), .c ({new_AGEMA_signal_1563, n2565}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2704 ( .a ({new_AGEMA_signal_1412, n2574}), .b ({new_AGEMA_signal_1440, n2573}), .clk ( clk ), .r ( Fresh[550] ), .c ({new_AGEMA_signal_1564, n2591}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2709 ( .a ({new_AGEMA_signal_1442, n2579}), .b ({new_AGEMA_signal_1277, n2578}), .clk ( clk ), .r ( Fresh[551] ), .c ({new_AGEMA_signal_1565, n2580}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2727 ( .a ({new_AGEMA_signal_1118, n2601}), .b ({new_AGEMA_signal_984, n2600}), .clk ( clk ), .r ( Fresh[552] ), .c ({new_AGEMA_signal_1282, n2602}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2738 ( .a ({new_AGEMA_signal_1448, n2618}), .b ({new_AGEMA_signal_1119, n2617}), .clk ( clk ), .r ( Fresh[553] ), .c ({new_AGEMA_signal_1567, n2619}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2744 ( .a ({new_AGEMA_signal_1048, n2627}), .b ({new_AGEMA_signal_1449, n2626}), .clk ( clk ), .r ( Fresh[554] ), .c ({new_AGEMA_signal_1568, n2628}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2753 ( .a ({new_AGEMA_signal_1450, n2644}), .b ({new_AGEMA_signal_994, n2643}), .clk ( clk ), .r ( Fresh[555] ), .c ({new_AGEMA_signal_1569, n2649}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2755 ( .a ({new_AGEMA_signal_1081, n2647}), .b ({new_AGEMA_signal_1288, n2646}), .clk ( clk ), .r ( Fresh[556] ), .c ({new_AGEMA_signal_1451, n2648}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2765 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1453, n2663}), .clk ( clk ), .r ( Fresh[557] ), .c ({new_AGEMA_signal_1570, n2664}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2771 ( .a ({new_AGEMA_signal_1290, n2675}), .b ({new_AGEMA_signal_1375, n2674}), .clk ( clk ), .r ( Fresh[558] ), .c ({new_AGEMA_signal_1571, n2681}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2773 ( .a ({new_AGEMA_signal_1066, n2679}), .b ({new_AGEMA_signal_1291, n2678}), .clk ( clk ), .r ( Fresh[559] ), .c ({new_AGEMA_signal_1454, n2680}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2776 ( .a ({new_AGEMA_signal_1325, n2684}), .b ({new_AGEMA_signal_1022, n2683}), .clk ( clk ), .r ( Fresh[560] ), .c ({new_AGEMA_signal_1572, n2685}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2778 ( .a ({new_AGEMA_signal_1320, n2687}), .b ({new_AGEMA_signal_1040, n2724}), .clk ( clk ), .r ( Fresh[561] ), .c ({new_AGEMA_signal_1573, n2698}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2779 ( .a ({new_AGEMA_signal_1415, n2689}), .b ({new_AGEMA_signal_1031, n2688}), .clk ( clk ), .r ( Fresh[562] ), .c ({new_AGEMA_signal_1574, n2692}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2793 ( .a ({new_AGEMA_signal_1439, n2715}), .b ({new_AGEMA_signal_1122, n2714}), .clk ( clk ), .r ( Fresh[563] ), .c ({new_AGEMA_signal_1575, n2716}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2800 ( .a ({new_AGEMA_signal_1296, n2727}), .b ({new_AGEMA_signal_1297, n2726}), .clk ( clk ), .r ( Fresh[564] ), .c ({new_AGEMA_signal_1457, n2728}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2804 ( .a ({new_AGEMA_signal_1133, n2734}), .b ({new_AGEMA_signal_1458, n2733}), .clk ( clk ), .r ( Fresh[565] ), .c ({new_AGEMA_signal_1577, n2735}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2808 ( .a ({new_AGEMA_signal_1153, n2741}), .b ({new_AGEMA_signal_1459, n2740}), .clk ( clk ), .r ( Fresh[566] ), .c ({new_AGEMA_signal_1578, n2743}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2813 ( .a ({new_AGEMA_signal_972, n2750}), .b ({new_AGEMA_signal_1299, n2749}), .clk ( clk ), .r ( Fresh[567] ), .c ({new_AGEMA_signal_1460, n2751}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2817 ( .a ({new_AGEMA_signal_1461, n2757}), .b ({new_AGEMA_signal_1300, n2756}), .clk ( clk ), .r ( Fresh[568] ), .c ({new_AGEMA_signal_1579, n2758}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2820 ( .a ({new_AGEMA_signal_1134, n2763}), .b ({new_AGEMA_signal_1462, n2762}), .clk ( clk ), .r ( Fresh[569] ), .c ({new_AGEMA_signal_1580, n2764}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2827 ( .a ({new_AGEMA_signal_1464, n2776}), .b ({new_AGEMA_signal_1465, n2775}), .clk ( clk ), .r ( Fresh[570] ), .c ({new_AGEMA_signal_1581, n2800}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2831 ( .a ({new_AGEMA_signal_1287, n2784}), .b ({new_AGEMA_signal_1302, n2783}), .clk ( clk ), .r ( Fresh[571] ), .c ({new_AGEMA_signal_1466, n2788}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2837 ( .a ({new_AGEMA_signal_943, n2796}), .b ({new_AGEMA_signal_1467, n2795}), .clk ( clk ), .r ( Fresh[572] ), .c ({new_AGEMA_signal_1583, n2797}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2846 ( .a ({new_AGEMA_signal_1468, n2814}), .b ({new_AGEMA_signal_953, n2813}), .clk ( clk ), .r ( Fresh[573] ), .c ({new_AGEMA_signal_1584, n2822}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2849 ( .a ({new_AGEMA_signal_1126, n2820}), .b ({new_AGEMA_signal_1307, n2819}), .clk ( clk ), .r ( Fresh[574] ), .c ({new_AGEMA_signal_1469, n2821}) ) ;

    /* cells in depth 9 */

    /* cells in depth 10 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1983 ( .a ({new_AGEMA_signal_1029, n2707}), .b ({new_AGEMA_signal_1471, n1928}), .clk ( clk ), .r ( Fresh[575] ), .c ({new_AGEMA_signal_1585, n1934}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U1998 ( .a ({new_AGEMA_signal_1472, n1931}), .b ({new_AGEMA_signal_1036, n1930}), .clk ( clk ), .r ( Fresh[576] ), .c ({new_AGEMA_signal_1586, n1932}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2015 ( .a ({new_AGEMA_signal_1473, n1939}), .b ({new_AGEMA_signal_1040, n2724}), .clk ( clk ), .r ( Fresh[577] ), .c ({new_AGEMA_signal_1587, n1940}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2033 ( .a ({new_AGEMA_signal_1474, n1948}), .b ({new_AGEMA_signal_1475, n1947}), .clk ( clk ), .r ( Fresh[578] ), .c ({new_AGEMA_signal_1588, n1961}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2050 ( .a ({new_AGEMA_signal_1476, n1954}), .b ({new_AGEMA_signal_1477, n1953}), .clk ( clk ), .r ( Fresh[579] ), .c ({new_AGEMA_signal_1589, n1955}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2066 ( .a ({new_AGEMA_signal_1321, n1966}), .b ({new_AGEMA_signal_1322, n1965}), .clk ( clk ), .r ( Fresh[580] ), .c ({new_AGEMA_signal_1479, n1967}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2085 ( .a ({new_AGEMA_signal_1591, n1970}), .b ({new_AGEMA_signal_1481, n1969}), .clk ( clk ), .r ( Fresh[581] ), .c ({new_AGEMA_signal_1669, n1984}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2103 ( .a ({new_AGEMA_signal_1060, n1976}), .b ({new_AGEMA_signal_1483, n1975}), .clk ( clk ), .r ( Fresh[582] ), .c ({new_AGEMA_signal_1592, n1977}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2108 ( .a ({SI_s1[1], SI_s0[1]}), .b ({new_AGEMA_signal_1484, n1980}), .clk ( clk ), .r ( Fresh[583] ), .c ({new_AGEMA_signal_1593, n1981}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2115 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_1329, n1986}), .clk ( clk ), .r ( Fresh[584] ), .c ({new_AGEMA_signal_1485, n1987}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2127 ( .a ({new_AGEMA_signal_1486, n1997}), .b ({new_AGEMA_signal_1331, n1996}), .clk ( clk ), .r ( Fresh[585] ), .c ({new_AGEMA_signal_1594, n1998}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2146 ( .a ({new_AGEMA_signal_1159, n2008}), .b ({new_AGEMA_signal_1488, n2007}), .clk ( clk ), .r ( Fresh[586] ), .c ({new_AGEMA_signal_1595, n2010}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2162 ( .a ({new_AGEMA_signal_1164, n2022}), .b ({new_AGEMA_signal_1336, n2021}), .clk ( clk ), .r ( Fresh[587] ), .c ({new_AGEMA_signal_1489, n2024}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2177 ( .a ({new_AGEMA_signal_1337, n2033}), .b ({new_AGEMA_signal_1490, n2032}), .clk ( clk ), .r ( Fresh[588] ), .c ({new_AGEMA_signal_1597, n2035}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2186 ( .a ({new_AGEMA_signal_1491, n2041}), .b ({new_AGEMA_signal_987, n2753}), .clk ( clk ), .r ( Fresh[589] ), .c ({new_AGEMA_signal_1598, n2054}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2190 ( .a ({new_AGEMA_signal_980, n2713}), .b ({new_AGEMA_signal_1492, n2043}), .clk ( clk ), .r ( Fresh[590] ), .c ({new_AGEMA_signal_1599, n2048}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2195 ( .a ({new_AGEMA_signal_1493, n2046}), .b ({new_AGEMA_signal_1023, n2672}), .clk ( clk ), .r ( Fresh[591] ), .c ({new_AGEMA_signal_1600, n2047}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2206 ( .a ({new_AGEMA_signal_1494, n2058}), .b ({new_AGEMA_signal_1177, n2057}), .clk ( clk ), .r ( Fresh[592] ), .c ({new_AGEMA_signal_1601, n2059}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2213 ( .a ({new_AGEMA_signal_1495, n2063}), .b ({new_AGEMA_signal_1179, n2062}), .clk ( clk ), .r ( Fresh[593] ), .c ({new_AGEMA_signal_1602, n2064}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2229 ( .a ({new_AGEMA_signal_1497, n2076}), .b ({new_AGEMA_signal_1075, n2075}), .clk ( clk ), .r ( Fresh[594] ), .c ({new_AGEMA_signal_1603, n2077}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2249 ( .a ({new_AGEMA_signal_1501, n2090}), .b ({new_AGEMA_signal_1352, n2089}), .clk ( clk ), .r ( Fresh[595] ), .c ({new_AGEMA_signal_1604, n2158}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2255 ( .a ({new_AGEMA_signal_1502, n2093}), .b ({new_AGEMA_signal_1354, n2092}), .clk ( clk ), .r ( Fresh[596] ), .c ({new_AGEMA_signal_1605, n2095}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2274 ( .a ({new_AGEMA_signal_1606, n2116}), .b ({new_AGEMA_signal_1190, n2115}), .clk ( clk ), .r ( Fresh[597] ), .c ({new_AGEMA_signal_1681, n2117}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2283 ( .a ({new_AGEMA_signal_1191, n2121}), .b ({new_AGEMA_signal_1505, n2120}), .clk ( clk ), .r ( Fresh[598] ), .c ({new_AGEMA_signal_1607, n2123}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2300 ( .a ({new_AGEMA_signal_1320, n2687}), .b ({new_AGEMA_signal_1360, n2134}), .clk ( clk ), .r ( Fresh[599] ), .c ({new_AGEMA_signal_1507, n2135}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2309 ( .a ({new_AGEMA_signal_1058, n2818}), .b ({new_AGEMA_signal_1509, n2140}), .clk ( clk ), .r ( Fresh[600] ), .c ({new_AGEMA_signal_1609, n2141}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2327 ( .a ({new_AGEMA_signal_1025, n2737}), .b ({new_AGEMA_signal_1511, n2161}), .clk ( clk ), .r ( Fresh[601] ), .c ({new_AGEMA_signal_1610, n2166}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2331 ( .a ({new_AGEMA_signal_978, n2694}), .b ({new_AGEMA_signal_1367, n2164}), .clk ( clk ), .r ( Fresh[602] ), .c ({new_AGEMA_signal_1512, n2165}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2346 ( .a ({new_AGEMA_signal_1513, n2179}), .b ({new_AGEMA_signal_1050, n2766}), .clk ( clk ), .r ( Fresh[603] ), .c ({new_AGEMA_signal_1611, n2180}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2360 ( .a ({new_AGEMA_signal_1372, n2193}), .b ({new_AGEMA_signal_1514, n2192}), .clk ( clk ), .r ( Fresh[604] ), .c ({new_AGEMA_signal_1612, n2194}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2372 ( .a ({new_AGEMA_signal_1613, n2203}), .b ({new_AGEMA_signal_1516, n2202}), .clk ( clk ), .r ( Fresh[605] ), .c ({new_AGEMA_signal_1688, n2204}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2389 ( .a ({new_AGEMA_signal_1517, n2224}), .b ({new_AGEMA_signal_1518, n2223}), .clk ( clk ), .r ( Fresh[606] ), .c ({new_AGEMA_signal_1614, n2225}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2394 ( .a ({new_AGEMA_signal_1379, n2229}), .b ({new_AGEMA_signal_1214, n2228}), .clk ( clk ), .r ( Fresh[607] ), .c ({new_AGEMA_signal_1519, n2230}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2400 ( .a ({new_AGEMA_signal_1315, n2235}), .b ({new_AGEMA_signal_1616, n2234}), .clk ( clk ), .r ( Fresh[608] ), .c ({new_AGEMA_signal_1690, n2236}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2412 ( .a ({new_AGEMA_signal_1521, n2246}), .b ({new_AGEMA_signal_1220, n2245}), .clk ( clk ), .r ( Fresh[609] ), .c ({new_AGEMA_signal_1617, n2247}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2419 ( .a ({new_AGEMA_signal_1522, n2254}), .b ({new_AGEMA_signal_989, n2785}), .clk ( clk ), .r ( Fresh[610] ), .c ({new_AGEMA_signal_1618, n2255}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2427 ( .a ({new_AGEMA_signal_1523, n2263}), .b ({new_AGEMA_signal_1091, n2262}), .clk ( clk ), .r ( Fresh[611] ), .c ({new_AGEMA_signal_1619, n2264}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2435 ( .a ({new_AGEMA_signal_1525, n2752}), .b ({new_AGEMA_signal_1385, n2267}), .clk ( clk ), .r ( Fresh[612] ), .c ({new_AGEMA_signal_1620, n2271}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2446 ( .a ({new_AGEMA_signal_983, n2815}), .b ({new_AGEMA_signal_1387, n2279}), .clk ( clk ), .r ( Fresh[613] ), .c ({new_AGEMA_signal_1526, n2280}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2451 ( .a ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_1388, n2283}), .clk ( clk ), .r ( Fresh[614] ), .c ({new_AGEMA_signal_1527, n2286}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2461 ( .a ({new_AGEMA_signal_1529, n2686}), .b ({new_AGEMA_signal_1530, n2289}), .clk ( clk ), .r ( Fresh[615] ), .c ({new_AGEMA_signal_1622, n2304}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2466 ( .a ({new_AGEMA_signal_1393, n2293}), .b ({new_AGEMA_signal_1532, n2292}), .clk ( clk ), .r ( Fresh[616] ), .c ({new_AGEMA_signal_1623, n2295}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2488 ( .a ({new_AGEMA_signal_1534, n2321}), .b ({new_AGEMA_signal_1233, n2320}), .clk ( clk ), .r ( Fresh[617] ), .c ({new_AGEMA_signal_1624, n2322}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2499 ( .a ({new_AGEMA_signal_1535, n2332}), .b ({new_AGEMA_signal_1536, n2331}), .clk ( clk ), .r ( Fresh[618] ), .c ({new_AGEMA_signal_1625, n2333}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2509 ( .a ({new_AGEMA_signal_1237, n2343}), .b ({new_AGEMA_signal_1538, n2342}), .clk ( clk ), .r ( Fresh[619] ), .c ({new_AGEMA_signal_1627, n2345}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2526 ( .a ({new_AGEMA_signal_1539, n2358}), .b ({new_AGEMA_signal_1402, n2357}), .clk ( clk ), .r ( Fresh[620] ), .c ({new_AGEMA_signal_1628, n2361}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2549 ( .a ({new_AGEMA_signal_1406, n2387}), .b ({new_AGEMA_signal_1407, n2386}), .clk ( clk ), .r ( Fresh[621] ), .c ({new_AGEMA_signal_1541, n2388}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2556 ( .a ({new_AGEMA_signal_949, n2760}), .b ({new_AGEMA_signal_1542, n2392}), .clk ( clk ), .r ( Fresh[622] ), .c ({new_AGEMA_signal_1630, n2393}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2567 ( .a ({new_AGEMA_signal_1027, n2789}), .b ({new_AGEMA_signal_1410, n2404}), .clk ( clk ), .r ( Fresh[623] ), .c ({new_AGEMA_signal_1543, n2405}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2571 ( .a ({new_AGEMA_signal_1544, n2409}), .b ({new_AGEMA_signal_982, n2725}), .clk ( clk ), .r ( Fresh[624] ), .c ({new_AGEMA_signal_1632, n2410}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2576 ( .a ({new_AGEMA_signal_955, n2630}), .b ({new_AGEMA_signal_1545, n2414}), .clk ( clk ), .r ( Fresh[625] ), .c ({new_AGEMA_signal_1633, n2421}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2579 ( .a ({new_AGEMA_signal_1413, n2418}), .b ({new_AGEMA_signal_1324, n2417}), .clk ( clk ), .r ( Fresh[626] ), .c ({new_AGEMA_signal_1546, n2419}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2590 ( .a ({new_AGEMA_signal_1414, n2433}), .b ({new_AGEMA_signal_1547, n2432}), .clk ( clk ), .r ( Fresh[627] ), .c ({new_AGEMA_signal_1635, n2436}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2604 ( .a ({new_AGEMA_signal_1548, n2449}), .b ({new_AGEMA_signal_1549, n2448}), .clk ( clk ), .r ( Fresh[628] ), .c ({new_AGEMA_signal_1636, n2450}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2610 ( .a ({new_AGEMA_signal_1063, n2823}), .b ({new_AGEMA_signal_1550, n2455}), .clk ( clk ), .r ( Fresh[629] ), .c ({new_AGEMA_signal_1637, n2456}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2613 ( .a ({new_AGEMA_signal_1551, n2460}), .b ({new_AGEMA_signal_1390, n2459}), .clk ( clk ), .r ( Fresh[630] ), .c ({new_AGEMA_signal_1638, n2461}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2619 ( .a ({new_AGEMA_signal_1246, n2467}), .b ({new_AGEMA_signal_1422, n2466}), .clk ( clk ), .r ( Fresh[631] ), .c ({new_AGEMA_signal_1552, n2469}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2630 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1423, n2477}), .clk ( clk ), .r ( Fresh[632] ), .c ({new_AGEMA_signal_1553, n2478}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2635 ( .a ({new_AGEMA_signal_1107, n2483}), .b ({new_AGEMA_signal_1554, n2482}), .clk ( clk ), .r ( Fresh[633] ), .c ({new_AGEMA_signal_1640, n2484}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2643 ( .a ({new_AGEMA_signal_1425, n2490}), .b ({new_AGEMA_signal_1266, n2489}), .clk ( clk ), .r ( Fresh[634] ), .c ({new_AGEMA_signal_1555, n2491}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2649 ( .a ({new_AGEMA_signal_1267, n2497}), .b ({new_AGEMA_signal_1556, n2496}), .clk ( clk ), .r ( Fresh[635] ), .c ({new_AGEMA_signal_1642, n2500}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2656 ( .a ({new_AGEMA_signal_1643, n2507}), .b ({new_AGEMA_signal_1427, n2506}), .clk ( clk ), .r ( Fresh[636] ), .c ({new_AGEMA_signal_1708, n2508}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2670 ( .a ({new_AGEMA_signal_1644, n2525}), .b ({new_AGEMA_signal_1559, n2524}), .clk ( clk ), .r ( Fresh[637] ), .c ({new_AGEMA_signal_1709, n2526}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2679 ( .a ({new_AGEMA_signal_1560, n2537}), .b ({new_AGEMA_signal_1561, n2536}), .clk ( clk ), .r ( Fresh[638] ), .c ({new_AGEMA_signal_1645, n2539}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2682 ( .a ({new_AGEMA_signal_1506, n2543}), .b ({new_AGEMA_signal_1433, n2542}), .clk ( clk ), .r ( Fresh[639] ), .c ({new_AGEMA_signal_1646, n2548}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2694 ( .a ({new_AGEMA_signal_1436, n2558}), .b ({new_AGEMA_signal_1562, n2557}), .clk ( clk ), .r ( Fresh[640] ), .c ({new_AGEMA_signal_1647, n2568}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2700 ( .a ({new_AGEMA_signal_1438, n2566}), .b ({new_AGEMA_signal_1563, n2565}), .clk ( clk ), .r ( Fresh[641] ), .c ({new_AGEMA_signal_1648, n2567}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2710 ( .a ({new_AGEMA_signal_1276, n2581}), .b ({new_AGEMA_signal_1565, n2580}), .clk ( clk ), .r ( Fresh[642] ), .c ({new_AGEMA_signal_1649, n2583}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2728 ( .a ({new_AGEMA_signal_1446, n2603}), .b ({new_AGEMA_signal_1282, n2602}), .clk ( clk ), .r ( Fresh[643] ), .c ({new_AGEMA_signal_1566, n2604}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2739 ( .a ({new_AGEMA_signal_1447, n2620}), .b ({new_AGEMA_signal_1567, n2619}), .clk ( clk ), .r ( Fresh[644] ), .c ({new_AGEMA_signal_1651, n2621}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2745 ( .a ({new_AGEMA_signal_1120, n2629}), .b ({new_AGEMA_signal_1568, n2628}), .clk ( clk ), .r ( Fresh[645] ), .c ({new_AGEMA_signal_1652, n2633}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2756 ( .a ({new_AGEMA_signal_1569, n2649}), .b ({new_AGEMA_signal_1451, n2648}), .clk ( clk ), .r ( Fresh[646] ), .c ({new_AGEMA_signal_1653, n2660}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2759 ( .a ({new_AGEMA_signal_1289, n2653}), .b ({new_AGEMA_signal_1496, n2652}), .clk ( clk ), .r ( Fresh[647] ), .c ({new_AGEMA_signal_1654, n2656}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2766 ( .a ({new_AGEMA_signal_1313, n2665}), .b ({new_AGEMA_signal_1570, n2664}), .clk ( clk ), .r ( Fresh[648] ), .c ({new_AGEMA_signal_1655, n2666}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2774 ( .a ({new_AGEMA_signal_1571, n2681}), .b ({new_AGEMA_signal_1454, n2680}), .clk ( clk ), .r ( Fresh[649] ), .c ({new_AGEMA_signal_1656, n2706}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2777 ( .a ({new_AGEMA_signal_1529, n2686}), .b ({new_AGEMA_signal_1572, n2685}), .clk ( clk ), .r ( Fresh[650] ), .c ({new_AGEMA_signal_1657, n2704}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2781 ( .a ({new_AGEMA_signal_1574, n2692}), .b ({new_AGEMA_signal_1292, n2691}), .clk ( clk ), .r ( Fresh[651] ), .c ({new_AGEMA_signal_1658, n2696}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2794 ( .a ({new_AGEMA_signal_1456, n2717}), .b ({new_AGEMA_signal_1575, n2716}), .clk ( clk ), .r ( Fresh[652] ), .c ({new_AGEMA_signal_1659, n2718}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2801 ( .a ({new_AGEMA_signal_1576, n2729}), .b ({new_AGEMA_signal_1457, n2728}), .clk ( clk ), .r ( Fresh[653] ), .c ({new_AGEMA_signal_1660, n2730}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2805 ( .a ({new_AGEMA_signal_1051, n2736}), .b ({new_AGEMA_signal_1577, n2735}), .clk ( clk ), .r ( Fresh[654] ), .c ({new_AGEMA_signal_1661, n2745}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2809 ( .a ({new_AGEMA_signal_1578, n2743}), .b ({new_AGEMA_signal_986, n2742}), .clk ( clk ), .r ( Fresh[655] ), .c ({new_AGEMA_signal_1662, n2744}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2814 ( .a ({new_AGEMA_signal_1525, n2752}), .b ({new_AGEMA_signal_1460, n2751}), .clk ( clk ), .r ( Fresh[656] ), .c ({new_AGEMA_signal_1663, n2759}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2821 ( .a ({new_AGEMA_signal_957, n2765}), .b ({new_AGEMA_signal_1580, n2764}), .clk ( clk ), .r ( Fresh[657] ), .c ({new_AGEMA_signal_1664, n2771}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2833 ( .a ({new_AGEMA_signal_1466, n2788}), .b ({new_AGEMA_signal_1303, n2787}), .clk ( clk ), .r ( Fresh[658] ), .c ({new_AGEMA_signal_1582, n2798}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2850 ( .a ({new_AGEMA_signal_1584, n2822}), .b ({new_AGEMA_signal_1469, n2821}), .clk ( clk ), .r ( Fresh[659] ), .c ({new_AGEMA_signal_1666, n2826}) ) ;

    /* cells in depth 11 */

    /* cells in depth 12 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2001 ( .a ({new_AGEMA_signal_1586, n1932}), .b ({new_AGEMA_signal_1037, n2577}), .clk ( clk ), .r ( Fresh[660] ), .c ({new_AGEMA_signal_1667, n1933}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2051 ( .a ({new_AGEMA_signal_1317, n1956}), .b ({new_AGEMA_signal_1589, n1955}), .clk ( clk ), .r ( Fresh[661] ), .c ({new_AGEMA_signal_1668, n1958}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2067 ( .a ({new_AGEMA_signal_1479, n1967}), .b ({new_AGEMA_signal_963, n2595}), .clk ( clk ), .r ( Fresh[662] ), .c ({new_AGEMA_signal_1590, n1990}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2104 ( .a ({new_AGEMA_signal_1482, n1978}), .b ({new_AGEMA_signal_1592, n1977}), .clk ( clk ), .r ( Fresh[663] ), .c ({new_AGEMA_signal_1670, n1982}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2128 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_1594, n1998}), .clk ( clk ), .r ( Fresh[664] ), .c ({new_AGEMA_signal_1671, n1999}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2148 ( .a ({new_AGEMA_signal_1595, n2010}), .b ({new_AGEMA_signal_1162, n2009}), .clk ( clk ), .r ( Fresh[665] ), .c ({new_AGEMA_signal_1672, n2011}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2165 ( .a ({new_AGEMA_signal_1489, n2024}), .b ({new_AGEMA_signal_1166, n2023}), .clk ( clk ), .r ( Fresh[666] ), .c ({new_AGEMA_signal_1596, n2025}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2179 ( .a ({new_AGEMA_signal_1597, n2035}), .b ({new_AGEMA_signal_1072, n2034}), .clk ( clk ), .r ( Fresh[667] ), .c ({new_AGEMA_signal_1674, n2036}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2196 ( .a ({new_AGEMA_signal_1599, n2048}), .b ({new_AGEMA_signal_1600, n2047}), .clk ( clk ), .r ( Fresh[668] ), .c ({new_AGEMA_signal_1675, n2049}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2207 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1601, n2059}), .clk ( clk ), .r ( Fresh[669] ), .c ({new_AGEMA_signal_1676, n2072}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2214 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1602, n2064}), .clk ( clk ), .r ( Fresh[670] ), .c ({new_AGEMA_signal_1677, n2067}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2230 ( .a ({new_AGEMA_signal_974, n2699}), .b ({new_AGEMA_signal_1603, n2077}), .clk ( clk ), .r ( Fresh[671] ), .c ({new_AGEMA_signal_1678, n2078}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2250 ( .a ({new_AGEMA_signal_1500, n2091}), .b ({new_AGEMA_signal_1604, n2158}), .clk ( clk ), .r ( Fresh[672] ), .c ({new_AGEMA_signal_1679, n2097}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2257 ( .a ({new_AGEMA_signal_1605, n2095}), .b ({new_AGEMA_signal_1355, n2094}), .clk ( clk ), .r ( Fresh[673] ), .c ({new_AGEMA_signal_1680, n2096}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2275 ( .a ({SI_s1[3], SI_s0[3]}), .b ({new_AGEMA_signal_1681, n2117}), .clk ( clk ), .r ( Fresh[674] ), .c ({new_AGEMA_signal_1735, n2128}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2285 ( .a ({new_AGEMA_signal_1607, n2123}), .b ({new_AGEMA_signal_1193, n2122}), .clk ( clk ), .r ( Fresh[675] ), .c ({new_AGEMA_signal_1682, n2124}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2301 ( .a ({new_AGEMA_signal_1506, n2543}), .b ({new_AGEMA_signal_1507, n2135}), .clk ( clk ), .r ( Fresh[676] ), .c ({new_AGEMA_signal_1608, n2148}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2310 ( .a ({new_AGEMA_signal_1199, n2220}), .b ({new_AGEMA_signal_1609, n2141}), .clk ( clk ), .r ( Fresh[677] ), .c ({new_AGEMA_signal_1683, n2142}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2325 ( .a ({new_AGEMA_signal_1510, n2159}), .b ({new_AGEMA_signal_1604, n2158}), .clk ( clk ), .r ( Fresh[678] ), .c ({new_AGEMA_signal_1684, n2168}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2332 ( .a ({new_AGEMA_signal_1610, n2166}), .b ({new_AGEMA_signal_1512, n2165}), .clk ( clk ), .r ( Fresh[679] ), .c ({new_AGEMA_signal_1685, n2167}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2347 ( .a ({new_AGEMA_signal_1369, n2181}), .b ({new_AGEMA_signal_1611, n2180}), .clk ( clk ), .r ( Fresh[680] ), .c ({new_AGEMA_signal_1686, n2184}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2361 ( .a ({new_AGEMA_signal_1371, n2195}), .b ({new_AGEMA_signal_1612, n2194}), .clk ( clk ), .r ( Fresh[681] ), .c ({new_AGEMA_signal_1687, n2197}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2373 ( .a ({new_AGEMA_signal_1063, n2823}), .b ({new_AGEMA_signal_1688, n2204}), .clk ( clk ), .r ( Fresh[682] ), .c ({new_AGEMA_signal_1741, n2205}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2390 ( .a ({new_AGEMA_signal_1065, n2828}), .b ({new_AGEMA_signal_1614, n2225}), .clk ( clk ), .r ( Fresh[683] ), .c ({new_AGEMA_signal_1689, n2232}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2395 ( .a ({new_AGEMA_signal_1519, n2230}), .b ({new_AGEMA_signal_1007, n2563}), .clk ( clk ), .r ( Fresh[684] ), .c ({new_AGEMA_signal_1615, n2231}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2401 ( .a ({new_AGEMA_signal_1215, n2237}), .b ({new_AGEMA_signal_1690, n2236}), .clk ( clk ), .r ( Fresh[685] ), .c ({new_AGEMA_signal_1743, n2239}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2413 ( .a ({new_AGEMA_signal_1380, n2248}), .b ({new_AGEMA_signal_1617, n2247}), .clk ( clk ), .r ( Fresh[686] ), .c ({new_AGEMA_signal_1691, n2250}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2428 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1619, n2264}), .clk ( clk ), .r ( Fresh[687] ), .c ({new_AGEMA_signal_1692, n2276}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2439 ( .a ({new_AGEMA_signal_1620, n2271}), .b ({new_AGEMA_signal_1386, n2270}), .clk ( clk ), .r ( Fresh[688] ), .c ({new_AGEMA_signal_1693, n2272}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2454 ( .a ({new_AGEMA_signal_1527, n2286}), .b ({new_AGEMA_signal_1528, n2285}), .clk ( clk ), .r ( Fresh[689] ), .c ({new_AGEMA_signal_1621, n2306}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2468 ( .a ({new_AGEMA_signal_1623, n2295}), .b ({new_AGEMA_signal_1230, n2294}), .clk ( clk ), .r ( Fresh[690] ), .c ({new_AGEMA_signal_1694, n2296}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2489 ( .a ({new_AGEMA_signal_1395, n2323}), .b ({new_AGEMA_signal_1624, n2322}), .clk ( clk ), .r ( Fresh[691] ), .c ({new_AGEMA_signal_1695, n2324}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2500 ( .a ({new_AGEMA_signal_1397, n2334}), .b ({new_AGEMA_signal_1625, n2333}), .clk ( clk ), .r ( Fresh[692] ), .c ({new_AGEMA_signal_1696, n2337}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2511 ( .a ({new_AGEMA_signal_1627, n2345}), .b ({new_AGEMA_signal_1239, n2344}), .clk ( clk ), .r ( Fresh[693] ), .c ({new_AGEMA_signal_1697, n2350}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2528 ( .a ({new_AGEMA_signal_1628, n2361}), .b ({new_AGEMA_signal_1403, n2360}), .clk ( clk ), .r ( Fresh[694] ), .c ({new_AGEMA_signal_1698, n2362}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2550 ( .a ({new_AGEMA_signal_1246, n2467}), .b ({new_AGEMA_signal_1541, n2388}), .clk ( clk ), .r ( Fresh[695] ), .c ({new_AGEMA_signal_1629, n2389}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2557 ( .a ({new_AGEMA_signal_1249, n2394}), .b ({new_AGEMA_signal_1630, n2393}), .clk ( clk ), .r ( Fresh[696] ), .c ({new_AGEMA_signal_1700, n2397}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2568 ( .a ({new_AGEMA_signal_1409, n2406}), .b ({new_AGEMA_signal_1543, n2405}), .clk ( clk ), .r ( Fresh[697] ), .c ({new_AGEMA_signal_1631, n2411}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2580 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1546, n2419}), .clk ( clk ), .r ( Fresh[698] ), .c ({new_AGEMA_signal_1634, n2420}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2593 ( .a ({new_AGEMA_signal_1635, n2436}), .b ({new_AGEMA_signal_1416, n2435}), .clk ( clk ), .r ( Fresh[699] ), .c ({new_AGEMA_signal_1703, n2440}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2614 ( .a ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1638, n2461}), .clk ( clk ), .r ( Fresh[700] ), .c ({new_AGEMA_signal_1704, n2516}) ) ;
    mux2_GHPC #(.low_latency(0), .pipeline(0)) U2621 ( .s ({SI_s1[2], SI_s0[2]}), .b ({new_AGEMA_signal_1552, n2469}), .a ({new_AGEMA_signal_1110, n2468}), .clk ( clk ), .r ( Fresh[701] ), .c ({new_AGEMA_signal_1639, n2471}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2636 ( .a ({new_AGEMA_signal_1144, n2761}), .b ({new_AGEMA_signal_1640, n2484}), .clk ( clk ), .r ( Fresh[702] ), .c ({new_AGEMA_signal_1706, n2485}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2644 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1555, n2491}), .clk ( clk ), .r ( Fresh[703] ), .c ({new_AGEMA_signal_1641, n2502}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2651 ( .a ({new_AGEMA_signal_1642, n2500}), .b ({new_AGEMA_signal_1269, n2499}), .clk ( clk ), .r ( Fresh[704] ), .c ({new_AGEMA_signal_1707, n2501}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2657 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1708, n2508}), .clk ( clk ), .r ( Fresh[705] ), .c ({new_AGEMA_signal_1757, n2509}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2671 ( .a ({new_AGEMA_signal_989, n2785}), .b ({new_AGEMA_signal_1709, n2526}), .clk ( clk ), .r ( Fresh[706] ), .c ({new_AGEMA_signal_1758, n2527}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2680 ( .a ({new_AGEMA_signal_1645, n2539}), .b ({new_AGEMA_signal_985, n2538}), .clk ( clk ), .r ( Fresh[707] ), .c ({new_AGEMA_signal_1710, n2550}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2685 ( .a ({new_AGEMA_signal_1646, n2548}), .b ({new_AGEMA_signal_1434, n2547}), .clk ( clk ), .r ( Fresh[708] ), .c ({new_AGEMA_signal_1711, n2549}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2701 ( .a ({new_AGEMA_signal_1647, n2568}), .b ({new_AGEMA_signal_1648, n2567}), .clk ( clk ), .r ( Fresh[709] ), .c ({new_AGEMA_signal_1712, n2569}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2712 ( .a ({new_AGEMA_signal_1649, n2583}), .b ({new_AGEMA_signal_1443, n2582}), .clk ( clk ), .r ( Fresh[710] ), .c ({new_AGEMA_signal_1713, n2584}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2729 ( .a ({new_AGEMA_signal_1445, n2605}), .b ({new_AGEMA_signal_1566, n2604}), .clk ( clk ), .r ( Fresh[711] ), .c ({new_AGEMA_signal_1650, n2606}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2740 ( .a ({new_AGEMA_signal_971, n2641}), .b ({new_AGEMA_signal_1651, n2621}), .clk ( clk ), .r ( Fresh[712] ), .c ({new_AGEMA_signal_1715, n2622}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2747 ( .a ({new_AGEMA_signal_1652, n2633}), .b ({new_AGEMA_signal_1286, n2632}), .clk ( clk ), .r ( Fresh[713] ), .c ({new_AGEMA_signal_1716, n2634}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2761 ( .a ({new_AGEMA_signal_1654, n2656}), .b ({new_AGEMA_signal_1452, n2655}), .clk ( clk ), .r ( Fresh[714] ), .c ({new_AGEMA_signal_1717, n2657}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2783 ( .a ({new_AGEMA_signal_1658, n2696}), .b ({new_AGEMA_signal_1455, n2695}), .clk ( clk ), .r ( Fresh[715] ), .c ({new_AGEMA_signal_1718, n2697}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2795 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1659, n2718}), .clk ( clk ), .r ( Fresh[716] ), .c ({new_AGEMA_signal_1719, n2808}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2802 ( .a ({new_AGEMA_signal_1660, n2730}), .b ({new_AGEMA_signal_1067, n2809}), .clk ( clk ), .r ( Fresh[717] ), .c ({new_AGEMA_signal_1720, n2747}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2810 ( .a ({new_AGEMA_signal_1661, n2745}), .b ({new_AGEMA_signal_1662, n2744}), .clk ( clk ), .r ( Fresh[718] ), .c ({new_AGEMA_signal_1721, n2746}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2818 ( .a ({new_AGEMA_signal_1663, n2759}), .b ({new_AGEMA_signal_1579, n2758}), .clk ( clk ), .r ( Fresh[719] ), .c ({new_AGEMA_signal_1722, n2804}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2824 ( .a ({new_AGEMA_signal_1664, n2771}), .b ({new_AGEMA_signal_1463, n2770}), .clk ( clk ), .r ( Fresh[720] ), .c ({new_AGEMA_signal_1723, n2802}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2838 ( .a ({new_AGEMA_signal_1582, n2798}), .b ({new_AGEMA_signal_1583, n2797}), .clk ( clk ), .r ( Fresh[721] ), .c ({new_AGEMA_signal_1665, n2799}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2852 ( .a ({new_AGEMA_signal_1666, n2826}), .b ({new_AGEMA_signal_1308, n2825}), .clk ( clk ), .r ( Fresh[722] ), .c ({new_AGEMA_signal_1725, n2827}) ) ;

    /* cells in depth 13 */

    /* cells in depth 14 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2002 ( .a ({new_AGEMA_signal_1585, n1934}), .b ({new_AGEMA_signal_1667, n1933}), .clk ( clk ), .r ( Fresh[723] ), .c ({new_AGEMA_signal_1726, n1935}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2054 ( .a ({new_AGEMA_signal_1668, n1958}), .b ({new_AGEMA_signal_1049, n1957}), .clk ( clk ), .r ( Fresh[724] ), .c ({new_AGEMA_signal_1727, n1959}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2109 ( .a ({new_AGEMA_signal_1670, n1982}), .b ({new_AGEMA_signal_1593, n1981}), .clk ( clk ), .r ( Fresh[725] ), .c ({new_AGEMA_signal_1728, n1983}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2149 ( .a ({new_AGEMA_signal_1487, n2012}), .b ({new_AGEMA_signal_1672, n2011}), .clk ( clk ), .r ( Fresh[726] ), .c ({new_AGEMA_signal_1729, n2014}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2166 ( .a ({new_AGEMA_signal_1069, n2026}), .b ({new_AGEMA_signal_1596, n2025}), .clk ( clk ), .r ( Fresh[727] ), .c ({new_AGEMA_signal_1673, n2029}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2180 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_1674, n2036}), .clk ( clk ), .r ( Fresh[728] ), .c ({new_AGEMA_signal_1731, n2037}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2197 ( .a ({new_AGEMA_signal_1171, n2050}), .b ({new_AGEMA_signal_1675, n2049}), .clk ( clk ), .r ( Fresh[729] ), .c ({new_AGEMA_signal_1732, n2052}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2219 ( .a ({new_AGEMA_signal_1677, n2067}), .b ({new_AGEMA_signal_1496, n2652}), .clk ( clk ), .r ( Fresh[730] ), .c ({new_AGEMA_signal_1733, n2070}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2258 ( .a ({new_AGEMA_signal_1679, n2097}), .b ({new_AGEMA_signal_1680, n2096}), .clk ( clk ), .r ( Fresh[731] ), .c ({new_AGEMA_signal_1734, n2098}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2287 ( .a ({new_AGEMA_signal_1682, n2124}), .b ({new_AGEMA_signal_1194, n2811}), .clk ( clk ), .r ( Fresh[732] ), .c ({new_AGEMA_signal_1736, n2125}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2311 ( .a ({new_AGEMA_signal_1508, n2143}), .b ({new_AGEMA_signal_1683, n2142}), .clk ( clk ), .r ( Fresh[733] ), .c ({new_AGEMA_signal_1737, n2145}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2333 ( .a ({new_AGEMA_signal_1684, n2168}), .b ({new_AGEMA_signal_1685, n2167}), .clk ( clk ), .r ( Fresh[734] ), .c ({new_AGEMA_signal_1738, n2169}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2350 ( .a ({new_AGEMA_signal_1686, n2184}), .b ({new_AGEMA_signal_1086, n2183}), .clk ( clk ), .r ( Fresh[735] ), .c ({new_AGEMA_signal_1739, n2185}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2365 ( .a ({new_AGEMA_signal_1687, n2197}), .b ({new_AGEMA_signal_1209, n2196}), .clk ( clk ), .r ( Fresh[736] ), .c ({new_AGEMA_signal_1740, n2198}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2396 ( .a ({new_AGEMA_signal_1689, n2232}), .b ({new_AGEMA_signal_1615, n2231}), .clk ( clk ), .r ( Fresh[737] ), .c ({new_AGEMA_signal_1742, n2312}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2404 ( .a ({new_AGEMA_signal_1743, n2239}), .b ({new_AGEMA_signal_1216, n2238}), .clk ( clk ), .r ( Fresh[738] ), .c ({new_AGEMA_signal_1781, n2258}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2415 ( .a ({new_AGEMA_signal_1691, n2250}), .b ({new_AGEMA_signal_1382, n2249}), .clk ( clk ), .r ( Fresh[739] ), .c ({new_AGEMA_signal_1744, n2251}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2440 ( .a ({new_AGEMA_signal_1524, n2273}), .b ({new_AGEMA_signal_1693, n2272}), .clk ( clk ), .r ( Fresh[740] ), .c ({new_AGEMA_signal_1745, n2274}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2469 ( .a ({new_AGEMA_signal_1531, n2297}), .b ({new_AGEMA_signal_1694, n2296}), .clk ( clk ), .r ( Fresh[741] ), .c ({new_AGEMA_signal_1746, n2302}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2490 ( .a ({new_AGEMA_signal_1695, n2324}), .b ({new_AGEMA_signal_1000, n2772}), .clk ( clk ), .r ( Fresh[742] ), .c ({new_AGEMA_signal_1747, n2339}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2503 ( .a ({new_AGEMA_signal_1696, n2337}), .b ({new_AGEMA_signal_1626, n2336}), .clk ( clk ), .r ( Fresh[743] ), .c ({new_AGEMA_signal_1748, n2338}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2515 ( .a ({new_AGEMA_signal_1697, n2350}), .b ({new_AGEMA_signal_1240, n2349}), .clk ( clk ), .r ( Fresh[744] ), .c ({new_AGEMA_signal_1749, n2351}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2529 ( .a ({new_AGEMA_signal_1102, n2363}), .b ({new_AGEMA_signal_1698, n2362}), .clk ( clk ), .r ( Fresh[745] ), .c ({new_AGEMA_signal_1750, n2365}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2551 ( .a ({new_AGEMA_signal_1629, n2389}), .b ({SI_s1[2], SI_s0[2]}), .clk ( clk ), .r ( Fresh[746] ), .c ({new_AGEMA_signal_1699, n2399}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2560 ( .a ({new_AGEMA_signal_1700, n2397}), .b ({new_AGEMA_signal_1251, n2396}), .clk ( clk ), .r ( Fresh[747] ), .c ({new_AGEMA_signal_1751, n2398}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2572 ( .a ({new_AGEMA_signal_1631, n2411}), .b ({new_AGEMA_signal_1632, n2410}), .clk ( clk ), .r ( Fresh[748] ), .c ({new_AGEMA_signal_1701, n2423}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2581 ( .a ({new_AGEMA_signal_1633, n2421}), .b ({new_AGEMA_signal_1634, n2420}), .clk ( clk ), .r ( Fresh[749] ), .c ({new_AGEMA_signal_1702, n2422}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2596 ( .a ({new_AGEMA_signal_1703, n2440}), .b ({new_AGEMA_signal_1417, n2439}), .clk ( clk ), .r ( Fresh[750] ), .c ({new_AGEMA_signal_1753, n2441}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2623 ( .a ({new_AGEMA_signal_1639, n2471}), .b ({new_AGEMA_signal_1261, n2470}), .clk ( clk ), .r ( Fresh[751] ), .c ({new_AGEMA_signal_1705, n2479}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2637 ( .a ({new_AGEMA_signal_1706, n2485}), .b ({new_AGEMA_signal_1026, n2767}), .clk ( clk ), .r ( Fresh[752] ), .c ({new_AGEMA_signal_1755, n2512}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2652 ( .a ({new_AGEMA_signal_1641, n2502}), .b ({new_AGEMA_signal_1707, n2501}), .clk ( clk ), .r ( Fresh[753] ), .c ({new_AGEMA_signal_1756, n2510}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2686 ( .a ({new_AGEMA_signal_1710, n2550}), .b ({new_AGEMA_signal_1711, n2549}), .clk ( clk ), .r ( Fresh[754] ), .c ({new_AGEMA_signal_1759, n2552}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2702 ( .a ({new_AGEMA_signal_1044, n2570}), .b ({new_AGEMA_signal_1712, n2569}), .clk ( clk ), .r ( Fresh[755] ), .c ({new_AGEMA_signal_1760, n2593}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2713 ( .a ({new_AGEMA_signal_1441, n2585}), .b ({new_AGEMA_signal_1713, n2584}), .clk ( clk ), .r ( Fresh[756] ), .c ({new_AGEMA_signal_1761, n2589}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2730 ( .a ({new_AGEMA_signal_1279, n2607}), .b ({new_AGEMA_signal_1650, n2606}), .clk ( clk ), .r ( Fresh[757] ), .c ({new_AGEMA_signal_1714, n2608}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2748 ( .a ({new_AGEMA_signal_958, n2635}), .b ({new_AGEMA_signal_1716, n2634}), .clk ( clk ), .r ( Fresh[758] ), .c ({new_AGEMA_signal_1763, n2636}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2762 ( .a ({new_AGEMA_signal_1478, n2658}), .b ({new_AGEMA_signal_1717, n2657}), .clk ( clk ), .r ( Fresh[759] ), .c ({new_AGEMA_signal_1764, n2659}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2784 ( .a ({new_AGEMA_signal_1573, n2698}), .b ({new_AGEMA_signal_1718, n2697}), .clk ( clk ), .r ( Fresh[760] ), .c ({new_AGEMA_signal_1765, n2702}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2811 ( .a ({new_AGEMA_signal_1720, n2747}), .b ({new_AGEMA_signal_1721, n2746}), .clk ( clk ), .r ( Fresh[761] ), .c ({new_AGEMA_signal_1766, n2806}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2839 ( .a ({new_AGEMA_signal_1581, n2800}), .b ({new_AGEMA_signal_1665, n2799}), .clk ( clk ), .r ( Fresh[762] ), .c ({new_AGEMA_signal_1724, n2801}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2853 ( .a ({new_AGEMA_signal_1065, n2828}), .b ({new_AGEMA_signal_1725, n2827}), .clk ( clk ), .r ( Fresh[763] ), .c ({new_AGEMA_signal_1768, n2829}) ) ;

    /* cells in depth 15 */

    /* cells in depth 16 */
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2003 ( .a ({new_AGEMA_signal_1470, n1936}), .b ({new_AGEMA_signal_1726, n1935}), .clk ( clk ), .r ( Fresh[764] ), .c ({new_AGEMA_signal_1769, n1941}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2059 ( .a ({new_AGEMA_signal_1727, n1959}), .b ({new_AGEMA_signal_1478, n2658}), .clk ( clk ), .r ( Fresh[765] ), .c ({new_AGEMA_signal_1770, n1960}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2110 ( .a ({new_AGEMA_signal_1669, n1984}), .b ({new_AGEMA_signal_1728, n1983}), .clk ( clk ), .r ( Fresh[766] ), .c ({new_AGEMA_signal_1771, n1988}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2153 ( .a ({new_AGEMA_signal_1729, n2014}), .b ({new_AGEMA_signal_1335, n2013}), .clk ( clk ), .r ( Fresh[767] ), .c ({new_AGEMA_signal_1772, n2015}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2169 ( .a ({new_AGEMA_signal_1673, n2029}), .b ({new_AGEMA_signal_1071, n2028}), .clk ( clk ), .r ( Fresh[768] ), .c ({new_AGEMA_signal_1730, n2030}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2200 ( .a ({new_AGEMA_signal_1732, n2052}), .b ({new_AGEMA_signal_1341, n2051}), .clk ( clk ), .r ( Fresh[769] ), .c ({new_AGEMA_signal_1774, n2053}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2222 ( .a ({new_AGEMA_signal_1733, n2070}), .b ({new_AGEMA_signal_1346, n2069}), .clk ( clk ), .r ( Fresh[770] ), .c ({new_AGEMA_signal_1775, n2071}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2259 ( .a ({new_AGEMA_signal_1499, n2099}), .b ({new_AGEMA_signal_1734, n2098}), .clk ( clk ), .r ( Fresh[771] ), .c ({new_AGEMA_signal_1776, n2103}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2288 ( .a ({new_AGEMA_signal_1079, n2544}), .b ({new_AGEMA_signal_1736, n2125}), .clk ( clk ), .r ( Fresh[772] ), .c ({new_AGEMA_signal_1777, n2126}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2314 ( .a ({new_AGEMA_signal_1737, n2145}), .b ({new_AGEMA_signal_1363, n2144}), .clk ( clk ), .r ( Fresh[773] ), .c ({new_AGEMA_signal_1778, n2146}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2334 ( .a ({new_AGEMA_signal_1365, n2170}), .b ({new_AGEMA_signal_1738, n2169}), .clk ( clk ), .r ( Fresh[774] ), .c ({new_AGEMA_signal_1779, n2173}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2351 ( .a ({new_AGEMA_signal_1084, n2186}), .b ({new_AGEMA_signal_1739, n2185}), .clk ( clk ), .r ( Fresh[775] ), .c ({new_AGEMA_signal_1780, n2187}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2416 ( .a ({new_AGEMA_signal_996, n2437}), .b ({new_AGEMA_signal_1744, n2251}), .clk ( clk ), .r ( Fresh[776] ), .c ({new_AGEMA_signal_1782, n2256}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2441 ( .a ({new_AGEMA_signal_1745, n2274}), .b ({SI_s1[0], SI_s0[0]}), .clk ( clk ), .r ( Fresh[777] ), .c ({new_AGEMA_signal_1783, n2275}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2474 ( .a ({new_AGEMA_signal_1746, n2302}), .b ({new_AGEMA_signal_1533, n2301}), .clk ( clk ), .r ( Fresh[778] ), .c ({new_AGEMA_signal_1784, n2303}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2504 ( .a ({new_AGEMA_signal_1747, n2339}), .b ({new_AGEMA_signal_1748, n2338}), .clk ( clk ), .r ( Fresh[779] ), .c ({new_AGEMA_signal_1785, n2382}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2516 ( .a ({new_AGEMA_signal_1749, n2351}), .b ({new_AGEMA_signal_971, n2641}), .clk ( clk ), .r ( Fresh[780] ), .c ({new_AGEMA_signal_1786, n2380}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2531 ( .a ({new_AGEMA_signal_1750, n2365}), .b ({new_AGEMA_signal_1245, n2364}), .clk ( clk ), .r ( Fresh[781] ), .c ({new_AGEMA_signal_1787, n2366}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2561 ( .a ({new_AGEMA_signal_1699, n2399}), .b ({new_AGEMA_signal_1751, n2398}), .clk ( clk ), .r ( Fresh[782] ), .c ({new_AGEMA_signal_1788, n2425}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2582 ( .a ({new_AGEMA_signal_1701, n2423}), .b ({new_AGEMA_signal_1702, n2422}), .clk ( clk ), .r ( Fresh[783] ), .c ({new_AGEMA_signal_1752, n2424}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2597 ( .a ({new_AGEMA_signal_1031, n2688}), .b ({new_AGEMA_signal_1753, n2441}), .clk ( clk ), .r ( Fresh[784] ), .c ({new_AGEMA_signal_1789, n2451}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2631 ( .a ({new_AGEMA_signal_1705, n2479}), .b ({new_AGEMA_signal_1553, n2478}), .clk ( clk ), .r ( Fresh[785] ), .c ({new_AGEMA_signal_1754, n2514}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2658 ( .a ({new_AGEMA_signal_1756, n2510}), .b ({new_AGEMA_signal_1757, n2509}), .clk ( clk ), .r ( Fresh[786] ), .c ({new_AGEMA_signal_1790, n2511}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2688 ( .a ({new_AGEMA_signal_1759, n2552}), .b ({new_AGEMA_signal_1435, n2551}), .clk ( clk ), .r ( Fresh[787] ), .c ({new_AGEMA_signal_1791, n2671}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2716 ( .a ({new_AGEMA_signal_1761, n2589}), .b ({new_AGEMA_signal_1444, n2588}), .clk ( clk ), .r ( Fresh[788] ), .c ({new_AGEMA_signal_1792, n2590}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2731 ( .a ({new_AGEMA_signal_1714, n2608}), .b ({new_AGEMA_signal_1050, n2766}), .clk ( clk ), .r ( Fresh[789] ), .c ({new_AGEMA_signal_1762, n2623}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2763 ( .a ({new_AGEMA_signal_1653, n2660}), .b ({new_AGEMA_signal_1764, n2659}), .clk ( clk ), .r ( Fresh[790] ), .c ({new_AGEMA_signal_1794, n2667}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2786 ( .a ({new_AGEMA_signal_1765, n2702}), .b ({new_AGEMA_signal_1293, n2701}), .clk ( clk ), .r ( Fresh[791] ), .c ({new_AGEMA_signal_1795, n2703}) ) ;
    mux2_GHPC #(.low_latency(0), .pipeline(0)) U2840 ( .s ({SI_s1[0], SI_s0[0]}), .b ({new_AGEMA_signal_1723, n2802}), .a ({new_AGEMA_signal_1724, n2801}), .clk ( clk ), .r ( Fresh[792] ), .c ({new_AGEMA_signal_1767, n2803}) ) ;

    /* cells in depth 17 */

    /* cells in depth 18 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2016 ( .a ({new_AGEMA_signal_1769, n1941}), .b ({new_AGEMA_signal_1587, n1940}), .clk ( clk ), .r ( Fresh[793] ), .c ({new_AGEMA_signal_1797, n2019}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2060 ( .a ({new_AGEMA_signal_1588, n1961}), .b ({new_AGEMA_signal_1770, n1960}), .clk ( clk ), .r ( Fresh[794] ), .c ({new_AGEMA_signal_1798, n2002}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2116 ( .a ({new_AGEMA_signal_1771, n1988}), .b ({new_AGEMA_signal_1485, n1987}), .clk ( clk ), .r ( Fresh[795] ), .c ({new_AGEMA_signal_1799, n1989}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2154 ( .a ({new_AGEMA_signal_1065, n2828}), .b ({new_AGEMA_signal_1772, n2015}), .clk ( clk ), .r ( Fresh[796] ), .c ({new_AGEMA_signal_1800, n2016}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2170 ( .a ({new_AGEMA_signal_986, n2742}), .b ({new_AGEMA_signal_1730, n2030}), .clk ( clk ), .r ( Fresh[797] ), .c ({new_AGEMA_signal_1773, n2038}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2201 ( .a ({new_AGEMA_signal_1598, n2054}), .b ({new_AGEMA_signal_1774, n2053}), .clk ( clk ), .r ( Fresh[798] ), .c ({new_AGEMA_signal_1802, n2111}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2223 ( .a ({new_AGEMA_signal_1676, n2072}), .b ({new_AGEMA_signal_1775, n2071}), .clk ( clk ), .r ( Fresh[799] ), .c ({new_AGEMA_signal_1803, n2079}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2263 ( .a ({new_AGEMA_signal_1776, n2103}), .b ({new_AGEMA_signal_1503, n2102}), .clk ( clk ), .r ( Fresh[800] ), .c ({new_AGEMA_signal_1804, n2104}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2289 ( .a ({new_AGEMA_signal_1023, n2672}), .b ({new_AGEMA_signal_1777, n2126}), .clk ( clk ), .r ( Fresh[801] ), .c ({new_AGEMA_signal_1805, n2127}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2315 ( .a ({new_AGEMA_signal_1065, n2828}), .b ({new_AGEMA_signal_1778, n2146}), .clk ( clk ), .r ( Fresh[802] ), .c ({new_AGEMA_signal_1806, n2147}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2336 ( .a ({new_AGEMA_signal_1779, n2173}), .b ({new_AGEMA_signal_1368, n2172}), .clk ( clk ), .r ( Fresh[803] ), .c ({new_AGEMA_signal_1807, n2208}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2352 ( .a ({new_AGEMA_signal_1780, n2187}), .b ({new_AGEMA_signal_955, n2630}), .clk ( clk ), .r ( Fresh[804] ), .c ({new_AGEMA_signal_1808, n2199}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2420 ( .a ({new_AGEMA_signal_1782, n2256}), .b ({new_AGEMA_signal_1618, n2255}), .clk ( clk ), .r ( Fresh[805] ), .c ({new_AGEMA_signal_1809, n2257}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2442 ( .a ({new_AGEMA_signal_1692, n2276}), .b ({new_AGEMA_signal_1783, n2275}), .clk ( clk ), .r ( Fresh[806] ), .c ({new_AGEMA_signal_1810, n2281}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2475 ( .a ({new_AGEMA_signal_1622, n2304}), .b ({new_AGEMA_signal_1784, n2303}), .clk ( clk ), .r ( Fresh[807] ), .c ({new_AGEMA_signal_1811, n2305}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2532 ( .a ({new_AGEMA_signal_1400, n2367}), .b ({new_AGEMA_signal_1787, n2366}), .clk ( clk ), .r ( Fresh[808] ), .c ({new_AGEMA_signal_1812, n2368}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2583 ( .a ({new_AGEMA_signal_1788, n2425}), .b ({new_AGEMA_signal_1752, n2424}), .clk ( clk ), .r ( Fresh[809] ), .c ({new_AGEMA_signal_1813, n2426}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2605 ( .a ({new_AGEMA_signal_1789, n2451}), .b ({new_AGEMA_signal_1636, n2450}), .clk ( clk ), .r ( Fresh[810] ), .c ({new_AGEMA_signal_1814, n2457}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2659 ( .a ({new_AGEMA_signal_1755, n2512}), .b ({new_AGEMA_signal_1790, n2511}), .clk ( clk ), .r ( Fresh[811] ), .c ({new_AGEMA_signal_1815, n2513}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2717 ( .a ({new_AGEMA_signal_1564, n2591}), .b ({new_AGEMA_signal_1792, n2590}), .clk ( clk ), .r ( Fresh[812] ), .c ({new_AGEMA_signal_1816, n2592}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2741 ( .a ({new_AGEMA_signal_1762, n2623}), .b ({new_AGEMA_signal_1715, n2622}), .clk ( clk ), .r ( Fresh[813] ), .c ({new_AGEMA_signal_1793, n2637}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2767 ( .a ({new_AGEMA_signal_1794, n2667}), .b ({new_AGEMA_signal_1655, n2666}), .clk ( clk ), .r ( Fresh[814] ), .c ({new_AGEMA_signal_1818, n2668}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2787 ( .a ({new_AGEMA_signal_1657, n2704}), .b ({new_AGEMA_signal_1795, n2703}), .clk ( clk ), .r ( Fresh[815] ), .c ({new_AGEMA_signal_1819, n2705}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2841 ( .a ({new_AGEMA_signal_1722, n2804}), .b ({new_AGEMA_signal_1767, n2803}), .clk ( clk ), .r ( Fresh[816] ), .c ({new_AGEMA_signal_1796, n2805}) ) ;

    /* cells in depth 19 */

    /* cells in depth 20 */
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2117 ( .a ({new_AGEMA_signal_1590, n1990}), .b ({new_AGEMA_signal_1799, n1989}), .clk ( clk ), .r ( Fresh[817] ), .c ({new_AGEMA_signal_1821, n2000}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2181 ( .a ({new_AGEMA_signal_1773, n2038}), .b ({new_AGEMA_signal_1731, n2037}), .clk ( clk ), .r ( Fresh[818] ), .c ({new_AGEMA_signal_1801, n2113}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2231 ( .a ({new_AGEMA_signal_1803, n2079}), .b ({new_AGEMA_signal_1678, n2078}), .clk ( clk ), .r ( Fresh[819] ), .c ({new_AGEMA_signal_1822, n2109}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2264 ( .a ({new_AGEMA_signal_1498, n2105}), .b ({new_AGEMA_signal_1804, n2104}), .clk ( clk ), .r ( Fresh[820] ), .c ({new_AGEMA_signal_1823, n2107}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2290 ( .a ({new_AGEMA_signal_1735, n2128}), .b ({new_AGEMA_signal_1805, n2127}), .clk ( clk ), .r ( Fresh[821] ), .c ({new_AGEMA_signal_1824, n2212}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2316 ( .a ({new_AGEMA_signal_1608, n2148}), .b ({new_AGEMA_signal_1806, n2147}), .clk ( clk ), .r ( Fresh[822] ), .c ({new_AGEMA_signal_1825, n2149}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2366 ( .a ({new_AGEMA_signal_1808, n2199}), .b ({new_AGEMA_signal_1740, n2198}), .clk ( clk ), .r ( Fresh[823] ), .c ({new_AGEMA_signal_1826, n2206}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2421 ( .a ({new_AGEMA_signal_1781, n2258}), .b ({new_AGEMA_signal_1809, n2257}), .clk ( clk ), .r ( Fresh[824] ), .c ({new_AGEMA_signal_1827, n2310}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2447 ( .a ({new_AGEMA_signal_1810, n2281}), .b ({new_AGEMA_signal_1526, n2280}), .clk ( clk ), .r ( Fresh[825] ), .c ({new_AGEMA_signal_1828, n2308}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2476 ( .a ({new_AGEMA_signal_1621, n2306}), .b ({new_AGEMA_signal_1811, n2305}), .clk ( clk ), .r ( Fresh[826] ), .c ({new_AGEMA_signal_1829, n2307}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2533 ( .a ({new_AGEMA_signal_970, n2719}), .b ({new_AGEMA_signal_1812, n2368}), .clk ( clk ), .r ( Fresh[827] ), .c ({new_AGEMA_signal_1830, n2370}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2611 ( .a ({new_AGEMA_signal_1814, n2457}), .b ({new_AGEMA_signal_1637, n2456}), .clk ( clk ), .r ( Fresh[828] ), .c ({new_AGEMA_signal_1831, n2530}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2660 ( .a ({new_AGEMA_signal_1754, n2514}), .b ({new_AGEMA_signal_1815, n2513}), .clk ( clk ), .r ( Fresh[829] ), .c ({new_AGEMA_signal_1832, n2515}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2718 ( .a ({new_AGEMA_signal_1760, n2593}), .b ({new_AGEMA_signal_1816, n2592}), .clk ( clk ), .r ( Fresh[830] ), .c ({new_AGEMA_signal_1833, n2639}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2749 ( .a ({new_AGEMA_signal_1793, n2637}), .b ({new_AGEMA_signal_1763, n2636}), .clk ( clk ), .r ( Fresh[831] ), .c ({new_AGEMA_signal_1817, n2638}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2788 ( .a ({new_AGEMA_signal_1656, n2706}), .b ({new_AGEMA_signal_1819, n2705}), .clk ( clk ), .r ( Fresh[832] ), .c ({new_AGEMA_signal_1834, n2832}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2842 ( .a ({new_AGEMA_signal_1766, n2806}), .b ({new_AGEMA_signal_1796, n2805}), .clk ( clk ), .r ( Fresh[833] ), .c ({new_AGEMA_signal_1820, n2807}) ) ;

    /* cells in depth 21 */

    /* cells in depth 22 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2129 ( .a ({new_AGEMA_signal_1821, n2000}), .b ({new_AGEMA_signal_1671, n1999}), .clk ( clk ), .r ( Fresh[834] ), .c ({new_AGEMA_signal_1836, n2001}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2267 ( .a ({new_AGEMA_signal_1823, n2107}), .b ({new_AGEMA_signal_1357, n2106}), .clk ( clk ), .r ( Fresh[835] ), .c ({new_AGEMA_signal_1837, n2108}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2317 ( .a ({new_AGEMA_signal_1197, n2150}), .b ({new_AGEMA_signal_1825, n2149}), .clk ( clk ), .r ( Fresh[836] ), .c ({new_AGEMA_signal_1838, n2153}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2374 ( .a ({new_AGEMA_signal_1826, n2206}), .b ({new_AGEMA_signal_1741, n2205}), .clk ( clk ), .r ( Fresh[837] ), .c ({new_AGEMA_signal_1839, n2207}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2477 ( .a ({new_AGEMA_signal_1828, n2308}), .b ({new_AGEMA_signal_1829, n2307}), .clk ( clk ), .r ( Fresh[838] ), .c ({new_AGEMA_signal_1840, n2309}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2535 ( .a ({new_AGEMA_signal_1830, n2370}), .b ({new_AGEMA_signal_1540, n2369}), .clk ( clk ), .r ( Fresh[839] ), .c ({new_AGEMA_signal_1841, n2373}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2661 ( .a ({new_AGEMA_signal_1704, n2516}), .b ({new_AGEMA_signal_1832, n2515}), .clk ( clk ), .r ( Fresh[840] ), .c ({new_AGEMA_signal_1842, n2528}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2750 ( .a ({new_AGEMA_signal_1833, n2639}), .b ({new_AGEMA_signal_1817, n2638}), .clk ( clk ), .r ( Fresh[841] ), .c ({new_AGEMA_signal_1843, n2669}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2843 ( .a ({new_AGEMA_signal_1719, n2808}), .b ({new_AGEMA_signal_1820, n2807}), .clk ( clk ), .r ( Fresh[842] ), .c ({new_AGEMA_signal_1835, n2830}) ) ;

    /* cells in depth 23 */

    /* cells in depth 24 */
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2130 ( .a ({new_AGEMA_signal_1798, n2002}), .b ({new_AGEMA_signal_1836, n2001}), .clk ( clk ), .r ( Fresh[843] ), .c ({new_AGEMA_signal_1845, n2017}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2268 ( .a ({new_AGEMA_signal_1822, n2109}), .b ({new_AGEMA_signal_1837, n2108}), .clk ( clk ), .r ( Fresh[844] ), .c ({new_AGEMA_signal_1846, n2110}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2319 ( .a ({new_AGEMA_signal_1838, n2153}), .b ({new_AGEMA_signal_1364, n2152}), .clk ( clk ), .r ( Fresh[845] ), .c ({new_AGEMA_signal_1847, n2154}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2375 ( .a ({new_AGEMA_signal_1807, n2208}), .b ({new_AGEMA_signal_1839, n2207}), .clk ( clk ), .r ( Fresh[846] ), .c ({new_AGEMA_signal_1848, n2209}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2478 ( .a ({new_AGEMA_signal_1827, n2310}), .b ({new_AGEMA_signal_1840, n2309}), .clk ( clk ), .r ( Fresh[847] ), .c ({new_AGEMA_signal_1849, n2311}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2537 ( .a ({new_AGEMA_signal_1841, n2373}), .b ({new_AGEMA_signal_1404, n2372}), .clk ( clk ), .r ( Fresh[848] ), .c ({new_AGEMA_signal_1850, n2374}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2672 ( .a ({new_AGEMA_signal_1842, n2528}), .b ({new_AGEMA_signal_1758, n2527}), .clk ( clk ), .r ( Fresh[849] ), .c ({new_AGEMA_signal_1851, n2529}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2768 ( .a ({new_AGEMA_signal_1843, n2669}), .b ({new_AGEMA_signal_1818, n2668}), .clk ( clk ), .r ( Fresh[850] ), .c ({new_AGEMA_signal_1852, n2670}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2854 ( .a ({new_AGEMA_signal_1835, n2830}), .b ({new_AGEMA_signal_1768, n2829}), .clk ( clk ), .r ( Fresh[851] ), .c ({new_AGEMA_signal_1844, n2831}) ) ;

    /* cells in depth 25 */

    /* cells in depth 26 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2155 ( .a ({new_AGEMA_signal_1845, n2017}), .b ({new_AGEMA_signal_1800, n2016}), .clk ( clk ), .r ( Fresh[852] ), .c ({new_AGEMA_signal_1854, n2018}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2269 ( .a ({new_AGEMA_signal_1802, n2111}), .b ({new_AGEMA_signal_1846, n2110}), .clk ( clk ), .r ( Fresh[853] ), .c ({new_AGEMA_signal_1855, n2112}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2320 ( .a ({new_AGEMA_signal_1359, n2155}), .b ({new_AGEMA_signal_1847, n2154}), .clk ( clk ), .r ( Fresh[854] ), .c ({new_AGEMA_signal_1856, n2210}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2479 ( .a ({new_AGEMA_signal_1742, n2312}), .b ({new_AGEMA_signal_1849, n2311}), .clk ( clk ), .r ( Fresh[855] ), .c ({new_AGEMA_signal_1857, N470}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2538 ( .a ({new_AGEMA_signal_1241, n2375}), .b ({new_AGEMA_signal_1850, n2374}), .clk ( clk ), .r ( Fresh[856] ), .c ({new_AGEMA_signal_1858, n2378}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2673 ( .a ({new_AGEMA_signal_1831, n2530}), .b ({new_AGEMA_signal_1851, n2529}), .clk ( clk ), .r ( Fresh[857] ), .c ({new_AGEMA_signal_1859, N639}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2769 ( .a ({new_AGEMA_signal_1791, n2671}), .b ({new_AGEMA_signal_1852, n2670}), .clk ( clk ), .r ( Fresh[858] ), .c ({new_AGEMA_signal_1860, N723}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2855 ( .a ({new_AGEMA_signal_1834, n2832}), .b ({new_AGEMA_signal_1844, n2831}), .clk ( clk ), .r ( Fresh[859] ), .c ({new_AGEMA_signal_1853, N789}) ) ;

    /* cells in depth 27 */

    /* cells in depth 28 */
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2156 ( .a ({new_AGEMA_signal_1797, n2019}), .b ({new_AGEMA_signal_1854, n2018}), .clk ( clk ), .r ( Fresh[860] ), .c ({new_AGEMA_signal_1861, N169}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2270 ( .a ({new_AGEMA_signal_1801, n2113}), .b ({new_AGEMA_signal_1855, n2112}), .clk ( clk ), .r ( Fresh[861] ), .c ({new_AGEMA_signal_1862, N277}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2376 ( .a ({new_AGEMA_signal_1856, n2210}), .b ({new_AGEMA_signal_1848, n2209}), .clk ( clk ), .r ( Fresh[862] ), .c ({new_AGEMA_signal_1863, n2211}) ) ;
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2540 ( .a ({new_AGEMA_signal_1858, n2378}), .b ({new_AGEMA_signal_1405, n2377}), .clk ( clk ), .r ( Fresh[863] ), .c ({new_AGEMA_signal_1864, n2379}) ) ;

    /* cells in depth 29 */

    /* cells in depth 30 */
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2377 ( .a ({new_AGEMA_signal_1824, n2212}), .b ({new_AGEMA_signal_1863, n2211}), .clk ( clk ), .r ( Fresh[864] ), .c ({new_AGEMA_signal_1865, N379}) ) ;
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2541 ( .a ({new_AGEMA_signal_1786, n2380}), .b ({new_AGEMA_signal_1864, n2379}), .clk ( clk ), .r ( Fresh[865] ), .c ({new_AGEMA_signal_1866, n2381}) ) ;

    /* cells in depth 31 */

    /* cells in depth 32 */
    nor_GHPC #(.low_latency(0), .pipeline(0)) U2542 ( .a ({new_AGEMA_signal_1785, n2382}), .b ({new_AGEMA_signal_1866, n2381}), .clk ( clk ), .r ( Fresh[866] ), .c ({new_AGEMA_signal_1867, n2427}) ) ;

    /* cells in depth 33 */

    /* cells in depth 34 */
    nand_GHPC #(.low_latency(0), .pipeline(0)) U2584 ( .a ({new_AGEMA_signal_1867, n2427}), .b ({new_AGEMA_signal_1813, n2426}), .clk ( clk ), .r ( Fresh[867] ), .c ({new_AGEMA_signal_1868, N563}) ) ;

    /* register cells */
    reg_masked #(.low_latency(0), .pipeline(0)) SO_reg_7_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1861, N169}), .Q ({SO_s1[7], SO_s0[7]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) SO_reg_6_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1862, N277}), .Q ({SO_s1[6], SO_s0[6]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) SO_reg_5_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1865, N379}), .Q ({SO_s1[5], SO_s0[5]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) SO_reg_4_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1857, N470}), .Q ({SO_s1[4], SO_s0[4]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) SO_reg_3_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1868, N563}), .Q ({SO_s1[3], SO_s0[3]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) SO_reg_2_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1859, N639}), .Q ({SO_s1[2], SO_s0[2]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) SO_reg_1_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1860, N723}), .Q ({SO_s1[1], SO_s0[1]}) ) ;
    reg_masked #(.low_latency(0), .pipeline(0)) SO_reg_0_ ( .clk ( clk_gated ), .D ({new_AGEMA_signal_1853, N789}), .Q ({SO_s1[0], SO_s0[0]}) ) ;
endmodule
