module Reg1(x, y);
 input [174:0] x;
 output [173:0] y;

  assign y[14] = x[3];
  assign y[15] = x[1];
  assign y[16] = x[2];
  assign y[17] = x[170];
  assign y[18] = x[99];
  assign y[19] = x[168];
  assign y[20] = x[169];
  assign y[21] = x[102];
  assign y[22] = x[103];
  assign y[23] = x[98];
  assign y[24] = x[100];
  assign y[25] = x[101];
  assign y[170] = x[171];
  assign y[171] = x[172];
  assign y[172] = x[173];
  assign y[173] = x[174];
  register_stage #(.WIDTH(158)) inst_0(.clk(x[0]), .D({x[4],x[5],x[6],x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[104],x[105],x[106],x[107],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[18],x[19],x[20],x[21],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[26],y[27],y[28],y[29],y[30],y[31],y[32],y[33],y[34],y[35],y[36],y[37],y[38],y[39],y[40],y[41],y[42],y[43],y[44],y[45],y[46],y[47],y[48],y[49],y[50],y[51],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169]}));
endmodule

module Reg2(x, y);
 input [348:0] x;
 output [347:0] y;

  assign y[28] = x[5];
  assign y[29] = x[6];
  assign y[30] = x[1];
  assign y[31] = x[2];
  assign y[32] = x[3];
  assign y[33] = x[4];
  assign y[34] = x[339];
  assign y[35] = x[340];
  assign y[36] = x[197];
  assign y[37] = x[198];
  assign y[38] = x[335];
  assign y[39] = x[336];
  assign y[40] = x[337];
  assign y[41] = x[338];
  assign y[42] = x[203];
  assign y[43] = x[204];
  assign y[44] = x[205];
  assign y[45] = x[206];
  assign y[46] = x[195];
  assign y[47] = x[196];
  assign y[48] = x[199];
  assign y[49] = x[200];
  assign y[50] = x[201];
  assign y[51] = x[202];
  assign y[340] = x[341];
  assign y[341] = x[342];
  assign y[342] = x[343];
  assign y[343] = x[344];
  assign y[344] = x[345];
  assign y[345] = x[346];
  assign y[346] = x[347];
  assign y[347] = x[348];
  register_stage #(.WIDTH(316)) inst_0(.clk(x[0]), .D({x[7],x[8],x[9],x[10],x[11],x[12],x[13],x[14],x[15],x[16],x[17],x[18],x[19],x[20],x[21],x[22],x[23],x[24],x[25],x[26],x[27],x[28],x[29],x[30],x[31],x[32],x[33],x[34],x[207],x[208],x[209],x[210],x[211],x[212],x[213],x[214],x[263],x[264],x[265],x[266],x[267],x[268],x[269],x[270],x[271],x[272],x[273],x[274],x[275],x[276],x[277],x[278],x[279],x[280],x[281],x[282],x[283],x[284],x[285],x[286],x[287],x[288],x[289],x[290],x[291],x[292],x[293],x[294],x[295],x[296],x[297],x[298],x[299],x[300],x[301],x[302],x[303],x[304],x[305],x[306],x[307],x[308],x[309],x[310],x[311],x[312],x[313],x[314],x[315],x[316],x[317],x[318],x[319],x[320],x[321],x[322],x[323],x[324],x[325],x[326],x[327],x[328],x[329],x[330],x[331],x[332],x[333],x[334],x[35],x[36],x[37],x[38],x[39],x[40],x[41],x[42],x[123],x[124],x[125],x[126],x[127],x[128],x[129],x[130],x[131],x[132],x[133],x[134],x[135],x[136],x[137],x[138],x[139],x[140],x[141],x[142],x[143],x[144],x[145],x[146],x[147],x[148],x[149],x[150],x[151],x[152],x[153],x[154],x[155],x[156],x[157],x[158],x[159],x[160],x[161],x[162],x[163],x[164],x[165],x[166],x[167],x[168],x[169],x[170],x[171],x[172],x[173],x[174],x[175],x[176],x[177],x[178],x[179],x[180],x[181],x[182],x[183],x[184],x[185],x[186],x[187],x[188],x[189],x[190],x[191],x[192],x[193],x[194],x[215],x[216],x[217],x[218],x[219],x[220],x[221],x[222],x[223],x[224],x[225],x[226],x[227],x[228],x[229],x[230],x[231],x[232],x[233],x[234],x[235],x[236],x[237],x[238],x[239],x[240],x[241],x[242],x[243],x[244],x[245],x[246],x[247],x[248],x[249],x[250],x[251],x[252],x[253],x[254],x[255],x[256],x[257],x[258],x[259],x[260],x[261],x[262],x[43],x[44],x[45],x[46],x[47],x[48],x[49],x[50],x[51],x[52],x[53],x[54],x[55],x[56],x[57],x[58],x[59],x[60],x[61],x[62],x[63],x[64],x[65],x[66],x[67],x[68],x[69],x[70],x[71],x[72],x[73],x[74],x[75],x[76],x[77],x[78],x[79],x[80],x[81],x[82],x[83],x[84],x[85],x[86],x[87],x[88],x[89],x[90],x[91],x[92],x[93],x[94],x[95],x[96],x[97],x[98],x[99],x[100],x[101],x[102],x[103],x[104],x[105],x[106],x[107],x[108],x[109],x[110],x[111],x[112],x[113],x[114],x[115],x[116],x[117],x[118],x[119],x[120],x[121],x[122]}), .Q({y[0],y[1],y[2],y[3],y[4],y[5],y[6],y[7],y[8],y[9],y[10],y[11],y[12],y[13],y[14],y[15],y[16],y[17],y[18],y[19],y[20],y[21],y[22],y[23],y[24],y[25],y[26],y[27],y[52],y[53],y[54],y[55],y[56],y[57],y[58],y[59],y[60],y[61],y[62],y[63],y[64],y[65],y[66],y[67],y[68],y[69],y[70],y[71],y[72],y[73],y[74],y[75],y[76],y[77],y[78],y[79],y[80],y[81],y[82],y[83],y[84],y[85],y[86],y[87],y[88],y[89],y[90],y[91],y[92],y[93],y[94],y[95],y[96],y[97],y[98],y[99],y[100],y[101],y[102],y[103],y[104],y[105],y[106],y[107],y[108],y[109],y[110],y[111],y[112],y[113],y[114],y[115],y[116],y[117],y[118],y[119],y[120],y[121],y[122],y[123],y[124],y[125],y[126],y[127],y[128],y[129],y[130],y[131],y[132],y[133],y[134],y[135],y[136],y[137],y[138],y[139],y[140],y[141],y[142],y[143],y[144],y[145],y[146],y[147],y[148],y[149],y[150],y[151],y[152],y[153],y[154],y[155],y[156],y[157],y[158],y[159],y[160],y[161],y[162],y[163],y[164],y[165],y[166],y[167],y[168],y[169],y[170],y[171],y[172],y[173],y[174],y[175],y[176],y[177],y[178],y[179],y[180],y[181],y[182],y[183],y[184],y[185],y[186],y[187],y[188],y[189],y[190],y[191],y[192],y[193],y[194],y[195],y[196],y[197],y[198],y[199],y[200],y[201],y[202],y[203],y[204],y[205],y[206],y[207],y[208],y[209],y[210],y[211],y[212],y[213],y[214],y[215],y[216],y[217],y[218],y[219],y[220],y[221],y[222],y[223],y[224],y[225],y[226],y[227],y[228],y[229],y[230],y[231],y[232],y[233],y[234],y[235],y[236],y[237],y[238],y[239],y[240],y[241],y[242],y[243],y[244],y[245],y[246],y[247],y[248],y[249],y[250],y[251],y[252],y[253],y[254],y[255],y[256],y[257],y[258],y[259],y[260],y[261],y[262],y[263],y[264],y[265],y[266],y[267],y[268],y[269],y[270],y[271],y[272],y[273],y[274],y[275],y[276],y[277],y[278],y[279],y[280],y[281],y[282],y[283],y[284],y[285],y[286],y[287],y[288],y[289],y[290],y[291],y[292],y[293],y[294],y[295],y[296],y[297],y[298],y[299],y[300],y[301],y[302],y[303],y[304],y[305],y[306],y[307],y[308],y[309],y[310],y[311],y[312],y[313],y[314],y[315],y[316],y[317],y[318],y[319],y[320],y[321],y[322],y[323],y[324],y[325],y[326],y[327],y[328],y[329],y[330],y[331],y[332],y[333],y[334],y[335],y[336],y[337],y[338],y[339]}));
endmodule

module Fx0(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx1(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx2(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx3(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx4(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx5(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx6(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx7(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx8(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx9(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx10(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx11(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx12(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx13(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx14(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx15(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx16(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx17(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx18(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx19(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx20(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx21(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx22(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx23(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx24(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx25(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx26(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx27(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx28(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx29(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx30(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx31(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx32(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx33(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx34(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx35(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx36(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx37(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx38(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx39(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx40(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx41(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx42(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx43(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx44(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx45(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx46(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx47(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx48(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx49(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx50(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx51(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx52(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx53(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx54(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx55(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx56(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx57(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx58(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx59(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx60(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx61(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx62(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx63(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx64(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx65(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx66(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx67(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx68(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx69(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx70(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx71(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx72(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx73(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx74(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx75(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx76(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx77(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx78(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx79(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx80(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx81(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx82(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx83(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx84(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx85(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx86(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx87(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx88(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx89(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx90(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx91(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx92(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx93(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx94(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx95(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx96(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx97(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx98(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx99(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx100(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx101(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx102(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx103(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx104(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx105(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx106(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx107(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx108(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx109(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx110(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx111(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx112(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx113(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx114(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx115(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx116(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx117(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx118(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx119(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx120(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx121(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx122(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx123(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx124(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx125(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx126(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx127(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx128(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx129(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx130(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx131(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx132(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx133(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx134(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx135(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx136(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx137(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx138(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx139(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx140(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx141(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx142(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx143(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx144(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx145(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx146(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx147(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx148(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx149(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx150(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx151(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx152(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx153(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx154(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx155(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx156(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx157(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx158(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx159(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx160(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx161(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx162(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx163(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx164(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx165(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx166(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx167(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx168(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx169(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx170(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx171(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx172(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx173(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx174(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx175(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx176(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx177(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx178(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx179(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx180(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx181(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx182(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx183(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx184(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx185(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx186(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx187(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx188(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx189(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx190(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx191(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx192(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx193(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx194(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx195(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx196(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx197(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx198(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx199(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx200(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx201(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx202(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx203(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx204(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx205(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx206(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx207(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx208(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx209(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx210(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx211(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx212(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx213(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx214(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx215(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx216(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx217(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx218(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx219(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx220(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx221(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx222(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx223(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx224(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx225(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx226(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx227(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx228(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx229(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx230(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx231(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx232(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx233(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx234(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx235(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx236(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx237(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx238(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx239(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx240(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx241(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx242(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx243(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx244(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx245(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx246(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx247(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx248(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx249(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx250(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx251(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx252(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx253(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx254(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx255(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx256(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx257(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx258(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx259(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx260(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx261(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx262(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx263(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx264(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx265(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx266(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx267(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx268(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx269(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx270(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx271(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx272(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx273(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx274(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx275(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx276(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx277(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx278(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx279(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx280(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx281(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx282(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx283(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx284(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx285(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx286(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx287(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx288(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx289(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx290(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx291(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx292(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx293(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx294(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx295(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx296(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx297(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx298(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx299(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx300(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx301(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx302(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx303(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx304(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx305(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx306(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx307(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx308(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx309(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx310(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx311(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx312(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx313(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx314(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx315(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx316(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx317(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx318(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx319(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx320(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx321(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx322(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx323(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx324(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx325(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx326(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx327(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx328(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx329(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx330(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx331(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx332(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx333(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx334(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx335(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx336(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx337(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx338(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx339(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx340(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx341(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx342(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx343(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx344(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx345(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx346(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module Fx347(x, y);
 input [1:0] x;
 output y;

 wire t;
  assign t = (x[0]);
  assign y = t ^ x[1];
endmodule

module FX(x, y);
 input [521:0] x;
 output [347:0] y;

  Fx0 Fx0_inst(.x({x[1], x[0]}), .y(y[0]));
  Fx1 Fx1_inst(.x({x[2], x[0]}), .y(y[1]));
  Fx2 Fx2_inst(.x({x[4], x[3]}), .y(y[2]));
  Fx3 Fx3_inst(.x({x[5], x[3]}), .y(y[3]));
  Fx4 Fx4_inst(.x({x[7], x[6]}), .y(y[4]));
  Fx5 Fx5_inst(.x({x[8], x[6]}), .y(y[5]));
  Fx6 Fx6_inst(.x({x[10], x[9]}), .y(y[6]));
  Fx7 Fx7_inst(.x({x[11], x[9]}), .y(y[7]));
  Fx8 Fx8_inst(.x({x[13], x[12]}), .y(y[8]));
  Fx9 Fx9_inst(.x({x[14], x[12]}), .y(y[9]));
  Fx10 Fx10_inst(.x({x[16], x[15]}), .y(y[10]));
  Fx11 Fx11_inst(.x({x[17], x[15]}), .y(y[11]));
  Fx12 Fx12_inst(.x({x[19], x[18]}), .y(y[12]));
  Fx13 Fx13_inst(.x({x[20], x[18]}), .y(y[13]));
  Fx14 Fx14_inst(.x({x[22], x[21]}), .y(y[14]));
  Fx15 Fx15_inst(.x({x[23], x[21]}), .y(y[15]));
  Fx16 Fx16_inst(.x({x[25], x[24]}), .y(y[16]));
  Fx17 Fx17_inst(.x({x[26], x[24]}), .y(y[17]));
  Fx18 Fx18_inst(.x({x[28], x[27]}), .y(y[18]));
  Fx19 Fx19_inst(.x({x[29], x[27]}), .y(y[19]));
  Fx20 Fx20_inst(.x({x[31], x[30]}), .y(y[20]));
  Fx21 Fx21_inst(.x({x[32], x[30]}), .y(y[21]));
  Fx22 Fx22_inst(.x({x[34], x[33]}), .y(y[22]));
  Fx23 Fx23_inst(.x({x[35], x[33]}), .y(y[23]));
  Fx24 Fx24_inst(.x({x[37], x[36]}), .y(y[24]));
  Fx25 Fx25_inst(.x({x[38], x[36]}), .y(y[25]));
  Fx26 Fx26_inst(.x({x[40], x[39]}), .y(y[26]));
  Fx27 Fx27_inst(.x({x[41], x[39]}), .y(y[27]));
  Fx28 Fx28_inst(.x({x[43], x[42]}), .y(y[28]));
  Fx29 Fx29_inst(.x({x[44], x[42]}), .y(y[29]));
  Fx30 Fx30_inst(.x({x[46], x[45]}), .y(y[30]));
  Fx31 Fx31_inst(.x({x[47], x[45]}), .y(y[31]));
  Fx32 Fx32_inst(.x({x[49], x[48]}), .y(y[32]));
  Fx33 Fx33_inst(.x({x[50], x[48]}), .y(y[33]));
  Fx34 Fx34_inst(.x({x[52], x[51]}), .y(y[34]));
  Fx35 Fx35_inst(.x({x[53], x[51]}), .y(y[35]));
  Fx36 Fx36_inst(.x({x[55], x[54]}), .y(y[36]));
  Fx37 Fx37_inst(.x({x[56], x[54]}), .y(y[37]));
  Fx38 Fx38_inst(.x({x[58], x[57]}), .y(y[38]));
  Fx39 Fx39_inst(.x({x[59], x[57]}), .y(y[39]));
  Fx40 Fx40_inst(.x({x[61], x[60]}), .y(y[40]));
  Fx41 Fx41_inst(.x({x[62], x[60]}), .y(y[41]));
  Fx42 Fx42_inst(.x({x[64], x[63]}), .y(y[42]));
  Fx43 Fx43_inst(.x({x[65], x[63]}), .y(y[43]));
  Fx44 Fx44_inst(.x({x[67], x[66]}), .y(y[44]));
  Fx45 Fx45_inst(.x({x[68], x[66]}), .y(y[45]));
  Fx46 Fx46_inst(.x({x[70], x[69]}), .y(y[46]));
  Fx47 Fx47_inst(.x({x[71], x[69]}), .y(y[47]));
  Fx48 Fx48_inst(.x({x[73], x[72]}), .y(y[48]));
  Fx49 Fx49_inst(.x({x[74], x[72]}), .y(y[49]));
  Fx50 Fx50_inst(.x({x[76], x[75]}), .y(y[50]));
  Fx51 Fx51_inst(.x({x[77], x[75]}), .y(y[51]));
  Fx52 Fx52_inst(.x({x[79], x[78]}), .y(y[52]));
  Fx53 Fx53_inst(.x({x[80], x[78]}), .y(y[53]));
  Fx54 Fx54_inst(.x({x[82], x[81]}), .y(y[54]));
  Fx55 Fx55_inst(.x({x[83], x[81]}), .y(y[55]));
  Fx56 Fx56_inst(.x({x[85], x[84]}), .y(y[56]));
  Fx57 Fx57_inst(.x({x[86], x[84]}), .y(y[57]));
  Fx58 Fx58_inst(.x({x[88], x[87]}), .y(y[58]));
  Fx59 Fx59_inst(.x({x[89], x[87]}), .y(y[59]));
  Fx60 Fx60_inst(.x({x[91], x[90]}), .y(y[60]));
  Fx61 Fx61_inst(.x({x[92], x[90]}), .y(y[61]));
  Fx62 Fx62_inst(.x({x[94], x[93]}), .y(y[62]));
  Fx63 Fx63_inst(.x({x[95], x[93]}), .y(y[63]));
  Fx64 Fx64_inst(.x({x[97], x[96]}), .y(y[64]));
  Fx65 Fx65_inst(.x({x[98], x[96]}), .y(y[65]));
  Fx66 Fx66_inst(.x({x[100], x[99]}), .y(y[66]));
  Fx67 Fx67_inst(.x({x[101], x[99]}), .y(y[67]));
  Fx68 Fx68_inst(.x({x[103], x[102]}), .y(y[68]));
  Fx69 Fx69_inst(.x({x[104], x[102]}), .y(y[69]));
  Fx70 Fx70_inst(.x({x[106], x[105]}), .y(y[70]));
  Fx71 Fx71_inst(.x({x[107], x[105]}), .y(y[71]));
  Fx72 Fx72_inst(.x({x[109], x[108]}), .y(y[72]));
  Fx73 Fx73_inst(.x({x[110], x[108]}), .y(y[73]));
  Fx74 Fx74_inst(.x({x[112], x[111]}), .y(y[74]));
  Fx75 Fx75_inst(.x({x[113], x[111]}), .y(y[75]));
  Fx76 Fx76_inst(.x({x[115], x[114]}), .y(y[76]));
  Fx77 Fx77_inst(.x({x[116], x[114]}), .y(y[77]));
  Fx78 Fx78_inst(.x({x[118], x[117]}), .y(y[78]));
  Fx79 Fx79_inst(.x({x[119], x[117]}), .y(y[79]));
  Fx80 Fx80_inst(.x({x[121], x[120]}), .y(y[80]));
  Fx81 Fx81_inst(.x({x[122], x[120]}), .y(y[81]));
  Fx82 Fx82_inst(.x({x[124], x[123]}), .y(y[82]));
  Fx83 Fx83_inst(.x({x[125], x[123]}), .y(y[83]));
  Fx84 Fx84_inst(.x({x[127], x[126]}), .y(y[84]));
  Fx85 Fx85_inst(.x({x[128], x[126]}), .y(y[85]));
  Fx86 Fx86_inst(.x({x[130], x[129]}), .y(y[86]));
  Fx87 Fx87_inst(.x({x[131], x[129]}), .y(y[87]));
  Fx88 Fx88_inst(.x({x[133], x[132]}), .y(y[88]));
  Fx89 Fx89_inst(.x({x[134], x[132]}), .y(y[89]));
  Fx90 Fx90_inst(.x({x[136], x[135]}), .y(y[90]));
  Fx91 Fx91_inst(.x({x[137], x[135]}), .y(y[91]));
  Fx92 Fx92_inst(.x({x[139], x[138]}), .y(y[92]));
  Fx93 Fx93_inst(.x({x[140], x[138]}), .y(y[93]));
  Fx94 Fx94_inst(.x({x[142], x[141]}), .y(y[94]));
  Fx95 Fx95_inst(.x({x[143], x[141]}), .y(y[95]));
  Fx96 Fx96_inst(.x({x[145], x[144]}), .y(y[96]));
  Fx97 Fx97_inst(.x({x[146], x[144]}), .y(y[97]));
  Fx98 Fx98_inst(.x({x[148], x[147]}), .y(y[98]));
  Fx99 Fx99_inst(.x({x[149], x[147]}), .y(y[99]));
  Fx100 Fx100_inst(.x({x[151], x[150]}), .y(y[100]));
  Fx101 Fx101_inst(.x({x[152], x[150]}), .y(y[101]));
  Fx102 Fx102_inst(.x({x[154], x[153]}), .y(y[102]));
  Fx103 Fx103_inst(.x({x[155], x[153]}), .y(y[103]));
  Fx104 Fx104_inst(.x({x[157], x[156]}), .y(y[104]));
  Fx105 Fx105_inst(.x({x[158], x[156]}), .y(y[105]));
  Fx106 Fx106_inst(.x({x[160], x[159]}), .y(y[106]));
  Fx107 Fx107_inst(.x({x[161], x[159]}), .y(y[107]));
  Fx108 Fx108_inst(.x({x[163], x[162]}), .y(y[108]));
  Fx109 Fx109_inst(.x({x[164], x[162]}), .y(y[109]));
  Fx110 Fx110_inst(.x({x[166], x[165]}), .y(y[110]));
  Fx111 Fx111_inst(.x({x[167], x[165]}), .y(y[111]));
  Fx112 Fx112_inst(.x({x[169], x[168]}), .y(y[112]));
  Fx113 Fx113_inst(.x({x[170], x[168]}), .y(y[113]));
  Fx114 Fx114_inst(.x({x[172], x[171]}), .y(y[114]));
  Fx115 Fx115_inst(.x({x[173], x[171]}), .y(y[115]));
  Fx116 Fx116_inst(.x({x[175], x[174]}), .y(y[116]));
  Fx117 Fx117_inst(.x({x[176], x[174]}), .y(y[117]));
  Fx118 Fx118_inst(.x({x[178], x[177]}), .y(y[118]));
  Fx119 Fx119_inst(.x({x[179], x[177]}), .y(y[119]));
  Fx120 Fx120_inst(.x({x[181], x[180]}), .y(y[120]));
  Fx121 Fx121_inst(.x({x[182], x[180]}), .y(y[121]));
  Fx122 Fx122_inst(.x({x[184], x[183]}), .y(y[122]));
  Fx123 Fx123_inst(.x({x[185], x[183]}), .y(y[123]));
  Fx124 Fx124_inst(.x({x[187], x[186]}), .y(y[124]));
  Fx125 Fx125_inst(.x({x[188], x[186]}), .y(y[125]));
  Fx126 Fx126_inst(.x({x[190], x[189]}), .y(y[126]));
  Fx127 Fx127_inst(.x({x[191], x[189]}), .y(y[127]));
  Fx128 Fx128_inst(.x({x[193], x[192]}), .y(y[128]));
  Fx129 Fx129_inst(.x({x[194], x[192]}), .y(y[129]));
  Fx130 Fx130_inst(.x({x[196], x[195]}), .y(y[130]));
  Fx131 Fx131_inst(.x({x[197], x[195]}), .y(y[131]));
  Fx132 Fx132_inst(.x({x[199], x[198]}), .y(y[132]));
  Fx133 Fx133_inst(.x({x[200], x[198]}), .y(y[133]));
  Fx134 Fx134_inst(.x({x[202], x[201]}), .y(y[134]));
  Fx135 Fx135_inst(.x({x[203], x[201]}), .y(y[135]));
  Fx136 Fx136_inst(.x({x[205], x[204]}), .y(y[136]));
  Fx137 Fx137_inst(.x({x[206], x[204]}), .y(y[137]));
  Fx138 Fx138_inst(.x({x[208], x[207]}), .y(y[138]));
  Fx139 Fx139_inst(.x({x[209], x[207]}), .y(y[139]));
  Fx140 Fx140_inst(.x({x[211], x[210]}), .y(y[140]));
  Fx141 Fx141_inst(.x({x[212], x[210]}), .y(y[141]));
  Fx142 Fx142_inst(.x({x[214], x[213]}), .y(y[142]));
  Fx143 Fx143_inst(.x({x[215], x[213]}), .y(y[143]));
  Fx144 Fx144_inst(.x({x[217], x[216]}), .y(y[144]));
  Fx145 Fx145_inst(.x({x[218], x[216]}), .y(y[145]));
  Fx146 Fx146_inst(.x({x[220], x[219]}), .y(y[146]));
  Fx147 Fx147_inst(.x({x[221], x[219]}), .y(y[147]));
  Fx148 Fx148_inst(.x({x[223], x[222]}), .y(y[148]));
  Fx149 Fx149_inst(.x({x[224], x[222]}), .y(y[149]));
  Fx150 Fx150_inst(.x({x[226], x[225]}), .y(y[150]));
  Fx151 Fx151_inst(.x({x[227], x[225]}), .y(y[151]));
  Fx152 Fx152_inst(.x({x[229], x[228]}), .y(y[152]));
  Fx153 Fx153_inst(.x({x[230], x[228]}), .y(y[153]));
  Fx154 Fx154_inst(.x({x[232], x[231]}), .y(y[154]));
  Fx155 Fx155_inst(.x({x[233], x[231]}), .y(y[155]));
  Fx156 Fx156_inst(.x({x[235], x[234]}), .y(y[156]));
  Fx157 Fx157_inst(.x({x[236], x[234]}), .y(y[157]));
  Fx158 Fx158_inst(.x({x[238], x[237]}), .y(y[158]));
  Fx159 Fx159_inst(.x({x[239], x[237]}), .y(y[159]));
  Fx160 Fx160_inst(.x({x[241], x[240]}), .y(y[160]));
  Fx161 Fx161_inst(.x({x[242], x[240]}), .y(y[161]));
  Fx162 Fx162_inst(.x({x[244], x[243]}), .y(y[162]));
  Fx163 Fx163_inst(.x({x[245], x[243]}), .y(y[163]));
  Fx164 Fx164_inst(.x({x[247], x[246]}), .y(y[164]));
  Fx165 Fx165_inst(.x({x[248], x[246]}), .y(y[165]));
  Fx166 Fx166_inst(.x({x[250], x[249]}), .y(y[166]));
  Fx167 Fx167_inst(.x({x[251], x[249]}), .y(y[167]));
  Fx168 Fx168_inst(.x({x[253], x[252]}), .y(y[168]));
  Fx169 Fx169_inst(.x({x[254], x[252]}), .y(y[169]));
  Fx170 Fx170_inst(.x({x[256], x[255]}), .y(y[170]));
  Fx171 Fx171_inst(.x({x[257], x[255]}), .y(y[171]));
  Fx172 Fx172_inst(.x({x[259], x[258]}), .y(y[172]));
  Fx173 Fx173_inst(.x({x[260], x[258]}), .y(y[173]));
  Fx174 Fx174_inst(.x({x[262], x[261]}), .y(y[174]));
  Fx175 Fx175_inst(.x({x[263], x[261]}), .y(y[175]));
  Fx176 Fx176_inst(.x({x[265], x[264]}), .y(y[176]));
  Fx177 Fx177_inst(.x({x[266], x[264]}), .y(y[177]));
  Fx178 Fx178_inst(.x({x[268], x[267]}), .y(y[178]));
  Fx179 Fx179_inst(.x({x[269], x[267]}), .y(y[179]));
  Fx180 Fx180_inst(.x({x[271], x[270]}), .y(y[180]));
  Fx181 Fx181_inst(.x({x[272], x[270]}), .y(y[181]));
  Fx182 Fx182_inst(.x({x[274], x[273]}), .y(y[182]));
  Fx183 Fx183_inst(.x({x[275], x[273]}), .y(y[183]));
  Fx184 Fx184_inst(.x({x[277], x[276]}), .y(y[184]));
  Fx185 Fx185_inst(.x({x[278], x[276]}), .y(y[185]));
  Fx186 Fx186_inst(.x({x[280], x[279]}), .y(y[186]));
  Fx187 Fx187_inst(.x({x[281], x[279]}), .y(y[187]));
  Fx188 Fx188_inst(.x({x[283], x[282]}), .y(y[188]));
  Fx189 Fx189_inst(.x({x[284], x[282]}), .y(y[189]));
  Fx190 Fx190_inst(.x({x[286], x[285]}), .y(y[190]));
  Fx191 Fx191_inst(.x({x[287], x[285]}), .y(y[191]));
  Fx192 Fx192_inst(.x({x[289], x[288]}), .y(y[192]));
  Fx193 Fx193_inst(.x({x[290], x[288]}), .y(y[193]));
  Fx194 Fx194_inst(.x({x[292], x[291]}), .y(y[194]));
  Fx195 Fx195_inst(.x({x[293], x[291]}), .y(y[195]));
  Fx196 Fx196_inst(.x({x[295], x[294]}), .y(y[196]));
  Fx197 Fx197_inst(.x({x[296], x[294]}), .y(y[197]));
  Fx198 Fx198_inst(.x({x[298], x[297]}), .y(y[198]));
  Fx199 Fx199_inst(.x({x[299], x[297]}), .y(y[199]));
  Fx200 Fx200_inst(.x({x[301], x[300]}), .y(y[200]));
  Fx201 Fx201_inst(.x({x[302], x[300]}), .y(y[201]));
  Fx202 Fx202_inst(.x({x[304], x[303]}), .y(y[202]));
  Fx203 Fx203_inst(.x({x[305], x[303]}), .y(y[203]));
  Fx204 Fx204_inst(.x({x[307], x[306]}), .y(y[204]));
  Fx205 Fx205_inst(.x({x[308], x[306]}), .y(y[205]));
  Fx206 Fx206_inst(.x({x[310], x[309]}), .y(y[206]));
  Fx207 Fx207_inst(.x({x[311], x[309]}), .y(y[207]));
  Fx208 Fx208_inst(.x({x[313], x[312]}), .y(y[208]));
  Fx209 Fx209_inst(.x({x[314], x[312]}), .y(y[209]));
  Fx210 Fx210_inst(.x({x[316], x[315]}), .y(y[210]));
  Fx211 Fx211_inst(.x({x[317], x[315]}), .y(y[211]));
  Fx212 Fx212_inst(.x({x[319], x[318]}), .y(y[212]));
  Fx213 Fx213_inst(.x({x[320], x[318]}), .y(y[213]));
  Fx214 Fx214_inst(.x({x[322], x[321]}), .y(y[214]));
  Fx215 Fx215_inst(.x({x[323], x[321]}), .y(y[215]));
  Fx216 Fx216_inst(.x({x[325], x[324]}), .y(y[216]));
  Fx217 Fx217_inst(.x({x[326], x[324]}), .y(y[217]));
  Fx218 Fx218_inst(.x({x[328], x[327]}), .y(y[218]));
  Fx219 Fx219_inst(.x({x[329], x[327]}), .y(y[219]));
  Fx220 Fx220_inst(.x({x[331], x[330]}), .y(y[220]));
  Fx221 Fx221_inst(.x({x[332], x[330]}), .y(y[221]));
  Fx222 Fx222_inst(.x({x[334], x[333]}), .y(y[222]));
  Fx223 Fx223_inst(.x({x[335], x[333]}), .y(y[223]));
  Fx224 Fx224_inst(.x({x[337], x[336]}), .y(y[224]));
  Fx225 Fx225_inst(.x({x[338], x[336]}), .y(y[225]));
  Fx226 Fx226_inst(.x({x[340], x[339]}), .y(y[226]));
  Fx227 Fx227_inst(.x({x[341], x[339]}), .y(y[227]));
  Fx228 Fx228_inst(.x({x[343], x[342]}), .y(y[228]));
  Fx229 Fx229_inst(.x({x[344], x[342]}), .y(y[229]));
  Fx230 Fx230_inst(.x({x[346], x[345]}), .y(y[230]));
  Fx231 Fx231_inst(.x({x[347], x[345]}), .y(y[231]));
  Fx232 Fx232_inst(.x({x[349], x[348]}), .y(y[232]));
  Fx233 Fx233_inst(.x({x[350], x[348]}), .y(y[233]));
  Fx234 Fx234_inst(.x({x[352], x[351]}), .y(y[234]));
  Fx235 Fx235_inst(.x({x[353], x[351]}), .y(y[235]));
  Fx236 Fx236_inst(.x({x[355], x[354]}), .y(y[236]));
  Fx237 Fx237_inst(.x({x[356], x[354]}), .y(y[237]));
  Fx238 Fx238_inst(.x({x[358], x[357]}), .y(y[238]));
  Fx239 Fx239_inst(.x({x[359], x[357]}), .y(y[239]));
  Fx240 Fx240_inst(.x({x[361], x[360]}), .y(y[240]));
  Fx241 Fx241_inst(.x({x[362], x[360]}), .y(y[241]));
  Fx242 Fx242_inst(.x({x[364], x[363]}), .y(y[242]));
  Fx243 Fx243_inst(.x({x[365], x[363]}), .y(y[243]));
  Fx244 Fx244_inst(.x({x[367], x[366]}), .y(y[244]));
  Fx245 Fx245_inst(.x({x[368], x[366]}), .y(y[245]));
  Fx246 Fx246_inst(.x({x[370], x[369]}), .y(y[246]));
  Fx247 Fx247_inst(.x({x[371], x[369]}), .y(y[247]));
  Fx248 Fx248_inst(.x({x[373], x[372]}), .y(y[248]));
  Fx249 Fx249_inst(.x({x[374], x[372]}), .y(y[249]));
  Fx250 Fx250_inst(.x({x[376], x[375]}), .y(y[250]));
  Fx251 Fx251_inst(.x({x[377], x[375]}), .y(y[251]));
  Fx252 Fx252_inst(.x({x[379], x[378]}), .y(y[252]));
  Fx253 Fx253_inst(.x({x[380], x[378]}), .y(y[253]));
  Fx254 Fx254_inst(.x({x[382], x[381]}), .y(y[254]));
  Fx255 Fx255_inst(.x({x[383], x[381]}), .y(y[255]));
  Fx256 Fx256_inst(.x({x[385], x[384]}), .y(y[256]));
  Fx257 Fx257_inst(.x({x[386], x[384]}), .y(y[257]));
  Fx258 Fx258_inst(.x({x[388], x[387]}), .y(y[258]));
  Fx259 Fx259_inst(.x({x[389], x[387]}), .y(y[259]));
  Fx260 Fx260_inst(.x({x[391], x[390]}), .y(y[260]));
  Fx261 Fx261_inst(.x({x[392], x[390]}), .y(y[261]));
  Fx262 Fx262_inst(.x({x[394], x[393]}), .y(y[262]));
  Fx263 Fx263_inst(.x({x[395], x[393]}), .y(y[263]));
  Fx264 Fx264_inst(.x({x[397], x[396]}), .y(y[264]));
  Fx265 Fx265_inst(.x({x[398], x[396]}), .y(y[265]));
  Fx266 Fx266_inst(.x({x[400], x[399]}), .y(y[266]));
  Fx267 Fx267_inst(.x({x[401], x[399]}), .y(y[267]));
  Fx268 Fx268_inst(.x({x[403], x[402]}), .y(y[268]));
  Fx269 Fx269_inst(.x({x[404], x[402]}), .y(y[269]));
  Fx270 Fx270_inst(.x({x[406], x[405]}), .y(y[270]));
  Fx271 Fx271_inst(.x({x[407], x[405]}), .y(y[271]));
  Fx272 Fx272_inst(.x({x[409], x[408]}), .y(y[272]));
  Fx273 Fx273_inst(.x({x[410], x[408]}), .y(y[273]));
  Fx274 Fx274_inst(.x({x[412], x[411]}), .y(y[274]));
  Fx275 Fx275_inst(.x({x[413], x[411]}), .y(y[275]));
  Fx276 Fx276_inst(.x({x[415], x[414]}), .y(y[276]));
  Fx277 Fx277_inst(.x({x[416], x[414]}), .y(y[277]));
  Fx278 Fx278_inst(.x({x[418], x[417]}), .y(y[278]));
  Fx279 Fx279_inst(.x({x[419], x[417]}), .y(y[279]));
  Fx280 Fx280_inst(.x({x[421], x[420]}), .y(y[280]));
  Fx281 Fx281_inst(.x({x[422], x[420]}), .y(y[281]));
  Fx282 Fx282_inst(.x({x[424], x[423]}), .y(y[282]));
  Fx283 Fx283_inst(.x({x[425], x[423]}), .y(y[283]));
  Fx284 Fx284_inst(.x({x[427], x[426]}), .y(y[284]));
  Fx285 Fx285_inst(.x({x[428], x[426]}), .y(y[285]));
  Fx286 Fx286_inst(.x({x[430], x[429]}), .y(y[286]));
  Fx287 Fx287_inst(.x({x[431], x[429]}), .y(y[287]));
  Fx288 Fx288_inst(.x({x[433], x[432]}), .y(y[288]));
  Fx289 Fx289_inst(.x({x[434], x[432]}), .y(y[289]));
  Fx290 Fx290_inst(.x({x[436], x[435]}), .y(y[290]));
  Fx291 Fx291_inst(.x({x[437], x[435]}), .y(y[291]));
  Fx292 Fx292_inst(.x({x[439], x[438]}), .y(y[292]));
  Fx293 Fx293_inst(.x({x[440], x[438]}), .y(y[293]));
  Fx294 Fx294_inst(.x({x[442], x[441]}), .y(y[294]));
  Fx295 Fx295_inst(.x({x[443], x[441]}), .y(y[295]));
  Fx296 Fx296_inst(.x({x[445], x[444]}), .y(y[296]));
  Fx297 Fx297_inst(.x({x[446], x[444]}), .y(y[297]));
  Fx298 Fx298_inst(.x({x[448], x[447]}), .y(y[298]));
  Fx299 Fx299_inst(.x({x[449], x[447]}), .y(y[299]));
  Fx300 Fx300_inst(.x({x[451], x[450]}), .y(y[300]));
  Fx301 Fx301_inst(.x({x[452], x[450]}), .y(y[301]));
  Fx302 Fx302_inst(.x({x[454], x[453]}), .y(y[302]));
  Fx303 Fx303_inst(.x({x[455], x[453]}), .y(y[303]));
  Fx304 Fx304_inst(.x({x[457], x[456]}), .y(y[304]));
  Fx305 Fx305_inst(.x({x[458], x[456]}), .y(y[305]));
  Fx306 Fx306_inst(.x({x[460], x[459]}), .y(y[306]));
  Fx307 Fx307_inst(.x({x[461], x[459]}), .y(y[307]));
  Fx308 Fx308_inst(.x({x[463], x[462]}), .y(y[308]));
  Fx309 Fx309_inst(.x({x[464], x[462]}), .y(y[309]));
  Fx310 Fx310_inst(.x({x[466], x[465]}), .y(y[310]));
  Fx311 Fx311_inst(.x({x[467], x[465]}), .y(y[311]));
  Fx312 Fx312_inst(.x({x[469], x[468]}), .y(y[312]));
  Fx313 Fx313_inst(.x({x[470], x[468]}), .y(y[313]));
  Fx314 Fx314_inst(.x({x[472], x[471]}), .y(y[314]));
  Fx315 Fx315_inst(.x({x[473], x[471]}), .y(y[315]));
  Fx316 Fx316_inst(.x({x[475], x[474]}), .y(y[316]));
  Fx317 Fx317_inst(.x({x[476], x[474]}), .y(y[317]));
  Fx318 Fx318_inst(.x({x[478], x[477]}), .y(y[318]));
  Fx319 Fx319_inst(.x({x[479], x[477]}), .y(y[319]));
  Fx320 Fx320_inst(.x({x[481], x[480]}), .y(y[320]));
  Fx321 Fx321_inst(.x({x[482], x[480]}), .y(y[321]));
  Fx322 Fx322_inst(.x({x[484], x[483]}), .y(y[322]));
  Fx323 Fx323_inst(.x({x[485], x[483]}), .y(y[323]));
  Fx324 Fx324_inst(.x({x[487], x[486]}), .y(y[324]));
  Fx325 Fx325_inst(.x({x[488], x[486]}), .y(y[325]));
  Fx326 Fx326_inst(.x({x[490], x[489]}), .y(y[326]));
  Fx327 Fx327_inst(.x({x[491], x[489]}), .y(y[327]));
  Fx328 Fx328_inst(.x({x[493], x[492]}), .y(y[328]));
  Fx329 Fx329_inst(.x({x[494], x[492]}), .y(y[329]));
  Fx330 Fx330_inst(.x({x[496], x[495]}), .y(y[330]));
  Fx331 Fx331_inst(.x({x[497], x[495]}), .y(y[331]));
  Fx332 Fx332_inst(.x({x[499], x[498]}), .y(y[332]));
  Fx333 Fx333_inst(.x({x[500], x[498]}), .y(y[333]));
  Fx334 Fx334_inst(.x({x[502], x[501]}), .y(y[334]));
  Fx335 Fx335_inst(.x({x[503], x[501]}), .y(y[335]));
  Fx336 Fx336_inst(.x({x[505], x[504]}), .y(y[336]));
  Fx337 Fx337_inst(.x({x[506], x[504]}), .y(y[337]));
  Fx338 Fx338_inst(.x({x[508], x[507]}), .y(y[338]));
  Fx339 Fx339_inst(.x({x[509], x[507]}), .y(y[339]));
  Fx340 Fx340_inst(.x({x[511], x[510]}), .y(y[340]));
  Fx341 Fx341_inst(.x({x[512], x[510]}), .y(y[341]));
  Fx342 Fx342_inst(.x({x[514], x[513]}), .y(y[342]));
  Fx343 Fx343_inst(.x({x[515], x[513]}), .y(y[343]));
  Fx344 Fx344_inst(.x({x[517], x[516]}), .y(y[344]));
  Fx345 Fx345_inst(.x({x[518], x[516]}), .y(y[345]));
  Fx346 Fx346_inst(.x({x[520], x[519]}), .y(y[346]));
  Fx347 Fx347_inst(.x({x[521], x[519]}), .y(y[347]));
endmodule

module R1ind0(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind1(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind2(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind3(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind4(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind5(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind6(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind7(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind8(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind9(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind10(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind11(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind12(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind13(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind14(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind15(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind16(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind17(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind18(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind19(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind20(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind21(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind22(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind23(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind24(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind25(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind26(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind27(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind28(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind29(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind30(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind31(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind32(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind33(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind34(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind35(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind36(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind37(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind38(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind39(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind40(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind41(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind42(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind43(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind44(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind45(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind46(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind47(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind48(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind49(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind50(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind51(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind52(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind53(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind54(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind55(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind56(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind57(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind58(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind59(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind60(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind61(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind62(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind63(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind64(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = t[0];
endmodule

module R1ind65(x, y);
 input [26:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = t[19] ^ x[8];
  assign t[11] = t[20] ^ x[11];
  assign t[12] = t[21] ^ x[14];
  assign t[13] = t[22] ^ x[17];
  assign t[14] = t[23] ^ x[20];
  assign t[15] = t[24] ^ x[23];
  assign t[16] = t[25] ^ x[26];
  assign t[17] = (x[0] & x[1]);
  assign t[18] = (x[3] & x[4]);
  assign t[19] = (x[6] & x[7]);
  assign t[1] = ~(t[8] & t[4]);
  assign t[20] = (x[9] & x[10]);
  assign t[21] = (x[12] & x[13]);
  assign t[22] = (x[15] & x[16]);
  assign t[23] = (x[18] & x[19]);
  assign t[24] = (x[21] & x[22]);
  assign t[25] = (x[24] & x[25]);
  assign t[2] = ~(t[9] | t[10]);
  assign t[3] = ~(t[5] | t[11]);
  assign t[4] = ~(t[6] | t[7]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13] & t[14]);
  assign t[7] = ~(t[15] & t[16]);
  assign t[8] = t[17] ^ x[2];
  assign t[9] = t[18] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind66(x, y);
 input [25:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[17] ^ t[18]);
  assign t[11] = ~(t[19]);
  assign t[12] = t[20] ^ x[2];
  assign t[13] = t[21] ^ x[5];
  assign t[14] = t[22] ^ x[8];
  assign t[15] = t[23] ^ x[11];
  assign t[16] = t[24] ^ x[16];
  assign t[17] = t[25] ^ x[19];
  assign t[18] = t[26] ^ x[22];
  assign t[19] = t[27] ^ x[25];
  assign t[1] = ~(t[5] & t[12]);
  assign t[20] = (x[0] & x[1]);
  assign t[21] = (x[3] & x[4]);
  assign t[22] = (x[6] & x[7]);
  assign t[23] = (x[9] & x[10]);
  assign t[24] = (x[14] & x[15]);
  assign t[25] = (x[17] & x[18]);
  assign t[26] = (x[20] & x[21]);
  assign t[27] = (x[23] & x[24]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[13]);
  assign t[4] = ~(t[14] & t[7]);
  assign t[5] = ~(t[14] | t[6]);
  assign t[6] = ~(t[15]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = ~(t[9] ^ t[10]);
  assign t[9] = ~(t[11] | t[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind67(x, y);
 input [25:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13] | t[14]);
  assign t[11] = ~(t[15] | t[13]);
  assign t[12] = t[23] ? t[16] : t[24];
  assign t[13] = ~(t[25]);
  assign t[14] = ~(t[23] ^ t[26]);
  assign t[15] = ~(t[23] | t[26]);
  assign t[16] = ~(t[24] & t[17]);
  assign t[17] = ~(t[18] & t[13]);
  assign t[18] = ~(t[26]);
  assign t[19] = t[27] ^ x[2];
  assign t[1] = ~(t[5] & t[19]);
  assign t[20] = t[28] ^ x[5];
  assign t[21] = t[29] ^ x[8];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = t[31] ^ x[16];
  assign t[24] = t[32] ^ x[19];
  assign t[25] = t[33] ^ x[22];
  assign t[26] = t[34] ^ x[25];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[3] & x[4]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[14] & x[15]);
  assign t[32] = (x[17] & x[18]);
  assign t[33] = (x[20] & x[21]);
  assign t[34] = (x[23] & x[24]);
  assign t[3] = ~(t[20]);
  assign t[4] = ~(t[21] & t[7]);
  assign t[5] = ~(t[21] | t[6]);
  assign t[6] = ~(t[22]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = ~(t[9] | t[10]);
  assign t[9] = ~(t[11] | t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind68(x, y);
 input [25:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[27] | t[15]);
  assign t[12] = ~(t[28] & t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = t[29] ? t[12] : t[28];
  assign t[15] = ~(t[19] | t[20]);
  assign t[16] = ~(t[21] & t[18]);
  assign t[17] = ~(t[29] | t[30]);
  assign t[18] = ~(t[27]);
  assign t[19] = ~(t[29]);
  assign t[1] = ~(t[5] & t[23]);
  assign t[20] = ~(t[21] & t[22]);
  assign t[21] = ~(t[30]);
  assign t[22] = ~(t[28]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[8];
  assign t[26] = t[34] ^ x[11];
  assign t[27] = t[35] ^ x[16];
  assign t[28] = t[36] ^ x[19];
  assign t[29] = t[37] ^ x[22];
  assign t[2] = ~(t[6]);
  assign t[30] = t[38] ^ x[25];
  assign t[31] = (x[0] & x[1]);
  assign t[32] = (x[3] & x[4]);
  assign t[33] = (x[6] & x[7]);
  assign t[34] = (x[9] & x[10]);
  assign t[35] = (x[14] & x[15]);
  assign t[36] = (x[17] & x[18]);
  assign t[37] = (x[20] & x[21]);
  assign t[38] = (x[23] & x[24]);
  assign t[3] = ~(t[24]);
  assign t[4] = ~(t[25] & t[7]);
  assign t[5] = ~(t[25] | t[6]);
  assign t[6] = ~(t[26]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[11] & t[12]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind69(x, y);
 input [25:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = ~(t[13] & t[14]);
  assign t[11] = ~(t[24] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(t[23] | t[25]);
  assign t[14] = ~(t[24]);
  assign t[15] = ~(t[18] & t[16]);
  assign t[16] = ~(t[26]);
  assign t[17] = ~(t[18] & t[14]);
  assign t[18] = ~(t[25]);
  assign t[19] = t[27] ^ x[2];
  assign t[1] = ~(t[5] & t[19]);
  assign t[20] = t[28] ^ x[5];
  assign t[21] = t[29] ^ x[8];
  assign t[22] = t[30] ^ x[11];
  assign t[23] = t[31] ^ x[16];
  assign t[24] = t[32] ^ x[19];
  assign t[25] = t[33] ^ x[22];
  assign t[26] = t[34] ^ x[25];
  assign t[27] = (x[0] & x[1]);
  assign t[28] = (x[3] & x[4]);
  assign t[29] = (x[6] & x[7]);
  assign t[2] = ~(t[6]);
  assign t[30] = (x[9] & x[10]);
  assign t[31] = (x[14] & x[15]);
  assign t[32] = (x[17] & x[18]);
  assign t[33] = (x[20] & x[21]);
  assign t[34] = (x[23] & x[24]);
  assign t[3] = ~(t[20]);
  assign t[4] = ~(t[21] & t[7]);
  assign t[5] = ~(t[21] | t[6]);
  assign t[6] = ~(t[22]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = t[23] ? t[12] : t[11];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind70(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind71(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind72(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind73(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind74(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind75(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind76(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind77(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind78(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind79(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind80(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind81(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind82(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind83(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind84(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind85(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind86(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind87(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind88(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind89(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind90(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind91(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind92(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind93(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind94(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind95(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind96(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind97(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind98(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind99(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind100(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind101(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind102(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind103(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind104(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind105(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind106(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind107(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind108(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind109(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind110(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind111(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind112(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind113(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind114(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind115(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind116(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind117(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind118(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind119(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind120(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind121(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind122(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind123(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind124(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind125(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind126(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind127(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind128(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind129(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind130(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind131(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind132(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind133(x, y);
 input [19:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[16] ^ x[5];
  assign t[11] = t[17] ^ x[8];
  assign t[12] = t[18] ^ x[11];
  assign t[13] = t[19] ^ x[16];
  assign t[14] = t[20] ^ x[19];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[14] & x[15]);
  assign t[1] = ~(t[5] & t[9]);
  assign t[20] = (x[17] & x[18]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[10]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[5] = ~(t[11] | t[6]);
  assign t[6] = ~(t[12]);
  assign t[7] = x[12] ? x[13] : t[8];
  assign t[8] = t[13] ^ t[14];
  assign t[9] = t[15] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind134(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind135(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind136(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind137(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind138(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind139(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind140(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind141(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind142(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind143(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind144(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind145(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind146(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind147(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind148(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind149(x, y);
 input [13:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[12] : t[11];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind150(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind151(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind152(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind153(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind154(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind155(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind156(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind157(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind158(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind159(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind160(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind161(x, y);
 input [16:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[8];
  assign t[11] = t[16] ^ x[11];
  assign t[12] = t[17] ^ x[15];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[13] & x[14]);
  assign t[1] = ~(t[5] & t[8]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[9]);
  assign t[4] = ~(t[10] & t[7]);
  assign t[5] = ~(t[10] | t[6]);
  assign t[6] = ~(t[11]);
  assign t[7] = x[12] ? x[16] : t[12];
  assign t[8] = t[13] ^ x[2];
  assign t[9] = t[14] ^ x[5];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind162(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind163(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind164(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind165(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind166(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind167(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind168(x, y);
 input [13:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[14] ^ x[5];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[11];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[12] : t[11];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[13]);
  assign t[9] = t[13] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind169(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind170(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind171(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind172(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind173(x, y);
 input [16:0] x;
 output y;

 wire [16:0] t;
  assign t[0] = t[7] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[11];
  assign t[11] = t[16] ^ x[15];
  assign t[12] = (x[0] & x[1]);
  assign t[13] = (x[3] & x[4]);
  assign t[14] = (x[6] & x[7]);
  assign t[15] = (x[9] & x[10]);
  assign t[16] = (x[13] & x[14]);
  assign t[1] = ~(t[4] & t[8]);
  assign t[2] = ~(t[9]);
  assign t[3] = ~(t[10] & t[5]);
  assign t[4] = ~(t[10] | t[6]);
  assign t[5] = x[12] ? x[16] : t[11];
  assign t[6] = ~(t[7]);
  assign t[7] = t[12] ^ x[2];
  assign t[8] = t[13] ^ x[5];
  assign t[9] = t[14] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind174(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind175(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind176(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind177(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind178(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind179(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind180(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind181(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind182(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind183(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind184(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind185(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind186(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind187(x, y);
 input [13:0] x;
 output y;

 wire [17:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[14] ^ x[2];
  assign t[11] = t[15] ^ x[5];
  assign t[12] = t[16] ^ x[8];
  assign t[13] = t[17] ^ x[11];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[12] : t[11];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[13]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind188(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind189(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind190(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind191(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind192(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind193(x, y);
 input [16:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = t[9] ? t[3] : t[2];
  assign t[10] = t[15] ^ x[5];
  assign t[11] = t[16] ^ x[8];
  assign t[12] = t[17] ^ x[11];
  assign t[13] = t[18] ^ x[14];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[1] = ~(t[4] & t[10]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12] & t[5]);
  assign t[4] = ~(t[12] | t[6]);
  assign t[5] = t[7] ? x[15] : t[13];
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(x[16]);
  assign t[9] = t[14] ^ x[2];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind194(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind195(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind196(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind197(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind198(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind199(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind200(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind201(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind202(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind203(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind204(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind205(x, y);
 input [16:0] x;
 output y;

 wire [19:0] t;
  assign t[0] = t[2] ? t[4] : t[3];
  assign t[10] = t[15] ^ x[2];
  assign t[11] = t[16] ^ x[5];
  assign t[12] = t[17] ^ x[8];
  assign t[13] = t[18] ^ x[11];
  assign t[14] = t[19] ^ x[14];
  assign t[15] = (x[0] & x[1]);
  assign t[16] = (x[3] & x[4]);
  assign t[17] = (x[6] & x[7]);
  assign t[18] = (x[9] & x[10]);
  assign t[19] = (x[12] & x[13]);
  assign t[1] = ~(t[5] & t[10]);
  assign t[2] = ~(t[6]);
  assign t[3] = ~(t[11]);
  assign t[4] = ~(t[12] & t[7]);
  assign t[5] = ~(t[12] | t[6]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[8] ? x[15] : t[14];
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind206(x, y);
 input [31:0] x;
 output y;

 wire [34:0] t;
  assign t[0] = t[15] ? t[3] : t[2];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[21]);
  assign t[12] = ~(t[22] ^ t[23]);
  assign t[13] = ~(x[28]);
  assign t[14] = ~(t[24]);
  assign t[15] = t[25] ^ x[2];
  assign t[16] = t[26] ^ x[5];
  assign t[17] = t[27] ^ x[8];
  assign t[18] = t[28] ^ x[11];
  assign t[19] = t[29] ^ x[15];
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = t[30] ^ x[18];
  assign t[21] = t[31] ^ x[21];
  assign t[22] = t[32] ^ x[24];
  assign t[23] = t[33] ^ x[27];
  assign t[24] = t[34] ^ x[31];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[6] & x[7]);
  assign t[28] = (x[9] & x[10]);
  assign t[29] = (x[13] & x[14]);
  assign t[2] = ~(t[16]);
  assign t[30] = (x[16] & x[17]);
  assign t[31] = (x[19] & x[20]);
  assign t[32] = (x[22] & x[23]);
  assign t[33] = (x[25] & x[26]);
  assign t[34] = (x[29] & x[30]);
  assign t[3] = ~(t[17] & t[6]);
  assign t[4] = ~(t[17] | t[7]);
  assign t[5] = t[18] ? t[9] : t[8];
  assign t[6] = t[10] ? x[12] : t[16];
  assign t[7] = ~(t[15]);
  assign t[8] = ~(t[11] ^ t[12]);
  assign t[9] = t[19] ^ t[20];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind207(x, y);
 input [34:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[22] ? t[3] : t[2];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[17]);
  assign t[13] = ~(x[22]);
  assign t[14] = ~(t[18] | t[16]);
  assign t[15] = t[29] ? t[19] : t[30];
  assign t[16] = ~(t[31]);
  assign t[17] = ~(t[29] ^ t[32]);
  assign t[18] = ~(t[29] | t[32]);
  assign t[19] = ~(t[30] & t[20]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[21] & t[16]);
  assign t[21] = ~(t[32]);
  assign t[22] = t[33] ^ x[2];
  assign t[23] = t[34] ^ x[5];
  assign t[24] = t[35] ^ x[8];
  assign t[25] = t[36] ^ x[11];
  assign t[26] = t[37] ^ x[14];
  assign t[27] = t[38] ^ x[18];
  assign t[28] = t[39] ^ x[21];
  assign t[29] = t[40] ^ x[25];
  assign t[2] = ~(t[23]);
  assign t[30] = t[41] ^ x[28];
  assign t[31] = t[42] ^ x[31];
  assign t[32] = t[43] ^ x[34];
  assign t[33] = (x[0] & x[1]);
  assign t[34] = (x[3] & x[4]);
  assign t[35] = (x[6] & x[7]);
  assign t[36] = (x[9] & x[10]);
  assign t[37] = (x[12] & x[13]);
  assign t[38] = (x[16] & x[17]);
  assign t[39] = (x[19] & x[20]);
  assign t[3] = ~(t[24] & t[6]);
  assign t[40] = (x[23] & x[24]);
  assign t[41] = (x[26] & x[27]);
  assign t[42] = (x[29] & x[30]);
  assign t[43] = (x[32] & x[33]);
  assign t[4] = ~(t[24] | t[7]);
  assign t[5] = t[25] ? t[9] : t[8];
  assign t[6] = t[10] ? x[15] : t[26];
  assign t[7] = ~(t[22]);
  assign t[8] = ~(t[11] | t[12]);
  assign t[9] = t[27] ^ t[28];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind208(x, y);
 input [34:0] x;
 output y;

 wire [47:0] t;
  assign t[0] = t[26] ? t[3] : t[2];
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(x[22]);
  assign t[14] = ~(t[33] | t[18]);
  assign t[15] = ~(t[34] & t[19]);
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = t[35] ? t[15] : t[34];
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[24] & t[21]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[35] | t[36]);
  assign t[21] = ~(t[33]);
  assign t[22] = ~(t[35]);
  assign t[23] = ~(t[24] & t[25]);
  assign t[24] = ~(t[36]);
  assign t[25] = ~(t[34]);
  assign t[26] = t[37] ^ x[2];
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[8];
  assign t[29] = t[40] ^ x[11];
  assign t[2] = ~(t[27]);
  assign t[30] = t[41] ^ x[14];
  assign t[31] = t[42] ^ x[18];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[25];
  assign t[34] = t[45] ^ x[28];
  assign t[35] = t[46] ^ x[31];
  assign t[36] = t[47] ^ x[34];
  assign t[37] = (x[0] & x[1]);
  assign t[38] = (x[3] & x[4]);
  assign t[39] = (x[6] & x[7]);
  assign t[3] = ~(t[28] & t[6]);
  assign t[40] = (x[9] & x[10]);
  assign t[41] = (x[12] & x[13]);
  assign t[42] = (x[16] & x[17]);
  assign t[43] = (x[19] & x[20]);
  assign t[44] = (x[23] & x[24]);
  assign t[45] = (x[26] & x[27]);
  assign t[46] = (x[29] & x[30]);
  assign t[47] = (x[32] & x[33]);
  assign t[4] = ~(t[28] | t[7]);
  assign t[5] = t[29] ? t[9] : t[8];
  assign t[6] = t[10] ? x[15] : t[30];
  assign t[7] = ~(t[26]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = t[31] ^ t[32];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind209(x, y);
 input [34:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = t[22] ? t[3] : t[2];
  assign t[10] = ~(t[13]);
  assign t[11] = t[29] ? t[15] : t[14];
  assign t[12] = ~(t[16] & t[17]);
  assign t[13] = ~(x[25]);
  assign t[14] = ~(t[30] & t[18]);
  assign t[15] = ~(t[19] & t[20]);
  assign t[16] = ~(t[29] | t[31]);
  assign t[17] = ~(t[30]);
  assign t[18] = ~(t[21] & t[19]);
  assign t[19] = ~(t[32]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[21] & t[17]);
  assign t[21] = ~(t[31]);
  assign t[22] = t[33] ^ x[2];
  assign t[23] = t[34] ^ x[5];
  assign t[24] = t[35] ^ x[8];
  assign t[25] = t[36] ^ x[11];
  assign t[26] = t[37] ^ x[14];
  assign t[27] = t[38] ^ x[18];
  assign t[28] = t[39] ^ x[21];
  assign t[29] = t[40] ^ x[24];
  assign t[2] = ~(t[23]);
  assign t[30] = t[41] ^ x[28];
  assign t[31] = t[42] ^ x[31];
  assign t[32] = t[43] ^ x[34];
  assign t[33] = (x[0] & x[1]);
  assign t[34] = (x[3] & x[4]);
  assign t[35] = (x[6] & x[7]);
  assign t[36] = (x[9] & x[10]);
  assign t[37] = (x[12] & x[13]);
  assign t[38] = (x[16] & x[17]);
  assign t[39] = (x[19] & x[20]);
  assign t[3] = ~(t[24] & t[6]);
  assign t[40] = (x[22] & x[23]);
  assign t[41] = (x[26] & x[27]);
  assign t[42] = (x[29] & x[30]);
  assign t[43] = (x[32] & x[33]);
  assign t[4] = ~(t[24] | t[7]);
  assign t[5] = t[25] ? t[9] : t[8];
  assign t[6] = t[10] ? x[15] : t[26];
  assign t[7] = ~(t[22]);
  assign t[8] = ~(t[11] & t[12]);
  assign t[9] = t[27] ^ t[28];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind210(x, y);
 input [24:0] x;
 output y;

 wire [25:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[18] ^ x[3];
  assign t[11] = t[19] ^ x[6];
  assign t[12] = t[20] ^ x[9];
  assign t[13] = t[21] ^ x[12];
  assign t[14] = t[22] ^ x[15];
  assign t[15] = t[23] ^ x[18];
  assign t[16] = t[24] ^ x[21];
  assign t[17] = t[25] ^ x[24];
  assign t[18] = (x[1] & x[2]);
  assign t[19] = (x[4] & x[5]);
  assign t[1] = ~(x[0]);
  assign t[20] = (x[7] & x[8]);
  assign t[21] = (x[10] & x[11]);
  assign t[22] = (x[13] & x[14]);
  assign t[23] = (x[16] & x[17]);
  assign t[24] = (x[19] & x[20]);
  assign t[25] = (x[22] & x[23]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[6]);
  assign t[4] = ~(t[10]);
  assign t[5] = t[7] & t[11];
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = ~(t[14] & t[15]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = t[0] & t[1];
endmodule

module R1ind211(x, y);
 input [29:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = ~(t[16] ^ t[2]);
  assign t[10] = ~(t[21] | t[11]);
  assign t[11] = ~(t[12]);
  assign t[12] = ~(t[13] & t[14]);
  assign t[13] = ~(t[22]);
  assign t[14] = t[15] & t[23];
  assign t[15] = ~(t[24] | t[25]);
  assign t[16] = t[26] ^ x[2];
  assign t[17] = t[27] ^ x[5];
  assign t[18] = t[28] ^ x[8];
  assign t[19] = t[29] ^ x[11];
  assign t[1] = ~(t[3]);
  assign t[20] = t[30] ^ x[14];
  assign t[21] = t[31] ^ x[17];
  assign t[22] = t[32] ^ x[20];
  assign t[23] = t[33] ^ x[23];
  assign t[24] = t[34] ^ x[26];
  assign t[25] = t[35] ^ x[29];
  assign t[26] = (x[0] & x[1]);
  assign t[27] = (x[3] & x[4]);
  assign t[28] = (x[6] & x[7]);
  assign t[29] = (x[9] & x[10]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[30] = (x[12] & x[13]);
  assign t[31] = (x[15] & x[16]);
  assign t[32] = (x[18] & x[19]);
  assign t[33] = (x[21] & x[22]);
  assign t[34] = (x[24] & x[25]);
  assign t[35] = (x[27] & x[28]);
  assign t[3] = ~(t[17]);
  assign t[4] = ~(t[18]);
  assign t[5] = ~(t[6] & t[19]);
  assign t[6] = ~(t[7] | t[8]);
  assign t[7] = ~(t[20]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[10]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind212(x, y);
 input [26:0] x;
 output y;

 wire [31:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[19]);
  assign t[12] = t[13] & t[20];
  assign t[13] = ~(t[21] | t[22]);
  assign t[14] = t[23] ^ x[2];
  assign t[15] = t[24] ^ x[5];
  assign t[16] = t[25] ^ x[8];
  assign t[17] = t[26] ^ x[11];
  assign t[18] = t[27] ^ x[14];
  assign t[19] = t[28] ^ x[17];
  assign t[1] = t[14] ^ t[3];
  assign t[20] = t[29] ^ x[20];
  assign t[21] = t[30] ^ x[23];
  assign t[22] = t[31] ^ x[26];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[6] & x[7]);
  assign t[26] = (x[9] & x[10]);
  assign t[27] = (x[12] & x[13]);
  assign t[28] = (x[15] & x[16]);
  assign t[29] = (x[18] & x[19]);
  assign t[2] = ~(t[15]);
  assign t[30] = (x[21] & x[22]);
  assign t[31] = (x[24] & x[25]);
  assign t[3] = ~(t[4] & t[16]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[17]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[18] | t[9]);
  assign t[9] = ~(t[10]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind213(x, y);
 input [23:0] x;
 output y;

 wire [28:0] t;
  assign t[0] = ~(t[2] ^ t[13]);
  assign t[10] = ~(t[17]);
  assign t[11] = t[12] & t[18];
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = t[21] ^ x[2];
  assign t[14] = t[22] ^ x[5];
  assign t[15] = t[23] ^ x[8];
  assign t[16] = t[24] ^ x[11];
  assign t[17] = t[25] ^ x[14];
  assign t[18] = t[26] ^ x[17];
  assign t[19] = t[27] ^ x[20];
  assign t[1] = ~(t[3]);
  assign t[20] = t[28] ^ x[23];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[3] & x[4]);
  assign t[23] = (x[6] & x[7]);
  assign t[24] = (x[9] & x[10]);
  assign t[25] = (x[12] & x[13]);
  assign t[26] = (x[15] & x[16]);
  assign t[27] = (x[18] & x[19]);
  assign t[28] = (x[21] & x[22]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(t[14]);
  assign t[4] = ~(t[15]);
  assign t[5] = ~(t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[16] | t[8]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[10] & t[11]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind214(x, y);
 input [20:0] x;
 output y;

 wire [24:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = t[18] ^ x[2];
  assign t[12] = t[19] ^ x[5];
  assign t[13] = t[20] ^ x[8];
  assign t[14] = t[21] ^ x[11];
  assign t[15] = t[22] ^ x[14];
  assign t[16] = t[23] ^ x[17];
  assign t[17] = t[24] ^ x[20];
  assign t[18] = (x[0] & x[1]);
  assign t[19] = (x[3] & x[4]);
  assign t[1] = t[3] ^ t[4];
  assign t[20] = (x[6] & x[7]);
  assign t[21] = (x[9] & x[10]);
  assign t[22] = (x[12] & x[13]);
  assign t[23] = (x[15] & x[16]);
  assign t[24] = (x[18] & x[19]);
  assign t[2] = ~(t[11]);
  assign t[3] = ~(t[12]);
  assign t[4] = ~(t[5]);
  assign t[5] = ~(t[13] | t[6]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[8] & t[9]);
  assign t[8] = ~(t[14]);
  assign t[9] = t[10] & t[15];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind215(x, y);
 input [39:0] x;
 output y;

 wire [46:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = ~(t[11] & t[24]);
  assign t[11] = t[25] & t[12];
  assign t[12] = ~(t[13] | t[14]);
  assign t[13] = ~(t[15] & t[16]);
  assign t[14] = ~(t[17]);
  assign t[15] = ~(t[26]);
  assign t[16] = t[18] & t[27];
  assign t[17] = ~(t[19] | t[20]);
  assign t[18] = ~(t[28] | t[29]);
  assign t[19] = ~(t[30] & t[31]);
  assign t[1] = t[21] ? t[4] : t[3];
  assign t[20] = ~(t[32] & t[33]);
  assign t[21] = t[34] ^ x[2];
  assign t[22] = t[35] ^ x[6];
  assign t[23] = t[36] ^ x[9];
  assign t[24] = t[37] ^ x[12];
  assign t[25] = t[38] ^ x[15];
  assign t[26] = t[39] ^ x[18];
  assign t[27] = t[40] ^ x[21];
  assign t[28] = t[41] ^ x[24];
  assign t[29] = t[42] ^ x[27];
  assign t[2] = ~(x[3]);
  assign t[30] = t[43] ^ x[30];
  assign t[31] = t[44] ^ x[33];
  assign t[32] = t[45] ^ x[36];
  assign t[33] = t[46] ^ x[39];
  assign t[34] = (x[0] & x[1]);
  assign t[35] = (x[4] & x[5]);
  assign t[36] = (x[7] & x[8]);
  assign t[37] = (x[10] & x[11]);
  assign t[38] = (x[13] & x[14]);
  assign t[39] = (x[16] & x[17]);
  assign t[3] = t[5] | t[6];
  assign t[40] = (x[19] & x[20]);
  assign t[41] = (x[22] & x[23]);
  assign t[42] = (x[25] & x[26]);
  assign t[43] = (x[28] & x[29]);
  assign t[44] = (x[31] & x[32]);
  assign t[45] = (x[34] & x[35]);
  assign t[46] = (x[37] & x[38]);
  assign t[4] = ~(t[5] | t[7]);
  assign t[5] = ~(t[22]);
  assign t[6] = ~(t[8] & t[23]);
  assign t[7] = t[9] | t[10];
  assign t[8] = ~(t[10]);
  assign t[9] = ~(t[23]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind216(x, y);
 input [36:0] x;
 output y;

 wire [39:0] t;
  assign t[0] = t[2] ^ t[16];
  assign t[10] = ~(t[20]);
  assign t[11] = t[13] & t[21];
  assign t[12] = ~(t[14] | t[15]);
  assign t[13] = ~(t[22] | t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = ~(t[26] & t[27]);
  assign t[16] = t[28] ^ x[2];
  assign t[17] = t[29] ^ x[6];
  assign t[18] = t[30] ^ x[9];
  assign t[19] = t[31] ^ x[12];
  assign t[1] = ~(t[3]);
  assign t[20] = t[32] ^ x[15];
  assign t[21] = t[33] ^ x[18];
  assign t[22] = t[34] ^ x[21];
  assign t[23] = t[35] ^ x[24];
  assign t[24] = t[36] ^ x[27];
  assign t[25] = t[37] ^ x[30];
  assign t[26] = t[38] ^ x[33];
  assign t[27] = t[39] ^ x[36];
  assign t[28] = (x[0] & x[1]);
  assign t[29] = (x[4] & x[5]);
  assign t[2] = t[4] | t[5];
  assign t[30] = (x[7] & x[8]);
  assign t[31] = (x[10] & x[11]);
  assign t[32] = (x[13] & x[14]);
  assign t[33] = (x[16] & x[17]);
  assign t[34] = (x[19] & x[20]);
  assign t[35] = (x[22] & x[23]);
  assign t[36] = (x[25] & x[26]);
  assign t[37] = (x[28] & x[29]);
  assign t[38] = (x[31] & x[32]);
  assign t[39] = (x[34] & x[35]);
  assign t[3] = ~(x[3]);
  assign t[4] = ~(t[17]);
  assign t[5] = ~(t[6] & t[18]);
  assign t[6] = t[19] & t[7];
  assign t[7] = ~(t[8] | t[9]);
  assign t[8] = ~(t[10] & t[11]);
  assign t[9] = ~(t[12]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind217(x, y);
 input [33:0] x;
 output y;

 wire [35:0] t;
  assign t[0] = t[2] ^ t[14];
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[19] | t[20]);
  assign t[12] = ~(t[21] & t[22]);
  assign t[13] = ~(t[23] & t[24]);
  assign t[14] = t[25] ^ x[2];
  assign t[15] = t[26] ^ x[5];
  assign t[16] = t[27] ^ x[9];
  assign t[17] = t[28] ^ x[12];
  assign t[18] = t[29] ^ x[15];
  assign t[19] = t[30] ^ x[18];
  assign t[1] = ~(t[3]);
  assign t[20] = t[31] ^ x[21];
  assign t[21] = t[32] ^ x[24];
  assign t[22] = t[33] ^ x[27];
  assign t[23] = t[34] ^ x[30];
  assign t[24] = t[35] ^ x[33];
  assign t[25] = (x[0] & x[1]);
  assign t[26] = (x[3] & x[4]);
  assign t[27] = (x[7] & x[8]);
  assign t[28] = (x[10] & x[11]);
  assign t[29] = (x[13] & x[14]);
  assign t[2] = ~(t[4] & t[15]);
  assign t[30] = (x[16] & x[17]);
  assign t[31] = (x[19] & x[20]);
  assign t[32] = (x[22] & x[23]);
  assign t[33] = (x[25] & x[26]);
  assign t[34] = (x[28] & x[29]);
  assign t[35] = (x[31] & x[32]);
  assign t[3] = ~(x[6]);
  assign t[4] = t[16] & t[5];
  assign t[5] = ~(t[6] | t[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[17]);
  assign t[9] = t[11] & t[18];
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind218(x, y);
 input [30:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[2] ^ t[13]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[11] = ~(t[19] & t[20]);
  assign t[12] = ~(t[21] & t[22]);
  assign t[13] = t[23] ^ x[2];
  assign t[14] = t[24] ^ x[5];
  assign t[15] = t[25] ^ x[9];
  assign t[16] = t[26] ^ x[12];
  assign t[17] = t[27] ^ x[15];
  assign t[18] = t[28] ^ x[18];
  assign t[19] = t[29] ^ x[21];
  assign t[1] = ~(t[3]);
  assign t[20] = t[30] ^ x[24];
  assign t[21] = t[31] ^ x[27];
  assign t[22] = t[32] ^ x[30];
  assign t[23] = (x[0] & x[1]);
  assign t[24] = (x[3] & x[4]);
  assign t[25] = (x[7] & x[8]);
  assign t[26] = (x[10] & x[11]);
  assign t[27] = (x[13] & x[14]);
  assign t[28] = (x[16] & x[17]);
  assign t[29] = (x[19] & x[20]);
  assign t[2] = t[14] & t[4];
  assign t[30] = (x[22] & x[23]);
  assign t[31] = (x[25] & x[26]);
  assign t[32] = (x[28] & x[29]);
  assign t[3] = ~(x[6]);
  assign t[4] = ~(t[5] | t[6]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[6] = ~(t[9]);
  assign t[7] = ~(t[15]);
  assign t[8] = t[10] & t[16];
  assign t[9] = ~(t[11] | t[12]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind219(x, y);
 input [27:0] x;
 output y;

 wire [29:0] t;
  assign t[0] = ~(t[12] ^ t[2]);
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = ~(t[19] & t[20]);
  assign t[12] = t[21] ^ x[2];
  assign t[13] = t[22] ^ x[6];
  assign t[14] = t[23] ^ x[9];
  assign t[15] = t[24] ^ x[12];
  assign t[16] = t[25] ^ x[15];
  assign t[17] = t[26] ^ x[18];
  assign t[18] = t[27] ^ x[21];
  assign t[19] = t[28] ^ x[24];
  assign t[1] = ~(t[3]);
  assign t[20] = t[29] ^ x[27];
  assign t[21] = (x[0] & x[1]);
  assign t[22] = (x[4] & x[5]);
  assign t[23] = (x[7] & x[8]);
  assign t[24] = (x[10] & x[11]);
  assign t[25] = (x[13] & x[14]);
  assign t[26] = (x[16] & x[17]);
  assign t[27] = (x[19] & x[20]);
  assign t[28] = (x[22] & x[23]);
  assign t[29] = (x[25] & x[26]);
  assign t[2] = ~(t[4] | t[5]);
  assign t[3] = ~(x[3]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[8]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[9] & t[14];
  assign t[8] = ~(t[10] | t[11]);
  assign t[9] = ~(t[15] | t[16]);
  assign y = ~(t[0] | t[1]);
endmodule

module R1ind220(x, y);
 input [27:0] x;
 output y;

 wire [27:0] t;
  assign t[0] = ~(x[0]);
  assign t[10] = t[19] ^ x[3];
  assign t[11] = t[20] ^ x[6];
  assign t[12] = t[21] ^ x[9];
  assign t[13] = t[22] ^ x[12];
  assign t[14] = t[23] ^ x[15];
  assign t[15] = t[24] ^ x[18];
  assign t[16] = t[25] ^ x[21];
  assign t[17] = t[26] ^ x[24];
  assign t[18] = t[27] ^ x[27];
  assign t[19] = (x[1] & x[2]);
  assign t[1] = ~(t[2] & t[3]);
  assign t[20] = (x[4] & x[5]);
  assign t[21] = (x[7] & x[8]);
  assign t[22] = (x[10] & x[11]);
  assign t[23] = (x[13] & x[14]);
  assign t[24] = (x[16] & x[17]);
  assign t[25] = (x[19] & x[20]);
  assign t[26] = (x[22] & x[23]);
  assign t[27] = (x[25] & x[26]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11] | t[12]);
  assign t[5] = ~(t[7] | t[13]);
  assign t[6] = ~(t[8] | t[9]);
  assign t[7] = ~(t[14]);
  assign t[8] = ~(t[15] & t[16]);
  assign t[9] = ~(t[17] & t[18]);
  assign y = t[0] & t[1];
endmodule

module R1ind221(x, y);
 input [42:0] x;
 output y;

 wire [54:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = ~(t[32]);
  assign t[11] = ~(t[13] & t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19] & t[10]);
  assign t[16] = ~(t[33] & t[20]);
  assign t[17] = ~(t[34] | t[21]);
  assign t[18] = ~(t[22] | t[23]);
  assign t[19] = ~(t[35]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[24]);
  assign t[22] = ~(t[37] & t[38]);
  assign t[23] = ~(t[39] & t[40]);
  assign t[24] = ~(t[19] & t[25]);
  assign t[25] = t[26] & t[36];
  assign t[26] = ~(t[33] | t[32]);
  assign t[27] = t[41] ^ x[3];
  assign t[28] = t[42] ^ x[6];
  assign t[29] = t[43] ^ x[9];
  assign t[2] = ~(t[6] | t[7]);
  assign t[30] = t[44] ^ x[12];
  assign t[31] = t[45] ^ x[15];
  assign t[32] = t[46] ^ x[18];
  assign t[33] = t[47] ^ x[21];
  assign t[34] = t[48] ^ x[24];
  assign t[35] = t[49] ^ x[27];
  assign t[36] = t[50] ^ x[30];
  assign t[37] = t[51] ^ x[33];
  assign t[38] = t[52] ^ x[36];
  assign t[39] = t[53] ^ x[39];
  assign t[3] = ~(t[8] | t[9]);
  assign t[40] = t[54] ^ x[42];
  assign t[41] = (x[1] & x[2]);
  assign t[42] = (x[4] & x[5]);
  assign t[43] = (x[7] & x[8]);
  assign t[44] = (x[10] & x[11]);
  assign t[45] = (x[13] & x[14]);
  assign t[46] = (x[16] & x[17]);
  assign t[47] = (x[19] & x[20]);
  assign t[48] = (x[22] & x[23]);
  assign t[49] = (x[25] & x[26]);
  assign t[4] = ~(t[10] | t[11]);
  assign t[50] = (x[28] & x[29]);
  assign t[51] = (x[31] & x[32]);
  assign t[52] = (x[34] & x[35]);
  assign t[53] = (x[37] & x[38]);
  assign t[54] = (x[40] & x[41]);
  assign t[5] = ~(x[0]);
  assign t[6] = ~(t[27] & t[28]);
  assign t[7] = ~(t[29] & t[30]);
  assign t[8] = ~(t[12]);
  assign t[9] = ~(t[31] & t[5]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind222(x, y);
 input [42:0] x;
 output y;

 wire [57:0] t;
  assign t[0] = ~(t[2] & t[3]);
  assign t[10] = ~(t[30]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[31] | t[20]);
  assign t[13] = ~(t[21] & t[22]);
  assign t[14] = ~(t[32] & t[33]);
  assign t[15] = ~(t[34] & t[35]);
  assign t[16] = ~(t[23]);
  assign t[17] = ~(t[36] & t[7]);
  assign t[18] = ~(t[37] & t[38]);
  assign t[19] = ~(t[39] & t[40]);
  assign t[1] = ~(t[4] & t[5]);
  assign t[20] = ~(t[24]);
  assign t[21] = ~(t[41] | t[42]);
  assign t[22] = ~(t[25] | t[30]);
  assign t[23] = ~(t[26] | t[27]);
  assign t[24] = ~(t[25] & t[28]);
  assign t[25] = ~(t[43]);
  assign t[26] = ~(t[25] & t[29]);
  assign t[27] = ~(t[41] & t[10]);
  assign t[28] = t[21] & t[30];
  assign t[29] = ~(t[42]);
  assign t[2] = ~(t[6] & t[7]);
  assign t[30] = t[44] ^ x[3];
  assign t[31] = t[45] ^ x[6];
  assign t[32] = t[46] ^ x[9];
  assign t[33] = t[47] ^ x[12];
  assign t[34] = t[48] ^ x[15];
  assign t[35] = t[49] ^ x[18];
  assign t[36] = t[50] ^ x[21];
  assign t[37] = t[51] ^ x[24];
  assign t[38] = t[52] ^ x[27];
  assign t[39] = t[53] ^ x[30];
  assign t[3] = ~(t[8] & t[9]);
  assign t[40] = t[54] ^ x[33];
  assign t[41] = t[55] ^ x[36];
  assign t[42] = t[56] ^ x[39];
  assign t[43] = t[57] ^ x[42];
  assign t[44] = (x[1] & x[2]);
  assign t[45] = (x[4] & x[5]);
  assign t[46] = (x[7] & x[8]);
  assign t[47] = (x[10] & x[11]);
  assign t[48] = (x[13] & x[14]);
  assign t[49] = (x[16] & x[17]);
  assign t[4] = ~(t[10]);
  assign t[50] = (x[19] & x[20]);
  assign t[51] = (x[22] & x[23]);
  assign t[52] = (x[25] & x[26]);
  assign t[53] = (x[28] & x[29]);
  assign t[54] = (x[31] & x[32]);
  assign t[55] = (x[34] & x[35]);
  assign t[56] = (x[37] & x[38]);
  assign t[57] = (x[40] & x[41]);
  assign t[5] = ~(t[11]);
  assign t[6] = ~(t[12] & t[13]);
  assign t[7] = ~(x[0]);
  assign t[8] = ~(t[14] | t[15]);
  assign t[9] = ~(t[16] | t[17]);
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind223(x, y);
 input [11:0] x;
 output y;

 wire [11:0] t;
  assign t[0] = ~(t[5] & t[1]);
  assign t[10] = (x[6] & x[7]);
  assign t[11] = (x[9] & x[10]);
  assign t[1] = ~(t[6] | t[2]);
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[7]);
  assign t[4] = t[8] ^ x[2];
  assign t[5] = t[9] ^ x[5];
  assign t[6] = t[10] ^ x[8];
  assign t[7] = t[11] ^ x[11];
  assign t[8] = (x[0] & x[1]);
  assign t[9] = (x[3] & x[4]);
  assign y = ~(t[4] | t[0]);
endmodule

module R1ind224(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind225(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind226(x, y);
 input [20:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[17] ^ x[11];
  assign t[11] = t[18] ^ x[14];
  assign t[12] = t[19] ^ x[17];
  assign t[13] = t[20] ^ x[20];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[19] = (x[15] & x[16]);
  assign t[1] = t[8] ^ t[9];
  assign t[20] = (x[18] & x[19]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[5];
  assign t[9] = t[16] ^ x[8];
  assign y = t[0] ? t[7] : t[1];
endmodule

module R1ind227(x, y);
 input [20:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[17] ^ x[11];
  assign t[11] = t[18] ^ x[14];
  assign t[12] = t[19] ^ x[17];
  assign t[13] = t[20] ^ x[20];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[19] = (x[15] & x[16]);
  assign t[1] = t[8] ^ t[9];
  assign t[20] = (x[18] & x[19]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[5];
  assign t[9] = t[16] ^ x[8];
  assign y = t[0] ? t[7] : t[1];
endmodule

module R1ind228(x, y);
 input [20:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[17] ^ x[11];
  assign t[11] = t[18] ^ x[14];
  assign t[12] = t[19] ^ x[17];
  assign t[13] = t[20] ^ x[20];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[19] = (x[15] & x[16]);
  assign t[1] = t[8] ^ t[9];
  assign t[20] = (x[18] & x[19]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[5];
  assign t[9] = t[16] ^ x[8];
  assign y = t[0] ? t[7] : t[1];
endmodule

module R1ind229(x, y);
 input [20:0] x;
 output y;

 wire [20:0] t;
  assign t[0] = ~(t[2] | t[3]);
  assign t[10] = t[17] ^ x[11];
  assign t[11] = t[18] ^ x[14];
  assign t[12] = t[19] ^ x[17];
  assign t[13] = t[20] ^ x[20];
  assign t[14] = (x[0] & x[1]);
  assign t[15] = (x[3] & x[4]);
  assign t[16] = (x[6] & x[7]);
  assign t[17] = (x[9] & x[10]);
  assign t[18] = (x[12] & x[13]);
  assign t[19] = (x[15] & x[16]);
  assign t[1] = t[8] ^ t[9];
  assign t[20] = (x[18] & x[19]);
  assign t[2] = ~(t[4] & t[5]);
  assign t[3] = ~(t[10] & t[6]);
  assign t[4] = ~(t[11]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = t[14] ^ x[2];
  assign t[8] = t[15] ^ x[5];
  assign t[9] = t[16] ^ x[8];
  assign y = t[0] ? t[7] : t[1];
endmodule

module R1ind230(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind231(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind232(x, y);
 input [12:0] x;
 output y;

 wire [15:0] t;
  assign t[0] = ~(t[2]);
  assign t[10] = t[14] ^ x[9];
  assign t[11] = t[15] ^ x[12];
  assign t[12] = (x[1] & x[2]);
  assign t[13] = (x[4] & x[5]);
  assign t[14] = (x[7] & x[8]);
  assign t[15] = (x[10] & x[11]);
  assign t[1] = ~(x[0]);
  assign t[2] = ~(t[3] | t[4]);
  assign t[3] = ~(t[5] & t[6]);
  assign t[4] = ~(t[8] & t[7]);
  assign t[5] = ~(t[9]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = t[12] ^ x[3];
  assign t[9] = t[13] ^ x[6];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind233(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind234(x, y);
 input [17:0] x;
 output y;

 wire [18:0] t;
  assign t[0] = ~(t[7] | t[2]);
  assign t[10] = t[16] ^ x[11];
  assign t[11] = t[17] ^ x[14];
  assign t[12] = t[18] ^ x[17];
  assign t[13] = (x[0] & x[1]);
  assign t[14] = (x[3] & x[4]);
  assign t[15] = (x[6] & x[7]);
  assign t[16] = (x[9] & x[10]);
  assign t[17] = (x[12] & x[13]);
  assign t[18] = (x[15] & x[16]);
  assign t[1] = ~(t[8]);
  assign t[2] = ~(t[3]);
  assign t[3] = ~(t[4] & t[5]);
  assign t[4] = ~(t[9]);
  assign t[5] = t[6] & t[10];
  assign t[6] = ~(t[11] | t[12]);
  assign t[7] = t[13] ^ x[2];
  assign t[8] = t[14] ^ x[5];
  assign t[9] = t[15] ^ x[8];
  assign y = ~(t[0] & t[1]);
endmodule

module R1ind235(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind236(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind237(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1ind238(x, y);
 input [2:0] x;
 output y;

 wire [1:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (x[0] & x[1]);
  assign y = ~(t[0]);
endmodule

module R1_ind(x, y);
 input [666:0] x;
 output [238:0] y;

  R1ind0 R1ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R1ind1 R1ind1_inst(.x({x[5], x[4], x[3]}), .y(y[1]));
  R1ind2 R1ind2_inst(.x({x[8], x[7], x[6]}), .y(y[2]));
  R1ind3 R1ind3_inst(.x({x[11], x[10], x[9]}), .y(y[3]));
  R1ind4 R1ind4_inst(.x({x[14], x[13], x[12]}), .y(y[4]));
  R1ind5 R1ind5_inst(.x({x[17], x[16], x[15]}), .y(y[5]));
  R1ind6 R1ind6_inst(.x({x[20], x[19], x[18]}), .y(y[6]));
  R1ind7 R1ind7_inst(.x({x[23], x[22], x[21]}), .y(y[7]));
  R1ind8 R1ind8_inst(.x({x[26], x[25], x[24]}), .y(y[8]));
  R1ind9 R1ind9_inst(.x({x[29], x[28], x[27]}), .y(y[9]));
  R1ind10 R1ind10_inst(.x({x[32], x[31], x[30]}), .y(y[10]));
  R1ind11 R1ind11_inst(.x({x[35], x[34], x[33]}), .y(y[11]));
  R1ind12 R1ind12_inst(.x({x[38], x[37], x[36]}), .y(y[12]));
  R1ind13 R1ind13_inst(.x({x[41], x[40], x[39]}), .y(y[13]));
  R1ind14 R1ind14_inst(.x({x[44], x[43], x[42]}), .y(y[14]));
  R1ind15 R1ind15_inst(.x({x[47], x[46], x[45]}), .y(y[15]));
  R1ind16 R1ind16_inst(.x({x[50], x[49], x[48]}), .y(y[16]));
  R1ind17 R1ind17_inst(.x({x[53], x[52], x[51]}), .y(y[17]));
  R1ind18 R1ind18_inst(.x({x[56], x[55], x[54]}), .y(y[18]));
  R1ind19 R1ind19_inst(.x({x[59], x[58], x[57]}), .y(y[19]));
  R1ind20 R1ind20_inst(.x({x[62], x[61], x[60]}), .y(y[20]));
  R1ind21 R1ind21_inst(.x({x[65], x[64], x[63]}), .y(y[21]));
  R1ind22 R1ind22_inst(.x({x[68], x[67], x[66]}), .y(y[22]));
  R1ind23 R1ind23_inst(.x({x[71], x[70], x[69]}), .y(y[23]));
  R1ind24 R1ind24_inst(.x({x[74], x[73], x[72]}), .y(y[24]));
  R1ind25 R1ind25_inst(.x({x[77], x[76], x[75]}), .y(y[25]));
  R1ind26 R1ind26_inst(.x({x[80], x[79], x[78]}), .y(y[26]));
  R1ind27 R1ind27_inst(.x({x[83], x[82], x[81]}), .y(y[27]));
  R1ind28 R1ind28_inst(.x({x[86], x[85], x[84]}), .y(y[28]));
  R1ind29 R1ind29_inst(.x({x[89], x[88], x[87]}), .y(y[29]));
  R1ind30 R1ind30_inst(.x({x[92], x[91], x[90]}), .y(y[30]));
  R1ind31 R1ind31_inst(.x({x[95], x[94], x[93]}), .y(y[31]));
  R1ind32 R1ind32_inst(.x({x[98], x[97], x[96]}), .y(y[32]));
  R1ind33 R1ind33_inst(.x({x[101], x[100], x[99]}), .y(y[33]));
  R1ind34 R1ind34_inst(.x({x[104], x[103], x[102]}), .y(y[34]));
  R1ind35 R1ind35_inst(.x({x[107], x[106], x[105]}), .y(y[35]));
  R1ind36 R1ind36_inst(.x({x[110], x[109], x[108]}), .y(y[36]));
  R1ind37 R1ind37_inst(.x({x[113], x[112], x[111]}), .y(y[37]));
  R1ind38 R1ind38_inst(.x({x[116], x[115], x[114]}), .y(y[38]));
  R1ind39 R1ind39_inst(.x({x[119], x[118], x[117]}), .y(y[39]));
  R1ind40 R1ind40_inst(.x({x[122], x[121], x[120]}), .y(y[40]));
  R1ind41 R1ind41_inst(.x({x[125], x[124], x[123]}), .y(y[41]));
  R1ind42 R1ind42_inst(.x({x[128], x[127], x[126]}), .y(y[42]));
  R1ind43 R1ind43_inst(.x({x[131], x[130], x[129]}), .y(y[43]));
  R1ind44 R1ind44_inst(.x({x[134], x[133], x[132]}), .y(y[44]));
  R1ind45 R1ind45_inst(.x({x[137], x[136], x[135]}), .y(y[45]));
  R1ind46 R1ind46_inst(.x({x[140], x[139], x[138]}), .y(y[46]));
  R1ind47 R1ind47_inst(.x({x[143], x[142], x[141]}), .y(y[47]));
  R1ind48 R1ind48_inst(.x({x[146], x[145], x[144]}), .y(y[48]));
  R1ind49 R1ind49_inst(.x({x[149], x[148], x[147]}), .y(y[49]));
  R1ind50 R1ind50_inst(.x({x[152], x[151], x[150]}), .y(y[50]));
  R1ind51 R1ind51_inst(.x({x[155], x[154], x[153]}), .y(y[51]));
  R1ind52 R1ind52_inst(.x({x[158], x[157], x[156]}), .y(y[52]));
  R1ind53 R1ind53_inst(.x({x[161], x[160], x[159]}), .y(y[53]));
  R1ind54 R1ind54_inst(.x({x[164], x[163], x[162]}), .y(y[54]));
  R1ind55 R1ind55_inst(.x({x[167], x[166], x[165]}), .y(y[55]));
  R1ind56 R1ind56_inst(.x({x[170], x[169], x[168]}), .y(y[56]));
  R1ind57 R1ind57_inst(.x({x[173], x[172], x[171]}), .y(y[57]));
  R1ind58 R1ind58_inst(.x({x[176], x[175], x[174]}), .y(y[58]));
  R1ind59 R1ind59_inst(.x({x[179], x[178], x[177]}), .y(y[59]));
  R1ind60 R1ind60_inst(.x({x[182], x[181], x[180]}), .y(y[60]));
  R1ind61 R1ind61_inst(.x({x[185], x[184], x[183]}), .y(y[61]));
  R1ind62 R1ind62_inst(.x({x[188], x[187], x[186]}), .y(y[62]));
  R1ind63 R1ind63_inst(.x({x[191], x[190], x[189]}), .y(y[63]));
  R1ind64 R1ind64_inst(.x({x[194], x[193], x[192]}), .y(y[64]));
  R1ind65 R1ind65_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195]}), .y(y[65]));
  R1ind66 R1ind66_inst(.x({x[247], x[246], x[245], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[235], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[227], x[226], x[225], x[224], x[223], x[222]}), .y(y[66]));
  R1ind67 R1ind67_inst(.x({x[244], x[243], x[242], x[247], x[246], x[245], x[238], x[237], x[236], x[241], x[240], x[239], x[254], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[253], x[252], x[251], x[250], x[249], x[248]}), .y(y[67]));
  R1ind68 R1ind68_inst(.x({x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[247], x[246], x[245], x[261], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[260], x[259], x[258], x[257], x[256], x[255]}), .y(y[68]));
  R1ind69 R1ind69_inst(.x({x[247], x[246], x[245], x[244], x[243], x[242], x[238], x[237], x[236], x[241], x[240], x[239], x[268], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[267], x[266], x[265], x[264], x[263], x[262]}), .y(y[69]));
  R1ind70 R1ind70_inst(.x({x[272], x[264], x[263], x[262], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[224], x[223], x[222], x[271], x[270], x[269]}), .y(y[70]));
  R1ind71 R1ind71_inst(.x({x[276], x[227], x[226], x[225], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[250], x[249], x[248], x[275], x[274], x[273]}), .y(y[71]));
  R1ind72 R1ind72_inst(.x({x[280], x[253], x[252], x[251], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[257], x[256], x[255], x[279], x[278], x[277]}), .y(y[72]));
  R1ind73 R1ind73_inst(.x({x[284], x[260], x[259], x[258], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[264], x[263], x[262], x[283], x[282], x[281]}), .y(y[73]));
  R1ind74 R1ind74_inst(.x({x[288], x[283], x[282], x[281], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[271], x[270], x[269], x[287], x[286], x[285]}), .y(y[74]));
  R1ind75 R1ind75_inst(.x({x[292], x[224], x[223], x[222], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[275], x[274], x[273], x[291], x[290], x[289]}), .y(y[75]));
  R1ind76 R1ind76_inst(.x({x[296], x[250], x[249], x[248], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[279], x[278], x[277], x[295], x[294], x[293]}), .y(y[76]));
  R1ind77 R1ind77_inst(.x({x[300], x[257], x[256], x[255], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[283], x[282], x[281], x[299], x[298], x[297]}), .y(y[77]));
  R1ind78 R1ind78_inst(.x({x[304], x[299], x[298], x[297], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[287], x[286], x[285], x[303], x[302], x[301]}), .y(y[78]));
  R1ind79 R1ind79_inst(.x({x[308], x[271], x[270], x[269], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[291], x[290], x[289], x[307], x[306], x[305]}), .y(y[79]));
  R1ind80 R1ind80_inst(.x({x[312], x[275], x[274], x[273], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[295], x[294], x[293], x[311], x[310], x[309]}), .y(y[80]));
  R1ind81 R1ind81_inst(.x({x[316], x[279], x[278], x[277], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[299], x[298], x[297], x[315], x[314], x[313]}), .y(y[81]));
  R1ind82 R1ind82_inst(.x({x[320], x[315], x[314], x[313], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[303], x[302], x[301], x[319], x[318], x[317]}), .y(y[82]));
  R1ind83 R1ind83_inst(.x({x[324], x[287], x[286], x[285], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[307], x[306], x[305], x[323], x[322], x[321]}), .y(y[83]));
  R1ind84 R1ind84_inst(.x({x[328], x[291], x[290], x[289], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[311], x[310], x[309], x[327], x[326], x[325]}), .y(y[84]));
  R1ind85 R1ind85_inst(.x({x[332], x[295], x[294], x[293], x[234], x[233], x[232], x[231], x[230], x[229], x[228], x[315], x[314], x[313], x[331], x[330], x[329]}), .y(y[85]));
  R1ind86 R1ind86_inst(.x({x[336], x[331], x[330], x[329], x[234], x[230], x[229], x[228], x[319], x[318], x[317], x[335], x[334], x[333], x[233], x[232], x[231]}), .y(y[86]));
  R1ind87 R1ind87_inst(.x({x[340], x[303], x[302], x[301], x[234], x[230], x[229], x[228], x[323], x[322], x[321], x[339], x[338], x[337], x[233], x[232], x[231]}), .y(y[87]));
  R1ind88 R1ind88_inst(.x({x[344], x[307], x[306], x[305], x[234], x[230], x[229], x[228], x[327], x[326], x[325], x[343], x[342], x[341], x[233], x[232], x[231]}), .y(y[88]));
  R1ind89 R1ind89_inst(.x({x[348], x[311], x[310], x[309], x[234], x[230], x[229], x[228], x[331], x[330], x[329], x[347], x[346], x[345], x[233], x[232], x[231]}), .y(y[89]));
  R1ind90 R1ind90_inst(.x({x[352], x[347], x[346], x[345], x[234], x[230], x[229], x[228], x[335], x[334], x[333], x[351], x[350], x[349], x[233], x[232], x[231]}), .y(y[90]));
  R1ind91 R1ind91_inst(.x({x[356], x[319], x[318], x[317], x[234], x[230], x[229], x[228], x[339], x[338], x[337], x[355], x[354], x[353], x[233], x[232], x[231]}), .y(y[91]));
  R1ind92 R1ind92_inst(.x({x[360], x[323], x[322], x[321], x[234], x[230], x[229], x[228], x[343], x[342], x[341], x[359], x[358], x[357], x[233], x[232], x[231]}), .y(y[92]));
  R1ind93 R1ind93_inst(.x({x[364], x[327], x[326], x[325], x[234], x[230], x[229], x[228], x[347], x[346], x[345], x[363], x[362], x[361], x[233], x[232], x[231]}), .y(y[93]));
  R1ind94 R1ind94_inst(.x({x[371], x[363], x[362], x[361], x[234], x[370], x[369], x[368], x[351], x[350], x[349], x[367], x[366], x[365], x[233], x[232], x[231]}), .y(y[94]));
  R1ind95 R1ind95_inst(.x({x[375], x[335], x[334], x[333], x[234], x[370], x[369], x[368], x[355], x[354], x[353], x[374], x[373], x[372], x[233], x[232], x[231]}), .y(y[95]));
  R1ind96 R1ind96_inst(.x({x[379], x[339], x[338], x[337], x[234], x[370], x[369], x[368], x[359], x[358], x[357], x[378], x[377], x[376], x[233], x[232], x[231]}), .y(y[96]));
  R1ind97 R1ind97_inst(.x({x[383], x[343], x[342], x[341], x[234], x[370], x[369], x[368], x[363], x[362], x[361], x[382], x[381], x[380], x[233], x[232], x[231]}), .y(y[97]));
  R1ind98 R1ind98_inst(.x({x[390], x[382], x[381], x[380], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[367], x[366], x[365], x[386], x[385], x[384]}), .y(y[98]));
  R1ind99 R1ind99_inst(.x({x[394], x[351], x[350], x[349], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[374], x[373], x[372], x[393], x[392], x[391]}), .y(y[99]));
  R1ind100 R1ind100_inst(.x({x[398], x[355], x[354], x[353], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[378], x[377], x[376], x[397], x[396], x[395]}), .y(y[100]));
  R1ind101 R1ind101_inst(.x({x[402], x[359], x[358], x[357], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[382], x[381], x[380], x[401], x[400], x[399]}), .y(y[101]));
  R1ind102 R1ind102_inst(.x({x[406], x[401], x[400], x[399], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[386], x[385], x[384], x[405], x[404], x[403]}), .y(y[102]));
  R1ind103 R1ind103_inst(.x({x[410], x[367], x[366], x[365], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[393], x[392], x[391], x[409], x[408], x[407]}), .y(y[103]));
  R1ind104 R1ind104_inst(.x({x[414], x[374], x[373], x[372], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[397], x[396], x[395], x[413], x[412], x[411]}), .y(y[104]));
  R1ind105 R1ind105_inst(.x({x[418], x[378], x[377], x[376], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[401], x[400], x[399], x[417], x[416], x[415]}), .y(y[105]));
  R1ind106 R1ind106_inst(.x({x[422], x[417], x[416], x[415], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[405], x[404], x[403], x[421], x[420], x[419]}), .y(y[106]));
  R1ind107 R1ind107_inst(.x({x[426], x[386], x[385], x[384], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[409], x[408], x[407], x[425], x[424], x[423]}), .y(y[107]));
  R1ind108 R1ind108_inst(.x({x[430], x[393], x[392], x[391], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[413], x[412], x[411], x[429], x[428], x[427]}), .y(y[108]));
  R1ind109 R1ind109_inst(.x({x[434], x[397], x[396], x[395], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[417], x[416], x[415], x[433], x[432], x[431]}), .y(y[109]));
  R1ind110 R1ind110_inst(.x({x[438], x[433], x[432], x[431], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[421], x[420], x[419], x[437], x[436], x[435]}), .y(y[110]));
  R1ind111 R1ind111_inst(.x({x[442], x[405], x[404], x[403], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[425], x[424], x[423], x[441], x[440], x[439]}), .y(y[111]));
  R1ind112 R1ind112_inst(.x({x[446], x[409], x[408], x[407], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[429], x[428], x[427], x[445], x[444], x[443]}), .y(y[112]));
  R1ind113 R1ind113_inst(.x({x[450], x[413], x[412], x[411], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[433], x[432], x[431], x[449], x[448], x[447]}), .y(y[113]));
  R1ind114 R1ind114_inst(.x({x[454], x[449], x[448], x[447], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[437], x[436], x[435], x[453], x[452], x[451]}), .y(y[114]));
  R1ind115 R1ind115_inst(.x({x[458], x[421], x[420], x[419], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[441], x[440], x[439], x[457], x[456], x[455]}), .y(y[115]));
  R1ind116 R1ind116_inst(.x({x[462], x[425], x[424], x[423], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[445], x[444], x[443], x[461], x[460], x[459]}), .y(y[116]));
  R1ind117 R1ind117_inst(.x({x[466], x[429], x[428], x[427], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[449], x[448], x[447], x[465], x[464], x[463]}), .y(y[117]));
  R1ind118 R1ind118_inst(.x({x[470], x[465], x[464], x[463], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[453], x[452], x[451], x[469], x[468], x[467]}), .y(y[118]));
  R1ind119 R1ind119_inst(.x({x[474], x[437], x[436], x[435], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[457], x[456], x[455], x[473], x[472], x[471]}), .y(y[119]));
  R1ind120 R1ind120_inst(.x({x[478], x[441], x[440], x[439], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[461], x[460], x[459], x[477], x[476], x[475]}), .y(y[120]));
  R1ind121 R1ind121_inst(.x({x[482], x[445], x[444], x[443], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[465], x[464], x[463], x[481], x[480], x[479]}), .y(y[121]));
  R1ind122 R1ind122_inst(.x({x[489], x[481], x[480], x[479], x[234], x[389], x[388], x[387], x[488], x[487], x[486], x[469], x[468], x[467], x[485], x[484], x[483]}), .y(y[122]));
  R1ind123 R1ind123_inst(.x({x[493], x[453], x[452], x[451], x[234], x[389], x[388], x[387], x[488], x[487], x[486], x[473], x[472], x[471], x[492], x[491], x[490]}), .y(y[123]));
  R1ind124 R1ind124_inst(.x({x[497], x[457], x[456], x[455], x[234], x[389], x[388], x[387], x[488], x[487], x[486], x[477], x[476], x[475], x[496], x[495], x[494]}), .y(y[124]));
  R1ind125 R1ind125_inst(.x({x[501], x[461], x[460], x[459], x[234], x[389], x[388], x[387], x[488], x[487], x[486], x[481], x[480], x[479], x[500], x[499], x[498]}), .y(y[125]));
  R1ind126 R1ind126_inst(.x({x[500], x[499], x[498], x[508], x[507], x[506], x[505], x[234], x[389], x[388], x[387], x[488], x[487], x[486], x[485], x[484], x[483], x[504], x[503], x[502]}), .y(y[126]));
  R1ind127 R1ind127_inst(.x({x[469], x[468], x[467], x[515], x[514], x[513], x[512], x[234], x[389], x[388], x[387], x[488], x[487], x[486], x[492], x[491], x[490], x[511], x[510], x[509]}), .y(y[127]));
  R1ind128 R1ind128_inst(.x({x[473], x[472], x[471], x[522], x[521], x[520], x[519], x[234], x[389], x[388], x[387], x[488], x[487], x[486], x[496], x[495], x[494], x[518], x[517], x[516]}), .y(y[128]));
  R1ind129 R1ind129_inst(.x({x[477], x[476], x[475], x[529], x[528], x[527], x[526], x[234], x[389], x[388], x[387], x[488], x[487], x[486], x[500], x[499], x[498], x[525], x[524], x[523]}), .y(y[129]));
  R1ind130 R1ind130_inst(.x({x[533], x[525], x[524], x[523], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[504], x[503], x[502], x[532], x[531], x[530]}), .y(y[130]));
  R1ind131 R1ind131_inst(.x({x[537], x[485], x[484], x[483], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[511], x[510], x[509], x[536], x[535], x[534]}), .y(y[131]));
  R1ind132 R1ind132_inst(.x({x[541], x[492], x[491], x[490], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[518], x[517], x[516], x[540], x[539], x[538]}), .y(y[132]));
  R1ind133 R1ind133_inst(.x({x[496], x[495], x[494], x[548], x[547], x[546], x[545], x[234], x[389], x[388], x[387], x[370], x[369], x[368], x[525], x[524], x[523], x[544], x[543], x[542]}), .y(y[133]));
  R1ind134 R1ind134_inst(.x({x[552], x[544], x[543], x[542], x[234], x[389], x[388], x[387], x[230], x[229], x[228], x[532], x[531], x[530], x[551], x[550], x[549]}), .y(y[134]));
  R1ind135 R1ind135_inst(.x({x[556], x[504], x[503], x[502], x[234], x[389], x[388], x[387], x[230], x[229], x[228], x[536], x[535], x[534], x[555], x[554], x[553]}), .y(y[135]));
  R1ind136 R1ind136_inst(.x({x[560], x[511], x[510], x[509], x[234], x[389], x[388], x[387], x[230], x[229], x[228], x[540], x[539], x[538], x[559], x[558], x[557]}), .y(y[136]));
  R1ind137 R1ind137_inst(.x({x[564], x[518], x[517], x[516], x[234], x[389], x[388], x[387], x[230], x[229], x[228], x[544], x[543], x[542], x[563], x[562], x[561]}), .y(y[137]));
  R1ind138 R1ind138_inst(.x({x[568], x[563], x[562], x[561], x[234], x[370], x[369], x[368], x[551], x[550], x[549], x[567], x[566], x[565], x[389], x[388], x[387]}), .y(y[138]));
  R1ind139 R1ind139_inst(.x({x[572], x[532], x[531], x[530], x[234], x[370], x[369], x[368], x[555], x[554], x[553], x[571], x[570], x[569], x[389], x[388], x[387]}), .y(y[139]));
  R1ind140 R1ind140_inst(.x({x[576], x[536], x[535], x[534], x[234], x[370], x[369], x[368], x[559], x[558], x[557], x[575], x[574], x[573], x[389], x[388], x[387]}), .y(y[140]));
  R1ind141 R1ind141_inst(.x({x[580], x[540], x[539], x[538], x[234], x[370], x[369], x[368], x[563], x[562], x[561], x[579], x[578], x[577], x[389], x[388], x[387]}), .y(y[141]));
  R1ind142 R1ind142_inst(.x({x[581], x[579], x[578], x[577], x[234], x[230], x[229], x[228], x[567], x[566], x[565], x[227], x[226], x[225], x[389], x[388], x[387]}), .y(y[142]));
  R1ind143 R1ind143_inst(.x({x[582], x[551], x[550], x[549], x[234], x[230], x[229], x[228], x[571], x[570], x[569], x[253], x[252], x[251], x[389], x[388], x[387]}), .y(y[143]));
  R1ind144 R1ind144_inst(.x({x[583], x[555], x[554], x[553], x[234], x[230], x[229], x[228], x[575], x[574], x[573], x[260], x[259], x[258], x[389], x[388], x[387]}), .y(y[144]));
  R1ind145 R1ind145_inst(.x({x[584], x[559], x[558], x[557], x[234], x[230], x[229], x[228], x[579], x[578], x[577], x[267], x[266], x[265], x[389], x[388], x[387]}), .y(y[145]));
  R1ind146 R1ind146_inst(.x({x[234], x[591], x[149], x[148], x[147], x[590], x[589], x[588], x[587], x[586], x[585], x[194], x[193], x[192], x[182], x[181], x[180]}), .y(y[146]));
  R1ind147 R1ind147_inst(.x({x[234], x[592], x[161], x[160], x[159], x[590], x[589], x[588], x[587], x[586], x[585], x[191], x[190], x[189], x[179], x[178], x[177]}), .y(y[147]));
  R1ind148 R1ind148_inst(.x({x[593], x[173], x[172], x[171], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[188], x[187], x[186], x[176], x[175], x[174]}), .y(y[148]));
  R1ind149 R1ind149_inst(.x({x[234], x[594], x[590], x[589], x[588], x[587], x[586], x[585], x[185], x[184], x[183], x[173], x[172], x[171]}), .y(y[149]));
  R1ind150 R1ind150_inst(.x({x[595], x[101], x[100], x[99], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[182], x[181], x[180], x[170], x[169], x[168]}), .y(y[150]));
  R1ind151 R1ind151_inst(.x({x[596], x[113], x[112], x[111], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[179], x[178], x[177], x[167], x[166], x[165]}), .y(y[151]));
  R1ind152 R1ind152_inst(.x({x[597], x[125], x[124], x[123], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[176], x[175], x[174], x[164], x[163], x[162]}), .y(y[152]));
  R1ind153 R1ind153_inst(.x({x[598], x[137], x[136], x[135], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[173], x[172], x[171], x[161], x[160], x[159]}), .y(y[153]));
  R1ind154 R1ind154_inst(.x({x[599], x[53], x[52], x[51], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[170], x[169], x[168], x[158], x[157], x[156]}), .y(y[154]));
  R1ind155 R1ind155_inst(.x({x[600], x[65], x[64], x[63], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[167], x[166], x[165], x[155], x[154], x[153]}), .y(y[155]));
  R1ind156 R1ind156_inst(.x({x[601], x[77], x[76], x[75], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[164], x[163], x[162], x[152], x[151], x[150]}), .y(y[156]));
  R1ind157 R1ind157_inst(.x({x[602], x[89], x[88], x[87], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[161], x[160], x[159], x[149], x[148], x[147]}), .y(y[157]));
  R1ind158 R1ind158_inst(.x({x[234], x[603], x[14], x[13], x[12], x[590], x[589], x[588], x[587], x[586], x[585], x[158], x[157], x[156], x[146], x[145], x[144]}), .y(y[158]));
  R1ind159 R1ind159_inst(.x({x[234], x[604], x[17], x[16], x[15], x[590], x[589], x[588], x[587], x[586], x[585], x[155], x[154], x[153], x[143], x[142], x[141]}), .y(y[159]));
  R1ind160 R1ind160_inst(.x({x[234], x[605], x[29], x[28], x[27], x[590], x[589], x[588], x[587], x[586], x[585], x[152], x[151], x[150], x[140], x[139], x[138]}), .y(y[160]));
  R1ind161 R1ind161_inst(.x({x[606], x[41], x[40], x[39], x[234], x[590], x[589], x[588], x[587], x[586], x[585], x[149], x[148], x[147], x[137], x[136], x[135]}), .y(y[161]));
  R1ind162 R1ind162_inst(.x({x[607], x[152], x[151], x[150], x[234], x[587], x[586], x[585], x[146], x[145], x[144], x[134], x[133], x[132], x[590], x[589], x[588]}), .y(y[162]));
  R1ind163 R1ind163_inst(.x({x[608], x[164], x[163], x[162], x[234], x[587], x[586], x[585], x[143], x[142], x[141], x[131], x[130], x[129], x[590], x[589], x[588]}), .y(y[163]));
  R1ind164 R1ind164_inst(.x({x[234], x[609], x[176], x[175], x[174], x[587], x[586], x[585], x[140], x[139], x[138], x[128], x[127], x[126], x[590], x[589], x[588]}), .y(y[164]));
  R1ind165 R1ind165_inst(.x({x[234], x[610], x[188], x[187], x[186], x[587], x[586], x[585], x[137], x[136], x[135], x[125], x[124], x[123], x[590], x[589], x[588]}), .y(y[165]));
  R1ind166 R1ind166_inst(.x({x[611], x[104], x[103], x[102], x[234], x[587], x[586], x[585], x[134], x[133], x[132], x[122], x[121], x[120], x[590], x[589], x[588]}), .y(y[166]));
  R1ind167 R1ind167_inst(.x({x[234], x[612], x[116], x[115], x[114], x[587], x[586], x[585], x[131], x[130], x[129], x[119], x[118], x[117], x[590], x[589], x[588]}), .y(y[167]));
  R1ind168 R1ind168_inst(.x({x[234], x[613], x[587], x[586], x[585], x[128], x[127], x[126], x[116], x[115], x[114], x[590], x[589], x[588]}), .y(y[168]));
  R1ind169 R1ind169_inst(.x({x[614], x[140], x[139], x[138], x[234], x[587], x[586], x[585], x[125], x[124], x[123], x[113], x[112], x[111], x[590], x[589], x[588]}), .y(y[169]));
  R1ind170 R1ind170_inst(.x({x[234], x[615], x[56], x[55], x[54], x[587], x[586], x[585], x[122], x[121], x[120], x[110], x[109], x[108], x[590], x[589], x[588]}), .y(y[170]));
  R1ind171 R1ind171_inst(.x({x[234], x[616], x[68], x[67], x[66], x[587], x[586], x[585], x[119], x[118], x[117], x[107], x[106], x[105], x[590], x[589], x[588]}), .y(y[171]));
  R1ind172 R1ind172_inst(.x({x[234], x[617], x[80], x[79], x[78], x[587], x[586], x[585], x[116], x[115], x[114], x[104], x[103], x[102], x[590], x[589], x[588]}), .y(y[172]));
  R1ind173 R1ind173_inst(.x({x[618], x[92], x[91], x[90], x[234], x[587], x[586], x[585], x[113], x[112], x[111], x[101], x[100], x[99], x[590], x[589], x[588]}), .y(y[173]));
  R1ind174 R1ind174_inst(.x({x[234], x[622], x[11], x[10], x[9], x[590], x[589], x[588], x[621], x[620], x[619], x[110], x[109], x[108], x[98], x[97], x[96]}), .y(y[174]));
  R1ind175 R1ind175_inst(.x({x[234], x[623], x[20], x[19], x[18], x[590], x[589], x[588], x[621], x[620], x[619], x[107], x[106], x[105], x[95], x[94], x[93]}), .y(y[175]));
  R1ind176 R1ind176_inst(.x({x[234], x[624], x[32], x[31], x[30], x[590], x[589], x[588], x[621], x[620], x[619], x[104], x[103], x[102], x[92], x[91], x[90]}), .y(y[176]));
  R1ind177 R1ind177_inst(.x({x[234], x[625], x[44], x[43], x[42], x[590], x[589], x[588], x[621], x[620], x[619], x[101], x[100], x[99], x[89], x[88], x[87]}), .y(y[177]));
  R1ind178 R1ind178_inst(.x({x[234], x[626], x[155], x[154], x[153], x[590], x[589], x[588], x[621], x[620], x[619], x[98], x[97], x[96], x[86], x[85], x[84]}), .y(y[178]));
  R1ind179 R1ind179_inst(.x({x[234], x[627], x[167], x[166], x[165], x[590], x[589], x[588], x[621], x[620], x[619], x[95], x[94], x[93], x[83], x[82], x[81]}), .y(y[179]));
  R1ind180 R1ind180_inst(.x({x[234], x[628], x[179], x[178], x[177], x[590], x[589], x[588], x[621], x[620], x[619], x[92], x[91], x[90], x[80], x[79], x[78]}), .y(y[180]));
  R1ind181 R1ind181_inst(.x({x[234], x[629], x[191], x[190], x[189], x[590], x[589], x[588], x[621], x[620], x[619], x[89], x[88], x[87], x[77], x[76], x[75]}), .y(y[181]));
  R1ind182 R1ind182_inst(.x({x[234], x[630], x[107], x[106], x[105], x[590], x[589], x[588], x[621], x[620], x[619], x[86], x[85], x[84], x[74], x[73], x[72]}), .y(y[182]));
  R1ind183 R1ind183_inst(.x({x[234], x[631], x[119], x[118], x[117], x[590], x[589], x[588], x[621], x[620], x[619], x[83], x[82], x[81], x[71], x[70], x[69]}), .y(y[183]));
  R1ind184 R1ind184_inst(.x({x[234], x[632], x[131], x[130], x[129], x[590], x[589], x[588], x[621], x[620], x[619], x[80], x[79], x[78], x[68], x[67], x[66]}), .y(y[184]));
  R1ind185 R1ind185_inst(.x({x[234], x[633], x[143], x[142], x[141], x[590], x[589], x[588], x[621], x[620], x[619], x[77], x[76], x[75], x[65], x[64], x[63]}), .y(y[185]));
  R1ind186 R1ind186_inst(.x({x[234], x[634], x[59], x[58], x[57], x[590], x[589], x[588], x[621], x[620], x[619], x[74], x[73], x[72], x[62], x[61], x[60]}), .y(y[186]));
  R1ind187 R1ind187_inst(.x({x[234], x[635], x[590], x[589], x[588], x[621], x[620], x[619], x[71], x[70], x[69], x[59], x[58], x[57]}), .y(y[187]));
  R1ind188 R1ind188_inst(.x({x[234], x[636], x[83], x[82], x[81], x[590], x[589], x[588], x[621], x[620], x[619], x[68], x[67], x[66], x[56], x[55], x[54]}), .y(y[188]));
  R1ind189 R1ind189_inst(.x({x[234], x[637], x[95], x[94], x[93], x[590], x[589], x[588], x[621], x[620], x[619], x[65], x[64], x[63], x[53], x[52], x[51]}), .y(y[189]));
  R1ind190 R1ind190_inst(.x({x[234], x[638], x[8], x[7], x[6], x[621], x[620], x[619], x[62], x[61], x[60], x[50], x[49], x[48], x[590], x[589], x[588]}), .y(y[190]));
  R1ind191 R1ind191_inst(.x({x[234], x[639], x[23], x[22], x[21], x[621], x[620], x[619], x[59], x[58], x[57], x[47], x[46], x[45], x[590], x[589], x[588]}), .y(y[191]));
  R1ind192 R1ind192_inst(.x({x[234], x[640], x[35], x[34], x[33], x[621], x[620], x[619], x[56], x[55], x[54], x[44], x[43], x[42], x[590], x[589], x[588]}), .y(y[192]));
  R1ind193 R1ind193_inst(.x({x[234], x[641], x[47], x[46], x[45], x[621], x[620], x[619], x[53], x[52], x[51], x[41], x[40], x[39], x[590], x[589], x[588]}), .y(y[193]));
  R1ind194 R1ind194_inst(.x({x[234], x[642], x[158], x[157], x[156], x[590], x[589], x[588], x[621], x[620], x[619], x[50], x[49], x[48], x[38], x[37], x[36]}), .y(y[194]));
  R1ind195 R1ind195_inst(.x({x[234], x[643], x[170], x[169], x[168], x[590], x[589], x[588], x[621], x[620], x[619], x[47], x[46], x[45], x[35], x[34], x[33]}), .y(y[195]));
  R1ind196 R1ind196_inst(.x({x[234], x[644], x[182], x[181], x[180], x[590], x[589], x[588], x[621], x[620], x[619], x[44], x[43], x[42], x[32], x[31], x[30]}), .y(y[196]));
  R1ind197 R1ind197_inst(.x({x[234], x[645], x[194], x[193], x[192], x[590], x[589], x[588], x[621], x[620], x[619], x[41], x[40], x[39], x[29], x[28], x[27]}), .y(y[197]));
  R1ind198 R1ind198_inst(.x({x[234], x[646], x[110], x[109], x[108], x[590], x[589], x[588], x[621], x[620], x[619], x[38], x[37], x[36], x[26], x[25], x[24]}), .y(y[198]));
  R1ind199 R1ind199_inst(.x({x[234], x[647], x[122], x[121], x[120], x[590], x[589], x[588], x[621], x[620], x[619], x[35], x[34], x[33], x[23], x[22], x[21]}), .y(y[199]));
  R1ind200 R1ind200_inst(.x({x[234], x[648], x[134], x[133], x[132], x[590], x[589], x[588], x[621], x[620], x[619], x[32], x[31], x[30], x[20], x[19], x[18]}), .y(y[200]));
  R1ind201 R1ind201_inst(.x({x[234], x[649], x[146], x[145], x[144], x[590], x[589], x[588], x[621], x[620], x[619], x[29], x[28], x[27], x[17], x[16], x[15]}), .y(y[201]));
  R1ind202 R1ind202_inst(.x({x[234], x[650], x[62], x[61], x[60], x[590], x[589], x[588], x[488], x[487], x[486], x[26], x[25], x[24], x[5], x[4], x[3]}), .y(y[202]));
  R1ind203 R1ind203_inst(.x({x[234], x[651], x[74], x[73], x[72], x[590], x[589], x[588], x[488], x[487], x[486], x[23], x[22], x[21], x[8], x[7], x[6]}), .y(y[203]));
  R1ind204 R1ind204_inst(.x({x[234], x[652], x[86], x[85], x[84], x[590], x[589], x[588], x[488], x[487], x[486], x[20], x[19], x[18], x[11], x[10], x[9]}), .y(y[204]));
  R1ind205 R1ind205_inst(.x({x[234], x[653], x[98], x[97], x[96], x[590], x[589], x[588], x[488], x[487], x[486], x[17], x[16], x[15], x[14], x[13], x[12]}), .y(y[205]));
  R1ind206 R1ind206_inst(.x({x[247], x[246], x[245], x[234], x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[194], x[193], x[192], x[227], x[226], x[225], x[654], x[197], x[196], x[195], x[488], x[487], x[486], x[5], x[4], x[3], x[590], x[589], x[588]}), .y(y[206]));
  R1ind207 R1ind207_inst(.x({x[244], x[243], x[242], x[247], x[246], x[245], x[238], x[237], x[236], x[241], x[240], x[239], x[234], x[191], x[190], x[189], x[253], x[252], x[251], x[655], x[26], x[25], x[24], x[197], x[196], x[195], x[488], x[487], x[486], x[8], x[7], x[6], x[590], x[589], x[588]}), .y(y[207]));
  R1ind208 R1ind208_inst(.x({x[244], x[243], x[242], x[241], x[240], x[239], x[238], x[237], x[236], x[247], x[246], x[245], x[234], x[188], x[187], x[186], x[260], x[259], x[258], x[656], x[38], x[37], x[36], x[197], x[196], x[195], x[488], x[487], x[486], x[11], x[10], x[9], x[590], x[589], x[588]}), .y(y[208]));
  R1ind209 R1ind209_inst(.x({x[247], x[246], x[245], x[244], x[243], x[242], x[238], x[237], x[236], x[234], x[241], x[240], x[239], x[185], x[184], x[183], x[267], x[266], x[265], x[657], x[50], x[49], x[48], x[197], x[196], x[195], x[488], x[487], x[486], x[14], x[13], x[12], x[590], x[589], x[588]}), .y(y[209]));
  R1ind210 R1ind210_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[234]}), .y(y[210]));
  R1ind211 R1ind211_inst(.x({x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[197], x[196], x[195], x[218], x[217], x[216], x[221], x[220], x[219], x[212], x[211], x[210], x[488], x[487], x[486], x[215], x[214], x[213]}), .y(y[211]));
  R1ind212 R1ind212_inst(.x({x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[197], x[196], x[195], x[218], x[217], x[216], x[221], x[220], x[219], x[488], x[487], x[486], x[212], x[211], x[210]}), .y(y[212]));
  R1ind213 R1ind213_inst(.x({x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[197], x[196], x[195], x[218], x[217], x[216], x[488], x[487], x[486], x[221], x[220], x[219]}), .y(y[213]));
  R1ind214 R1ind214_inst(.x({x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[197], x[196], x[195], x[218], x[217], x[216], x[488], x[487], x[486]}), .y(y[214]));
  R1ind215 R1ind215_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[548], x[547], x[546], x[508], x[507], x[506], x[515], x[514], x[513], x[522], x[521], x[520], x[234], x[529], x[528], x[527]}), .y(y[215]));
  R1ind216 R1ind216_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[548], x[547], x[546], x[508], x[507], x[506], x[515], x[514], x[513], x[234], x[522], x[521], x[520]}), .y(y[216]));
  R1ind217 R1ind217_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[548], x[547], x[546], x[234], x[508], x[507], x[506], x[515], x[514], x[513]}), .y(y[217]));
  R1ind218 R1ind218_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[234], x[548], x[547], x[546], x[508], x[507], x[506]}), .y(y[218]));
  R1ind219 R1ind219_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[234], x[548], x[547], x[546]}), .y(y[219]));
  R1ind220 R1ind220_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[209], x[208], x[207], x[206], x[205], x[204], x[203], x[202], x[201], x[200], x[199], x[198], x[197], x[196], x[195], x[234]}), .y(y[220]));
  R1ind221 R1ind221_inst(.x({x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[206], x[205], x[204], x[209], x[208], x[207], x[197], x[196], x[195], x[200], x[199], x[198], x[203], x[202], x[201], x[548], x[547], x[546], x[529], x[528], x[527], x[515], x[514], x[513], x[522], x[521], x[520], x[508], x[507], x[506], x[234]}), .y(y[221]));
  R1ind222 R1ind222_inst(.x({x[209], x[208], x[207], x[203], x[202], x[201], x[200], x[199], x[198], x[221], x[220], x[219], x[218], x[217], x[216], x[215], x[214], x[213], x[212], x[211], x[210], x[548], x[547], x[546], x[529], x[528], x[527], x[515], x[514], x[513], x[522], x[521], x[520], x[508], x[507], x[506], x[197], x[196], x[195], x[206], x[205], x[204], x[234]}), .y(y[222]));
  R1ind223 R1ind223_inst(.x({x[206], x[205], x[204], x[209], x[208], x[207], x[203], x[202], x[201], x[200], x[199], x[198]}), .y(y[223]));
  R1ind224 R1ind224_inst(.x({x[660], x[659], x[658]}), .y(y[224]));
  R1ind225 R1ind225_inst(.x({x[663], x[662], x[661]}), .y(y[225]));
  R1ind226 R1ind226_inst(.x({x[206], x[205], x[204], x[203], x[202], x[201], x[209], x[208], x[207], x[200], x[199], x[198], x[191], x[190], x[189], x[253], x[252], x[251], x[567], x[566], x[565]}), .y(y[226]));
  R1ind227 R1ind227_inst(.x({x[206], x[205], x[204], x[203], x[202], x[201], x[209], x[208], x[207], x[200], x[199], x[198], x[185], x[184], x[183], x[267], x[266], x[265], x[575], x[574], x[573]}), .y(y[227]));
  R1ind228 R1ind228_inst(.x({x[206], x[205], x[204], x[203], x[202], x[201], x[209], x[208], x[207], x[200], x[199], x[198], x[194], x[193], x[192], x[227], x[226], x[225], x[267], x[266], x[265]}), .y(y[228]));
  R1ind229 R1ind229_inst(.x({x[206], x[205], x[204], x[203], x[202], x[201], x[209], x[208], x[207], x[200], x[199], x[198], x[188], x[187], x[186], x[260], x[259], x[258], x[571], x[570], x[569]}), .y(y[229]));
  R1ind230 R1ind230_inst(.x({x[660], x[659], x[658]}), .y(y[230]));
  R1ind231 R1ind231_inst(.x({x[663], x[662], x[661]}), .y(y[231]));
  R1ind232 R1ind232_inst(.x({x[206], x[205], x[204], x[203], x[202], x[201], x[209], x[208], x[207], x[200], x[199], x[198], x[234]}), .y(y[232]));
  R1ind233 R1ind233_inst(.x({x[666], x[665], x[664]}), .y(y[233]));
  R1ind234 R1ind234_inst(.x({x[203], x[202], x[201], x[200], x[199], x[198], x[206], x[205], x[204], x[209], x[208], x[207], x[488], x[487], x[486], x[197], x[196], x[195]}), .y(y[234]));
  R1ind235 R1ind235_inst(.x({x[666], x[665], x[664]}), .y(y[235]));
  R1ind236 R1ind236_inst(.x({x[488], x[487], x[486]}), .y(y[236]));
  R1ind237 R1ind237_inst(.x({x[590], x[589], x[588]}), .y(y[237]));
  R1ind238 R1ind238_inst(.x({x[488], x[487], x[486]}), .y(y[238]));
endmodule

module R2ind0(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (t[2] & ~t[3]);
  assign t[2] = t[4] ^ x[2];
  assign t[3] = t[5] ^ x[1];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind1(x, y);
 input [2:0] x;
 output y;

 wire [5:0] t;
  assign t[0] = t[1] ^ x[2];
  assign t[1] = (~t[2] & t[3]);
  assign t[2] = t[4] ^ x[1];
  assign t[3] = t[5] ^ x[2];
  assign t[4] = (x[0]);
  assign t[5] = (x[0]);
  assign y = t[0];
endmodule

module R2ind2(x, y);
 input [26:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[5];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[29] ^ x[8];
  assign t[21] = t[30] ^ x[11];
  assign t[22] = t[31] ^ x[14];
  assign t[23] = t[32] ^ x[17];
  assign t[24] = t[33] ^ x[20];
  assign t[25] = t[34] ^ x[23];
  assign t[26] = t[35] ^ x[26];
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = (t[38] & ~t[39]);
  assign t[29] = (t[40] & ~t[41]);
  assign t[2] = ~(t[9] & t[5]);
  assign t[30] = (t[42] & ~t[43]);
  assign t[31] = (t[44] & ~t[45]);
  assign t[32] = (t[46] & ~t[47]);
  assign t[33] = (t[48] & ~t[49]);
  assign t[34] = (t[50] & ~t[51]);
  assign t[35] = (t[52] & ~t[53]);
  assign t[36] = t[54] ^ x[2];
  assign t[37] = t[55] ^ x[1];
  assign t[38] = t[56] ^ x[5];
  assign t[39] = t[57] ^ x[4];
  assign t[3] = ~(t[10] | t[11]);
  assign t[40] = t[58] ^ x[8];
  assign t[41] = t[59] ^ x[7];
  assign t[42] = t[60] ^ x[11];
  assign t[43] = t[61] ^ x[10];
  assign t[44] = t[62] ^ x[14];
  assign t[45] = t[63] ^ x[13];
  assign t[46] = t[64] ^ x[17];
  assign t[47] = t[65] ^ x[16];
  assign t[48] = t[66] ^ x[20];
  assign t[49] = t[67] ^ x[19];
  assign t[4] = ~(t[6] | t[12]);
  assign t[50] = t[68] ^ x[23];
  assign t[51] = t[69] ^ x[22];
  assign t[52] = t[70] ^ x[26];
  assign t[53] = t[71] ^ x[25];
  assign t[54] = (x[0]);
  assign t[55] = (x[0]);
  assign t[56] = (x[3]);
  assign t[57] = (x[3]);
  assign t[58] = (x[6]);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[9]);
  assign t[61] = (x[9]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[15]);
  assign t[65] = (x[15]);
  assign t[66] = (x[18]);
  assign t[67] = (x[18]);
  assign t[68] = (x[21]);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[13]);
  assign t[70] = (x[24]);
  assign t[71] = (x[24]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[8] = ~(t[16] & t[17]);
  assign t[9] = (t[18]);
  assign y = (t[0]);
endmodule

module R2ind3(x, y);
 input [26:0] x;
 output y;

 wire [71:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = t[27] ^ x[2];
  assign t[19] = t[28] ^ x[5];
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = t[29] ^ x[8];
  assign t[21] = t[30] ^ x[11];
  assign t[22] = t[31] ^ x[14];
  assign t[23] = t[32] ^ x[17];
  assign t[24] = t[33] ^ x[20];
  assign t[25] = t[34] ^ x[23];
  assign t[26] = t[35] ^ x[26];
  assign t[27] = (t[36] & ~t[37]);
  assign t[28] = (t[38] & ~t[39]);
  assign t[29] = (t[40] & ~t[41]);
  assign t[2] = ~(t[9] & t[5]);
  assign t[30] = (t[42] & ~t[43]);
  assign t[31] = (t[44] & ~t[45]);
  assign t[32] = (t[46] & ~t[47]);
  assign t[33] = (t[48] & ~t[49]);
  assign t[34] = (t[50] & ~t[51]);
  assign t[35] = (t[52] & ~t[53]);
  assign t[36] = t[54] ^ x[2];
  assign t[37] = t[55] ^ x[1];
  assign t[38] = t[56] ^ x[5];
  assign t[39] = t[57] ^ x[4];
  assign t[3] = ~(t[10] | t[11]);
  assign t[40] = t[58] ^ x[8];
  assign t[41] = t[59] ^ x[7];
  assign t[42] = t[60] ^ x[11];
  assign t[43] = t[61] ^ x[10];
  assign t[44] = t[62] ^ x[14];
  assign t[45] = t[63] ^ x[13];
  assign t[46] = t[64] ^ x[17];
  assign t[47] = t[65] ^ x[16];
  assign t[48] = t[66] ^ x[20];
  assign t[49] = t[67] ^ x[19];
  assign t[4] = ~(t[6] | t[12]);
  assign t[50] = t[68] ^ x[23];
  assign t[51] = t[69] ^ x[22];
  assign t[52] = t[70] ^ x[26];
  assign t[53] = t[71] ^ x[25];
  assign t[54] = (x[0]);
  assign t[55] = (x[0]);
  assign t[56] = (x[3]);
  assign t[57] = (x[3]);
  assign t[58] = (x[6]);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[7] | t[8]);
  assign t[60] = (x[9]);
  assign t[61] = (x[9]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[15]);
  assign t[65] = (x[15]);
  assign t[66] = (x[18]);
  assign t[67] = (x[18]);
  assign t[68] = (x[21]);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[13]);
  assign t[70] = (x[24]);
  assign t[71] = (x[24]);
  assign t[7] = ~(t[14] & t[15]);
  assign t[8] = ~(t[16] & t[17]);
  assign t[9] = (t[18]);
  assign y = (t[0]);
endmodule

module R2ind4(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = (t[19]);
  assign t[12] = (t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = t[27] ^ x[3];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[28] ^ x[6];
  assign t[21] = t[29] ^ x[9];
  assign t[22] = t[30] ^ x[12];
  assign t[23] = t[31] ^ x[15];
  assign t[24] = t[32] ^ x[18];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = t[34] ^ x[24];
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = (t[39] & ~t[40]);
  assign t[2] = ~(x[0]);
  assign t[30] = (t[41] & ~t[42]);
  assign t[31] = (t[43] & ~t[44]);
  assign t[32] = (t[45] & ~t[46]);
  assign t[33] = (t[47] & ~t[48]);
  assign t[34] = (t[49] & ~t[50]);
  assign t[35] = t[51] ^ x[3];
  assign t[36] = t[52] ^ x[2];
  assign t[37] = t[53] ^ x[6];
  assign t[38] = t[54] ^ x[5];
  assign t[39] = t[55] ^ x[9];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[56] ^ x[8];
  assign t[41] = t[57] ^ x[12];
  assign t[42] = t[58] ^ x[11];
  assign t[43] = t[59] ^ x[15];
  assign t[44] = t[60] ^ x[14];
  assign t[45] = t[61] ^ x[18];
  assign t[46] = t[62] ^ x[17];
  assign t[47] = t[63] ^ x[21];
  assign t[48] = t[64] ^ x[20];
  assign t[49] = t[65] ^ x[24];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[23];
  assign t[51] = (x[1]);
  assign t[52] = (x[1]);
  assign t[53] = (x[4]);
  assign t[54] = (x[4]);
  assign t[55] = (x[7]);
  assign t[56] = (x[7]);
  assign t[57] = (x[10]);
  assign t[58] = (x[10]);
  assign t[59] = (x[13]);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[13]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[19]);
  assign t[64] = (x[19]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[6] = t[8] & t[12];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[13] | t[14]);
  assign t[9] = ~(t[15] & t[16]);
  assign y = (t[0]);
endmodule

module R2ind5(x, y);
 input [24:0] x;
 output y;

 wire [66:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[17] & t[18]);
  assign t[11] = (t[19]);
  assign t[12] = (t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = t[27] ^ x[3];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[28] ^ x[6];
  assign t[21] = t[29] ^ x[9];
  assign t[22] = t[30] ^ x[12];
  assign t[23] = t[31] ^ x[15];
  assign t[24] = t[32] ^ x[18];
  assign t[25] = t[33] ^ x[21];
  assign t[26] = t[34] ^ x[24];
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = (t[39] & ~t[40]);
  assign t[2] = ~(x[0]);
  assign t[30] = (t[41] & ~t[42]);
  assign t[31] = (t[43] & ~t[44]);
  assign t[32] = (t[45] & ~t[46]);
  assign t[33] = (t[47] & ~t[48]);
  assign t[34] = (t[49] & ~t[50]);
  assign t[35] = t[51] ^ x[3];
  assign t[36] = t[52] ^ x[2];
  assign t[37] = t[53] ^ x[6];
  assign t[38] = t[54] ^ x[5];
  assign t[39] = t[55] ^ x[9];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[56] ^ x[8];
  assign t[41] = t[57] ^ x[12];
  assign t[42] = t[58] ^ x[11];
  assign t[43] = t[59] ^ x[15];
  assign t[44] = t[60] ^ x[14];
  assign t[45] = t[61] ^ x[18];
  assign t[46] = t[62] ^ x[17];
  assign t[47] = t[63] ^ x[21];
  assign t[48] = t[64] ^ x[20];
  assign t[49] = t[65] ^ x[24];
  assign t[4] = ~(t[7]);
  assign t[50] = t[66] ^ x[23];
  assign t[51] = (x[1]);
  assign t[52] = (x[1]);
  assign t[53] = (x[4]);
  assign t[54] = (x[4]);
  assign t[55] = (x[7]);
  assign t[56] = (x[7]);
  assign t[57] = (x[10]);
  assign t[58] = (x[10]);
  assign t[59] = (x[13]);
  assign t[5] = ~(t[11]);
  assign t[60] = (x[13]);
  assign t[61] = (x[16]);
  assign t[62] = (x[16]);
  assign t[63] = (x[19]);
  assign t[64] = (x[19]);
  assign t[65] = (x[22]);
  assign t[66] = (x[22]);
  assign t[6] = t[8] & t[12];
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[13] | t[14]);
  assign t[9] = ~(t[15] & t[16]);
  assign y = (t[0]);
endmodule

module R2ind6(x, y);
 input [42:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[4]);
  assign t[101] = (x[4]);
  assign t[102] = (x[7]);
  assign t[103] = (x[7]);
  assign t[104] = (x[10]);
  assign t[105] = (x[10]);
  assign t[106] = (x[13]);
  assign t[107] = (x[13]);
  assign t[108] = (x[16]);
  assign t[109] = (x[16]);
  assign t[10] = ~(t[32] & t[6]);
  assign t[110] = (x[19]);
  assign t[111] = (x[19]);
  assign t[112] = (x[22]);
  assign t[113] = (x[22]);
  assign t[114] = (x[25]);
  assign t[115] = (x[25]);
  assign t[116] = (x[28]);
  assign t[117] = (x[28]);
  assign t[118] = (x[31]);
  assign t[119] = (x[31]);
  assign t[11] = ~(t[33]);
  assign t[120] = (x[34]);
  assign t[121] = (x[34]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[40]);
  assign t[125] = (x[40]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20] & t[11]);
  assign t[17] = ~(t[34] & t[21]);
  assign t[18] = ~(t[35] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[38] & t[39]);
  assign t[24] = ~(t[40] & t[41]);
  assign t[25] = ~(t[20] & t[26]);
  assign t[26] = t[27] & t[37];
  assign t[27] = ~(t[34] | t[33]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = t[56] ^ x[3];
  assign t[43] = t[57] ^ x[6];
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[12];
  assign t[46] = t[60] ^ x[15];
  assign t[47] = t[61] ^ x[18];
  assign t[48] = t[62] ^ x[21];
  assign t[49] = t[63] ^ x[24];
  assign t[4] = ~(t[9] | t[10]);
  assign t[50] = t[64] ^ x[27];
  assign t[51] = t[65] ^ x[30];
  assign t[52] = t[66] ^ x[33];
  assign t[53] = t[67] ^ x[36];
  assign t[54] = t[68] ^ x[39];
  assign t[55] = t[69] ^ x[42];
  assign t[56] = (t[70] & ~t[71]);
  assign t[57] = (t[72] & ~t[73]);
  assign t[58] = (t[74] & ~t[75]);
  assign t[59] = (t[76] & ~t[77]);
  assign t[5] = ~(t[11] | t[12]);
  assign t[60] = (t[78] & ~t[79]);
  assign t[61] = (t[80] & ~t[81]);
  assign t[62] = (t[82] & ~t[83]);
  assign t[63] = (t[84] & ~t[85]);
  assign t[64] = (t[86] & ~t[87]);
  assign t[65] = (t[88] & ~t[89]);
  assign t[66] = (t[90] & ~t[91]);
  assign t[67] = (t[92] & ~t[93]);
  assign t[68] = (t[94] & ~t[95]);
  assign t[69] = (t[96] & ~t[97]);
  assign t[6] = ~(x[0]);
  assign t[70] = t[98] ^ x[3];
  assign t[71] = t[99] ^ x[2];
  assign t[72] = t[100] ^ x[6];
  assign t[73] = t[101] ^ x[5];
  assign t[74] = t[102] ^ x[9];
  assign t[75] = t[103] ^ x[8];
  assign t[76] = t[104] ^ x[12];
  assign t[77] = t[105] ^ x[11];
  assign t[78] = t[106] ^ x[15];
  assign t[79] = t[107] ^ x[14];
  assign t[7] = ~(t[28] & t[29]);
  assign t[80] = t[108] ^ x[18];
  assign t[81] = t[109] ^ x[17];
  assign t[82] = t[110] ^ x[21];
  assign t[83] = t[111] ^ x[20];
  assign t[84] = t[112] ^ x[24];
  assign t[85] = t[113] ^ x[23];
  assign t[86] = t[114] ^ x[27];
  assign t[87] = t[115] ^ x[26];
  assign t[88] = t[116] ^ x[30];
  assign t[89] = t[117] ^ x[29];
  assign t[8] = ~(t[30] & t[31]);
  assign t[90] = t[118] ^ x[33];
  assign t[91] = t[119] ^ x[32];
  assign t[92] = t[120] ^ x[36];
  assign t[93] = t[121] ^ x[35];
  assign t[94] = t[122] ^ x[39];
  assign t[95] = t[123] ^ x[38];
  assign t[96] = t[124] ^ x[42];
  assign t[97] = t[125] ^ x[41];
  assign t[98] = (x[1]);
  assign t[99] = (x[1]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind7(x, y);
 input [42:0] x;
 output y;

 wire [125:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[4]);
  assign t[101] = (x[4]);
  assign t[102] = (x[7]);
  assign t[103] = (x[7]);
  assign t[104] = (x[10]);
  assign t[105] = (x[10]);
  assign t[106] = (x[13]);
  assign t[107] = (x[13]);
  assign t[108] = (x[16]);
  assign t[109] = (x[16]);
  assign t[10] = ~(t[32] & t[6]);
  assign t[110] = (x[19]);
  assign t[111] = (x[19]);
  assign t[112] = (x[22]);
  assign t[113] = (x[22]);
  assign t[114] = (x[25]);
  assign t[115] = (x[25]);
  assign t[116] = (x[28]);
  assign t[117] = (x[28]);
  assign t[118] = (x[31]);
  assign t[119] = (x[31]);
  assign t[11] = ~(t[33]);
  assign t[120] = (x[34]);
  assign t[121] = (x[34]);
  assign t[122] = (x[37]);
  assign t[123] = (x[37]);
  assign t[124] = (x[40]);
  assign t[125] = (x[40]);
  assign t[12] = ~(t[14] & t[15]);
  assign t[13] = ~(t[16] | t[17]);
  assign t[14] = ~(t[18]);
  assign t[15] = ~(t[19]);
  assign t[16] = ~(t[20] & t[11]);
  assign t[17] = ~(t[34] & t[21]);
  assign t[18] = ~(t[35] | t[22]);
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[36]);
  assign t[21] = ~(t[37]);
  assign t[22] = ~(t[25]);
  assign t[23] = ~(t[38] & t[39]);
  assign t[24] = ~(t[40] & t[41]);
  assign t[25] = ~(t[20] & t[26]);
  assign t[26] = t[27] & t[37];
  assign t[27] = ~(t[34] | t[33]);
  assign t[28] = (t[42]);
  assign t[29] = (t[43]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[44]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7] | t[8]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = t[56] ^ x[3];
  assign t[43] = t[57] ^ x[6];
  assign t[44] = t[58] ^ x[9];
  assign t[45] = t[59] ^ x[12];
  assign t[46] = t[60] ^ x[15];
  assign t[47] = t[61] ^ x[18];
  assign t[48] = t[62] ^ x[21];
  assign t[49] = t[63] ^ x[24];
  assign t[4] = ~(t[9] | t[10]);
  assign t[50] = t[64] ^ x[27];
  assign t[51] = t[65] ^ x[30];
  assign t[52] = t[66] ^ x[33];
  assign t[53] = t[67] ^ x[36];
  assign t[54] = t[68] ^ x[39];
  assign t[55] = t[69] ^ x[42];
  assign t[56] = (t[70] & ~t[71]);
  assign t[57] = (t[72] & ~t[73]);
  assign t[58] = (t[74] & ~t[75]);
  assign t[59] = (t[76] & ~t[77]);
  assign t[5] = ~(t[11] | t[12]);
  assign t[60] = (t[78] & ~t[79]);
  assign t[61] = (t[80] & ~t[81]);
  assign t[62] = (t[82] & ~t[83]);
  assign t[63] = (t[84] & ~t[85]);
  assign t[64] = (t[86] & ~t[87]);
  assign t[65] = (t[88] & ~t[89]);
  assign t[66] = (t[90] & ~t[91]);
  assign t[67] = (t[92] & ~t[93]);
  assign t[68] = (t[94] & ~t[95]);
  assign t[69] = (t[96] & ~t[97]);
  assign t[6] = ~(x[0]);
  assign t[70] = t[98] ^ x[3];
  assign t[71] = t[99] ^ x[2];
  assign t[72] = t[100] ^ x[6];
  assign t[73] = t[101] ^ x[5];
  assign t[74] = t[102] ^ x[9];
  assign t[75] = t[103] ^ x[8];
  assign t[76] = t[104] ^ x[12];
  assign t[77] = t[105] ^ x[11];
  assign t[78] = t[106] ^ x[15];
  assign t[79] = t[107] ^ x[14];
  assign t[7] = ~(t[28] & t[29]);
  assign t[80] = t[108] ^ x[18];
  assign t[81] = t[109] ^ x[17];
  assign t[82] = t[110] ^ x[21];
  assign t[83] = t[111] ^ x[20];
  assign t[84] = t[112] ^ x[24];
  assign t[85] = t[113] ^ x[23];
  assign t[86] = t[114] ^ x[27];
  assign t[87] = t[115] ^ x[26];
  assign t[88] = t[116] ^ x[30];
  assign t[89] = t[117] ^ x[29];
  assign t[8] = ~(t[30] & t[31]);
  assign t[90] = t[118] ^ x[33];
  assign t[91] = t[119] ^ x[32];
  assign t[92] = t[120] ^ x[36];
  assign t[93] = t[121] ^ x[35];
  assign t[94] = t[122] ^ x[39];
  assign t[95] = t[123] ^ x[38];
  assign t[96] = t[124] ^ x[42];
  assign t[97] = t[125] ^ x[41];
  assign t[98] = (x[1]);
  assign t[99] = (x[1]);
  assign t[9] = ~(t[13]);
  assign y = (t[0]);
endmodule

module R2ind8(x, y);
 input [27:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[18] & t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(x[0]);
  assign t[20] = t[29] ^ x[3];
  assign t[21] = t[30] ^ x[6];
  assign t[22] = t[31] ^ x[9];
  assign t[23] = t[32] ^ x[12];
  assign t[24] = t[33] ^ x[15];
  assign t[25] = t[34] ^ x[18];
  assign t[26] = t[35] ^ x[21];
  assign t[27] = t[36] ^ x[24];
  assign t[28] = t[37] ^ x[27];
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (t[40] & ~t[41]);
  assign t[31] = (t[42] & ~t[43]);
  assign t[32] = (t[44] & ~t[45]);
  assign t[33] = (t[46] & ~t[47]);
  assign t[34] = (t[48] & ~t[49]);
  assign t[35] = (t[50] & ~t[51]);
  assign t[36] = (t[52] & ~t[53]);
  assign t[37] = (t[54] & ~t[55]);
  assign t[38] = t[56] ^ x[3];
  assign t[39] = t[57] ^ x[2];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[58] ^ x[6];
  assign t[41] = t[59] ^ x[5];
  assign t[42] = t[60] ^ x[9];
  assign t[43] = t[61] ^ x[8];
  assign t[44] = t[62] ^ x[12];
  assign t[45] = t[63] ^ x[11];
  assign t[46] = t[64] ^ x[15];
  assign t[47] = t[65] ^ x[14];
  assign t[48] = t[66] ^ x[18];
  assign t[49] = t[67] ^ x[17];
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = t[68] ^ x[21];
  assign t[51] = t[69] ^ x[20];
  assign t[52] = t[70] ^ x[24];
  assign t[53] = t[71] ^ x[23];
  assign t[54] = t[72] ^ x[27];
  assign t[55] = t[73] ^ x[26];
  assign t[56] = (x[1]);
  assign t[57] = (x[1]);
  assign t[58] = (x[4]);
  assign t[59] = (x[4]);
  assign t[5] = ~(t[12] | t[13]);
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[10]);
  assign t[63] = (x[10]);
  assign t[64] = (x[13]);
  assign t[65] = (x[13]);
  assign t[66] = (x[16]);
  assign t[67] = (x[16]);
  assign t[68] = (x[19]);
  assign t[69] = (x[19]);
  assign t[6] = ~(t[8] | t[14]);
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[25]);
  assign t[73] = (x[25]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = (t[0]);
endmodule

module R2ind9(x, y);
 input [27:0] x;
 output y;

 wire [73:0] t;
  assign t[0] = t[1] & t[2];
  assign t[10] = ~(t[18] & t[19]);
  assign t[11] = (t[20]);
  assign t[12] = (t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(x[0]);
  assign t[20] = t[29] ^ x[3];
  assign t[21] = t[30] ^ x[6];
  assign t[22] = t[31] ^ x[9];
  assign t[23] = t[32] ^ x[12];
  assign t[24] = t[33] ^ x[15];
  assign t[25] = t[34] ^ x[18];
  assign t[26] = t[35] ^ x[21];
  assign t[27] = t[36] ^ x[24];
  assign t[28] = t[37] ^ x[27];
  assign t[29] = (t[38] & ~t[39]);
  assign t[2] = ~(t[3] & t[4]);
  assign t[30] = (t[40] & ~t[41]);
  assign t[31] = (t[42] & ~t[43]);
  assign t[32] = (t[44] & ~t[45]);
  assign t[33] = (t[46] & ~t[47]);
  assign t[34] = (t[48] & ~t[49]);
  assign t[35] = (t[50] & ~t[51]);
  assign t[36] = (t[52] & ~t[53]);
  assign t[37] = (t[54] & ~t[55]);
  assign t[38] = t[56] ^ x[3];
  assign t[39] = t[57] ^ x[2];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[58] ^ x[6];
  assign t[41] = t[59] ^ x[5];
  assign t[42] = t[60] ^ x[9];
  assign t[43] = t[61] ^ x[8];
  assign t[44] = t[62] ^ x[12];
  assign t[45] = t[63] ^ x[11];
  assign t[46] = t[64] ^ x[15];
  assign t[47] = t[65] ^ x[14];
  assign t[48] = t[66] ^ x[18];
  assign t[49] = t[67] ^ x[17];
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = t[68] ^ x[21];
  assign t[51] = t[69] ^ x[20];
  assign t[52] = t[70] ^ x[24];
  assign t[53] = t[71] ^ x[23];
  assign t[54] = t[72] ^ x[27];
  assign t[55] = t[73] ^ x[26];
  assign t[56] = (x[1]);
  assign t[57] = (x[1]);
  assign t[58] = (x[4]);
  assign t[59] = (x[4]);
  assign t[5] = ~(t[12] | t[13]);
  assign t[60] = (x[7]);
  assign t[61] = (x[7]);
  assign t[62] = (x[10]);
  assign t[63] = (x[10]);
  assign t[64] = (x[13]);
  assign t[65] = (x[13]);
  assign t[66] = (x[16]);
  assign t[67] = (x[16]);
  assign t[68] = (x[19]);
  assign t[69] = (x[19]);
  assign t[6] = ~(t[8] | t[14]);
  assign t[70] = (x[22]);
  assign t[71] = (x[22]);
  assign t[72] = (x[25]);
  assign t[73] = (x[25]);
  assign t[7] = ~(t[9] | t[10]);
  assign t[8] = ~(t[15]);
  assign t[9] = ~(t[16] & t[17]);
  assign y = (t[0]);
endmodule

module R2ind10(x, y);
 input [42:0] x;
 output y;

 wire [128:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[128] ^ x[41];
  assign t[101] = (x[1]);
  assign t[102] = (x[1]);
  assign t[103] = (x[4]);
  assign t[104] = (x[4]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[10]);
  assign t[108] = (x[10]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = (x[13]);
  assign t[111] = (x[16]);
  assign t[112] = (x[16]);
  assign t[113] = (x[19]);
  assign t[114] = (x[19]);
  assign t[115] = (x[22]);
  assign t[116] = (x[22]);
  assign t[117] = (x[25]);
  assign t[118] = (x[25]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[31]);
  assign t[120] = (x[28]);
  assign t[121] = (x[31]);
  assign t[122] = (x[31]);
  assign t[123] = (x[34]);
  assign t[124] = (x[34]);
  assign t[125] = (x[37]);
  assign t[126] = (x[37]);
  assign t[127] = (x[40]);
  assign t[128] = (x[40]);
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[32] | t[21]);
  assign t[14] = ~(t[22] & t[23]);
  assign t[15] = ~(t[33] & t[34]);
  assign t[16] = ~(t[35] & t[36]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[37] & t[8]);
  assign t[19] = ~(t[38] & t[39]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[40] & t[41]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[26] | t[31]);
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[26] & t[29]);
  assign t[26] = ~(t[44]);
  assign t[27] = ~(t[26] & t[30]);
  assign t[28] = ~(t[42] & t[11]);
  assign t[29] = t[22] & t[31];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[43]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = t[59] ^ x[3];
  assign t[46] = t[60] ^ x[6];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[15];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[21];
  assign t[52] = t[66] ^ x[24];
  assign t[53] = t[67] ^ x[27];
  assign t[54] = t[68] ^ x[30];
  assign t[55] = t[69] ^ x[33];
  assign t[56] = t[70] ^ x[36];
  assign t[57] = t[71] ^ x[39];
  assign t[58] = t[72] ^ x[42];
  assign t[59] = (t[73] & ~t[74]);
  assign t[5] = ~(t[11]);
  assign t[60] = (t[75] & ~t[76]);
  assign t[61] = (t[77] & ~t[78]);
  assign t[62] = (t[79] & ~t[80]);
  assign t[63] = (t[81] & ~t[82]);
  assign t[64] = (t[83] & ~t[84]);
  assign t[65] = (t[85] & ~t[86]);
  assign t[66] = (t[87] & ~t[88]);
  assign t[67] = (t[89] & ~t[90]);
  assign t[68] = (t[91] & ~t[92]);
  assign t[69] = (t[93] & ~t[94]);
  assign t[6] = ~(t[12]);
  assign t[70] = (t[95] & ~t[96]);
  assign t[71] = (t[97] & ~t[98]);
  assign t[72] = (t[99] & ~t[100]);
  assign t[73] = t[101] ^ x[3];
  assign t[74] = t[102] ^ x[2];
  assign t[75] = t[103] ^ x[6];
  assign t[76] = t[104] ^ x[5];
  assign t[77] = t[105] ^ x[9];
  assign t[78] = t[106] ^ x[8];
  assign t[79] = t[107] ^ x[12];
  assign t[7] = ~(t[13] & t[14]);
  assign t[80] = t[108] ^ x[11];
  assign t[81] = t[109] ^ x[15];
  assign t[82] = t[110] ^ x[14];
  assign t[83] = t[111] ^ x[18];
  assign t[84] = t[112] ^ x[17];
  assign t[85] = t[113] ^ x[21];
  assign t[86] = t[114] ^ x[20];
  assign t[87] = t[115] ^ x[24];
  assign t[88] = t[116] ^ x[23];
  assign t[89] = t[117] ^ x[27];
  assign t[8] = ~(x[0]);
  assign t[90] = t[118] ^ x[26];
  assign t[91] = t[119] ^ x[30];
  assign t[92] = t[120] ^ x[29];
  assign t[93] = t[121] ^ x[33];
  assign t[94] = t[122] ^ x[32];
  assign t[95] = t[123] ^ x[36];
  assign t[96] = t[124] ^ x[35];
  assign t[97] = t[125] ^ x[39];
  assign t[98] = t[126] ^ x[38];
  assign t[99] = t[127] ^ x[42];
  assign t[9] = ~(t[15] | t[16]);
  assign y = (t[0]);
endmodule

module R2ind11(x, y);
 input [42:0] x;
 output y;

 wire [128:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = t[128] ^ x[41];
  assign t[101] = (x[1]);
  assign t[102] = (x[1]);
  assign t[103] = (x[4]);
  assign t[104] = (x[4]);
  assign t[105] = (x[7]);
  assign t[106] = (x[7]);
  assign t[107] = (x[10]);
  assign t[108] = (x[10]);
  assign t[109] = (x[13]);
  assign t[10] = ~(t[17] | t[18]);
  assign t[110] = (x[13]);
  assign t[111] = (x[16]);
  assign t[112] = (x[16]);
  assign t[113] = (x[19]);
  assign t[114] = (x[19]);
  assign t[115] = (x[22]);
  assign t[116] = (x[22]);
  assign t[117] = (x[25]);
  assign t[118] = (x[25]);
  assign t[119] = (x[28]);
  assign t[11] = ~(t[31]);
  assign t[120] = (x[28]);
  assign t[121] = (x[31]);
  assign t[122] = (x[31]);
  assign t[123] = (x[34]);
  assign t[124] = (x[34]);
  assign t[125] = (x[37]);
  assign t[126] = (x[37]);
  assign t[127] = (x[40]);
  assign t[128] = (x[40]);
  assign t[12] = ~(t[19] | t[20]);
  assign t[13] = ~(t[32] | t[21]);
  assign t[14] = ~(t[22] & t[23]);
  assign t[15] = ~(t[33] & t[34]);
  assign t[16] = ~(t[35] & t[36]);
  assign t[17] = ~(t[24]);
  assign t[18] = ~(t[37] & t[8]);
  assign t[19] = ~(t[38] & t[39]);
  assign t[1] = ~(t[3] & t[4]);
  assign t[20] = ~(t[40] & t[41]);
  assign t[21] = ~(t[25]);
  assign t[22] = ~(t[42] | t[43]);
  assign t[23] = ~(t[26] | t[31]);
  assign t[24] = ~(t[27] | t[28]);
  assign t[25] = ~(t[26] & t[29]);
  assign t[26] = ~(t[44]);
  assign t[27] = ~(t[26] & t[30]);
  assign t[28] = ~(t[42] & t[11]);
  assign t[29] = t[22] & t[31];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = ~(t[43]);
  assign t[31] = (t[45]);
  assign t[32] = (t[46]);
  assign t[33] = (t[47]);
  assign t[34] = (t[48]);
  assign t[35] = (t[49]);
  assign t[36] = (t[50]);
  assign t[37] = (t[51]);
  assign t[38] = (t[52]);
  assign t[39] = (t[53]);
  assign t[3] = ~(t[7] & t[8]);
  assign t[40] = (t[54]);
  assign t[41] = (t[55]);
  assign t[42] = (t[56]);
  assign t[43] = (t[57]);
  assign t[44] = (t[58]);
  assign t[45] = t[59] ^ x[3];
  assign t[46] = t[60] ^ x[6];
  assign t[47] = t[61] ^ x[9];
  assign t[48] = t[62] ^ x[12];
  assign t[49] = t[63] ^ x[15];
  assign t[4] = ~(t[9] & t[10]);
  assign t[50] = t[64] ^ x[18];
  assign t[51] = t[65] ^ x[21];
  assign t[52] = t[66] ^ x[24];
  assign t[53] = t[67] ^ x[27];
  assign t[54] = t[68] ^ x[30];
  assign t[55] = t[69] ^ x[33];
  assign t[56] = t[70] ^ x[36];
  assign t[57] = t[71] ^ x[39];
  assign t[58] = t[72] ^ x[42];
  assign t[59] = (t[73] & ~t[74]);
  assign t[5] = ~(t[11]);
  assign t[60] = (t[75] & ~t[76]);
  assign t[61] = (t[77] & ~t[78]);
  assign t[62] = (t[79] & ~t[80]);
  assign t[63] = (t[81] & ~t[82]);
  assign t[64] = (t[83] & ~t[84]);
  assign t[65] = (t[85] & ~t[86]);
  assign t[66] = (t[87] & ~t[88]);
  assign t[67] = (t[89] & ~t[90]);
  assign t[68] = (t[91] & ~t[92]);
  assign t[69] = (t[93] & ~t[94]);
  assign t[6] = ~(t[12]);
  assign t[70] = (t[95] & ~t[96]);
  assign t[71] = (t[97] & ~t[98]);
  assign t[72] = (t[99] & ~t[100]);
  assign t[73] = t[101] ^ x[3];
  assign t[74] = t[102] ^ x[2];
  assign t[75] = t[103] ^ x[6];
  assign t[76] = t[104] ^ x[5];
  assign t[77] = t[105] ^ x[9];
  assign t[78] = t[106] ^ x[8];
  assign t[79] = t[107] ^ x[12];
  assign t[7] = ~(t[13] & t[14]);
  assign t[80] = t[108] ^ x[11];
  assign t[81] = t[109] ^ x[15];
  assign t[82] = t[110] ^ x[14];
  assign t[83] = t[111] ^ x[18];
  assign t[84] = t[112] ^ x[17];
  assign t[85] = t[113] ^ x[21];
  assign t[86] = t[114] ^ x[20];
  assign t[87] = t[115] ^ x[24];
  assign t[88] = t[116] ^ x[23];
  assign t[89] = t[117] ^ x[27];
  assign t[8] = ~(x[0]);
  assign t[90] = t[118] ^ x[26];
  assign t[91] = t[119] ^ x[30];
  assign t[92] = t[120] ^ x[29];
  assign t[93] = t[121] ^ x[33];
  assign t[94] = t[122] ^ x[32];
  assign t[95] = t[123] ^ x[36];
  assign t[96] = t[124] ^ x[35];
  assign t[97] = t[125] ^ x[39];
  assign t[98] = t[126] ^ x[38];
  assign t[99] = t[127] ^ x[42];
  assign t[9] = ~(t[15] | t[16]);
  assign y = (t[0]);
endmodule

module R2ind12(x, y);
 input [39:0] x;
 output y;

 wire [112:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[19]);
  assign t[101] = (x[22]);
  assign t[102] = (x[22]);
  assign t[103] = (x[25]);
  assign t[104] = (x[25]);
  assign t[105] = (x[28]);
  assign t[106] = (x[28]);
  assign t[107] = (x[31]);
  assign t[108] = (x[31]);
  assign t[109] = (x[34]);
  assign t[10] = ~(t[24]);
  assign t[110] = (x[34]);
  assign t[111] = (x[37]);
  assign t[112] = (x[37]);
  assign t[11] = ~(t[12] & t[25]);
  assign t[12] = t[26] & t[13];
  assign t[13] = ~(t[14] | t[15]);
  assign t[14] = ~(t[16] & t[17]);
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[27]);
  assign t[17] = t[19] & t[28];
  assign t[18] = ~(t[20] | t[21]);
  assign t[19] = ~(t[29] | t[30]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[31] & t[32]);
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = (t[35]);
  assign t[23] = (t[36]);
  assign t[24] = (t[37]);
  assign t[25] = (t[38]);
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = t[22] ? t[5] : t[4];
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = t[48] ^ x[2];
  assign t[36] = t[49] ^ x[6];
  assign t[37] = t[50] ^ x[9];
  assign t[38] = t[51] ^ x[12];
  assign t[39] = t[52] ^ x[15];
  assign t[3] = ~(x[3]);
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[24];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[30];
  assign t[45] = t[58] ^ x[33];
  assign t[46] = t[59] ^ x[36];
  assign t[47] = t[60] ^ x[39];
  assign t[48] = (t[61] & ~t[62]);
  assign t[49] = (t[63] & ~t[64]);
  assign t[4] = t[6] | t[7];
  assign t[50] = (t[65] & ~t[66]);
  assign t[51] = (t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[70]);
  assign t[53] = (t[71] & ~t[72]);
  assign t[54] = (t[73] & ~t[74]);
  assign t[55] = (t[75] & ~t[76]);
  assign t[56] = (t[77] & ~t[78]);
  assign t[57] = (t[79] & ~t[80]);
  assign t[58] = (t[81] & ~t[82]);
  assign t[59] = (t[83] & ~t[84]);
  assign t[5] = ~(t[6] | t[8]);
  assign t[60] = (t[85] & ~t[86]);
  assign t[61] = t[87] ^ x[2];
  assign t[62] = t[88] ^ x[1];
  assign t[63] = t[89] ^ x[6];
  assign t[64] = t[90] ^ x[5];
  assign t[65] = t[91] ^ x[9];
  assign t[66] = t[92] ^ x[8];
  assign t[67] = t[93] ^ x[12];
  assign t[68] = t[94] ^ x[11];
  assign t[69] = t[95] ^ x[15];
  assign t[6] = ~(t[23]);
  assign t[70] = t[96] ^ x[14];
  assign t[71] = t[97] ^ x[18];
  assign t[72] = t[98] ^ x[17];
  assign t[73] = t[99] ^ x[21];
  assign t[74] = t[100] ^ x[20];
  assign t[75] = t[101] ^ x[24];
  assign t[76] = t[102] ^ x[23];
  assign t[77] = t[103] ^ x[27];
  assign t[78] = t[104] ^ x[26];
  assign t[79] = t[105] ^ x[30];
  assign t[7] = ~(t[9] & t[24]);
  assign t[80] = t[106] ^ x[29];
  assign t[81] = t[107] ^ x[33];
  assign t[82] = t[108] ^ x[32];
  assign t[83] = t[109] ^ x[36];
  assign t[84] = t[110] ^ x[35];
  assign t[85] = t[111] ^ x[39];
  assign t[86] = t[112] ^ x[38];
  assign t[87] = (x[0]);
  assign t[88] = (x[0]);
  assign t[89] = (x[4]);
  assign t[8] = t[10] | t[11];
  assign t[90] = (x[4]);
  assign t[91] = (x[7]);
  assign t[92] = (x[7]);
  assign t[93] = (x[10]);
  assign t[94] = (x[10]);
  assign t[95] = (x[13]);
  assign t[96] = (x[13]);
  assign t[97] = (x[16]);
  assign t[98] = (x[16]);
  assign t[99] = (x[19]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind13(x, y);
 input [39:0] x;
 output y;

 wire [112:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[19]);
  assign t[101] = (x[22]);
  assign t[102] = (x[22]);
  assign t[103] = (x[25]);
  assign t[104] = (x[25]);
  assign t[105] = (x[28]);
  assign t[106] = (x[28]);
  assign t[107] = (x[31]);
  assign t[108] = (x[31]);
  assign t[109] = (x[34]);
  assign t[10] = ~(t[24]);
  assign t[110] = (x[34]);
  assign t[111] = (x[37]);
  assign t[112] = (x[37]);
  assign t[11] = ~(t[12] & t[25]);
  assign t[12] = t[26] & t[13];
  assign t[13] = ~(t[14] | t[15]);
  assign t[14] = ~(t[16] & t[17]);
  assign t[15] = ~(t[18]);
  assign t[16] = ~(t[27]);
  assign t[17] = t[19] & t[28];
  assign t[18] = ~(t[20] | t[21]);
  assign t[19] = ~(t[29] | t[30]);
  assign t[1] = ~(t[3]);
  assign t[20] = ~(t[31] & t[32]);
  assign t[21] = ~(t[33] & t[34]);
  assign t[22] = (t[35]);
  assign t[23] = (t[36]);
  assign t[24] = (t[37]);
  assign t[25] = (t[38]);
  assign t[26] = (t[39]);
  assign t[27] = (t[40]);
  assign t[28] = (t[41]);
  assign t[29] = (t[42]);
  assign t[2] = t[22] ? t[5] : t[4];
  assign t[30] = (t[43]);
  assign t[31] = (t[44]);
  assign t[32] = (t[45]);
  assign t[33] = (t[46]);
  assign t[34] = (t[47]);
  assign t[35] = t[48] ^ x[2];
  assign t[36] = t[49] ^ x[6];
  assign t[37] = t[50] ^ x[9];
  assign t[38] = t[51] ^ x[12];
  assign t[39] = t[52] ^ x[15];
  assign t[3] = ~(x[3]);
  assign t[40] = t[53] ^ x[18];
  assign t[41] = t[54] ^ x[21];
  assign t[42] = t[55] ^ x[24];
  assign t[43] = t[56] ^ x[27];
  assign t[44] = t[57] ^ x[30];
  assign t[45] = t[58] ^ x[33];
  assign t[46] = t[59] ^ x[36];
  assign t[47] = t[60] ^ x[39];
  assign t[48] = (t[61] & ~t[62]);
  assign t[49] = (t[63] & ~t[64]);
  assign t[4] = t[6] | t[7];
  assign t[50] = (t[65] & ~t[66]);
  assign t[51] = (t[67] & ~t[68]);
  assign t[52] = (t[69] & ~t[70]);
  assign t[53] = (t[71] & ~t[72]);
  assign t[54] = (t[73] & ~t[74]);
  assign t[55] = (t[75] & ~t[76]);
  assign t[56] = (t[77] & ~t[78]);
  assign t[57] = (t[79] & ~t[80]);
  assign t[58] = (t[81] & ~t[82]);
  assign t[59] = (t[83] & ~t[84]);
  assign t[5] = ~(t[6] | t[8]);
  assign t[60] = (t[85] & ~t[86]);
  assign t[61] = t[87] ^ x[2];
  assign t[62] = t[88] ^ x[1];
  assign t[63] = t[89] ^ x[6];
  assign t[64] = t[90] ^ x[5];
  assign t[65] = t[91] ^ x[9];
  assign t[66] = t[92] ^ x[8];
  assign t[67] = t[93] ^ x[12];
  assign t[68] = t[94] ^ x[11];
  assign t[69] = t[95] ^ x[15];
  assign t[6] = ~(t[23]);
  assign t[70] = t[96] ^ x[14];
  assign t[71] = t[97] ^ x[18];
  assign t[72] = t[98] ^ x[17];
  assign t[73] = t[99] ^ x[21];
  assign t[74] = t[100] ^ x[20];
  assign t[75] = t[101] ^ x[24];
  assign t[76] = t[102] ^ x[23];
  assign t[77] = t[103] ^ x[27];
  assign t[78] = t[104] ^ x[26];
  assign t[79] = t[105] ^ x[30];
  assign t[7] = ~(t[9] & t[24]);
  assign t[80] = t[106] ^ x[29];
  assign t[81] = t[107] ^ x[33];
  assign t[82] = t[108] ^ x[32];
  assign t[83] = t[109] ^ x[36];
  assign t[84] = t[110] ^ x[35];
  assign t[85] = t[111] ^ x[39];
  assign t[86] = t[112] ^ x[38];
  assign t[87] = (x[0]);
  assign t[88] = (x[0]);
  assign t[89] = (x[4]);
  assign t[8] = t[10] | t[11];
  assign t[90] = (x[4]);
  assign t[91] = (x[7]);
  assign t[92] = (x[7]);
  assign t[93] = (x[10]);
  assign t[94] = (x[10]);
  assign t[95] = (x[13]);
  assign t[96] = (x[13]);
  assign t[97] = (x[16]);
  assign t[98] = (x[16]);
  assign t[99] = (x[19]);
  assign t[9] = ~(t[11]);
  assign y = (t[0]);
endmodule

module R2ind14(x, y);
 input [33:0] x;
 output y;

 wire [91:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[12] & t[19];
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = (t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = t[3] ^ t[15];
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = t[37] ^ x[2];
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[9];
  assign t[29] = t[40] ^ x[12];
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] ^ x[15];
  assign t[31] = t[42] ^ x[18];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[24];
  assign t[34] = t[45] ^ x[27];
  assign t[35] = t[46] ^ x[30];
  assign t[36] = t[47] ^ x[33];
  assign t[37] = (t[48] & ~t[49]);
  assign t[38] = (t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[53]);
  assign t[3] = ~(t[5] & t[16]);
  assign t[40] = (t[54] & ~t[55]);
  assign t[41] = (t[56] & ~t[57]);
  assign t[42] = (t[58] & ~t[59]);
  assign t[43] = (t[60] & ~t[61]);
  assign t[44] = (t[62] & ~t[63]);
  assign t[45] = (t[64] & ~t[65]);
  assign t[46] = (t[66] & ~t[67]);
  assign t[47] = (t[68] & ~t[69]);
  assign t[48] = t[70] ^ x[2];
  assign t[49] = t[71] ^ x[1];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[5];
  assign t[51] = t[73] ^ x[4];
  assign t[52] = t[74] ^ x[9];
  assign t[53] = t[75] ^ x[8];
  assign t[54] = t[76] ^ x[12];
  assign t[55] = t[77] ^ x[11];
  assign t[56] = t[78] ^ x[15];
  assign t[57] = t[79] ^ x[14];
  assign t[58] = t[80] ^ x[18];
  assign t[59] = t[81] ^ x[17];
  assign t[5] = t[17] & t[6];
  assign t[60] = t[82] ^ x[21];
  assign t[61] = t[83] ^ x[20];
  assign t[62] = t[84] ^ x[24];
  assign t[63] = t[85] ^ x[23];
  assign t[64] = t[86] ^ x[27];
  assign t[65] = t[87] ^ x[26];
  assign t[66] = t[88] ^ x[30];
  assign t[67] = t[89] ^ x[29];
  assign t[68] = t[90] ^ x[33];
  assign t[69] = t[91] ^ x[32];
  assign t[6] = ~(t[7] | t[8]);
  assign t[70] = (x[0]);
  assign t[71] = (x[0]);
  assign t[72] = (x[3]);
  assign t[73] = (x[3]);
  assign t[74] = (x[7]);
  assign t[75] = (x[7]);
  assign t[76] = (x[10]);
  assign t[77] = (x[10]);
  assign t[78] = (x[13]);
  assign t[79] = (x[13]);
  assign t[7] = ~(t[9] & t[10]);
  assign t[80] = (x[16]);
  assign t[81] = (x[16]);
  assign t[82] = (x[19]);
  assign t[83] = (x[19]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[25]);
  assign t[87] = (x[25]);
  assign t[88] = (x[28]);
  assign t[89] = (x[28]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[31]);
  assign t[91] = (x[31]);
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind15(x, y);
 input [33:0] x;
 output y;

 wire [91:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[12] & t[19];
  assign t[11] = ~(t[13] | t[14]);
  assign t[12] = ~(t[20] | t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = ~(t[24] & t[25]);
  assign t[15] = (t[26]);
  assign t[16] = (t[27]);
  assign t[17] = (t[28]);
  assign t[18] = (t[29]);
  assign t[19] = (t[30]);
  assign t[1] = t[3] ^ t[15];
  assign t[20] = (t[31]);
  assign t[21] = (t[32]);
  assign t[22] = (t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = t[37] ^ x[2];
  assign t[27] = t[38] ^ x[5];
  assign t[28] = t[39] ^ x[9];
  assign t[29] = t[40] ^ x[12];
  assign t[2] = ~(t[4]);
  assign t[30] = t[41] ^ x[15];
  assign t[31] = t[42] ^ x[18];
  assign t[32] = t[43] ^ x[21];
  assign t[33] = t[44] ^ x[24];
  assign t[34] = t[45] ^ x[27];
  assign t[35] = t[46] ^ x[30];
  assign t[36] = t[47] ^ x[33];
  assign t[37] = (t[48] & ~t[49]);
  assign t[38] = (t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[53]);
  assign t[3] = ~(t[5] & t[16]);
  assign t[40] = (t[54] & ~t[55]);
  assign t[41] = (t[56] & ~t[57]);
  assign t[42] = (t[58] & ~t[59]);
  assign t[43] = (t[60] & ~t[61]);
  assign t[44] = (t[62] & ~t[63]);
  assign t[45] = (t[64] & ~t[65]);
  assign t[46] = (t[66] & ~t[67]);
  assign t[47] = (t[68] & ~t[69]);
  assign t[48] = t[70] ^ x[2];
  assign t[49] = t[71] ^ x[1];
  assign t[4] = ~(x[6]);
  assign t[50] = t[72] ^ x[5];
  assign t[51] = t[73] ^ x[4];
  assign t[52] = t[74] ^ x[9];
  assign t[53] = t[75] ^ x[8];
  assign t[54] = t[76] ^ x[12];
  assign t[55] = t[77] ^ x[11];
  assign t[56] = t[78] ^ x[15];
  assign t[57] = t[79] ^ x[14];
  assign t[58] = t[80] ^ x[18];
  assign t[59] = t[81] ^ x[17];
  assign t[5] = t[17] & t[6];
  assign t[60] = t[82] ^ x[21];
  assign t[61] = t[83] ^ x[20];
  assign t[62] = t[84] ^ x[24];
  assign t[63] = t[85] ^ x[23];
  assign t[64] = t[86] ^ x[27];
  assign t[65] = t[87] ^ x[26];
  assign t[66] = t[88] ^ x[30];
  assign t[67] = t[89] ^ x[29];
  assign t[68] = t[90] ^ x[33];
  assign t[69] = t[91] ^ x[32];
  assign t[6] = ~(t[7] | t[8]);
  assign t[70] = (x[0]);
  assign t[71] = (x[0]);
  assign t[72] = (x[3]);
  assign t[73] = (x[3]);
  assign t[74] = (x[7]);
  assign t[75] = (x[7]);
  assign t[76] = (x[10]);
  assign t[77] = (x[10]);
  assign t[78] = (x[13]);
  assign t[79] = (x[13]);
  assign t[7] = ~(t[9] & t[10]);
  assign t[80] = (x[16]);
  assign t[81] = (x[16]);
  assign t[82] = (x[19]);
  assign t[83] = (x[19]);
  assign t[84] = (x[22]);
  assign t[85] = (x[22]);
  assign t[86] = (x[25]);
  assign t[87] = (x[25]);
  assign t[88] = (x[28]);
  assign t[89] = (x[28]);
  assign t[8] = ~(t[11]);
  assign t[90] = (x[31]);
  assign t[91] = (x[31]);
  assign t[9] = ~(t[18]);
  assign y = (t[0]);
endmodule

module R2ind16(x, y);
 input [30:0] x;
 output y;

 wire [83:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = (t[24]);
  assign t[15] = (t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[9];
  assign t[27] = t[37] ^ x[12];
  assign t[28] = t[38] ^ x[15];
  assign t[29] = t[39] ^ x[18];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[24];
  assign t[32] = t[42] ^ x[27];
  assign t[33] = t[43] ^ x[30];
  assign t[34] = (t[44] & ~t[45]);
  assign t[35] = (t[46] & ~t[47]);
  assign t[36] = (t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[51]);
  assign t[38] = (t[52] & ~t[53]);
  assign t[39] = (t[54] & ~t[55]);
  assign t[3] = t[15] & t[5];
  assign t[40] = (t[56] & ~t[57]);
  assign t[41] = (t[58] & ~t[59]);
  assign t[42] = (t[60] & ~t[61]);
  assign t[43] = (t[62] & ~t[63]);
  assign t[44] = t[64] ^ x[2];
  assign t[45] = t[65] ^ x[1];
  assign t[46] = t[66] ^ x[5];
  assign t[47] = t[67] ^ x[4];
  assign t[48] = t[68] ^ x[9];
  assign t[49] = t[69] ^ x[8];
  assign t[4] = ~(x[6]);
  assign t[50] = t[70] ^ x[12];
  assign t[51] = t[71] ^ x[11];
  assign t[52] = t[72] ^ x[15];
  assign t[53] = t[73] ^ x[14];
  assign t[54] = t[74] ^ x[18];
  assign t[55] = t[75] ^ x[17];
  assign t[56] = t[76] ^ x[21];
  assign t[57] = t[77] ^ x[20];
  assign t[58] = t[78] ^ x[24];
  assign t[59] = t[79] ^ x[23];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[80] ^ x[27];
  assign t[61] = t[81] ^ x[26];
  assign t[62] = t[82] ^ x[30];
  assign t[63] = t[83] ^ x[29];
  assign t[64] = (x[0]);
  assign t[65] = (x[0]);
  assign t[66] = (x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[70] = (x[10]);
  assign t[71] = (x[10]);
  assign t[72] = (x[13]);
  assign t[73] = (x[13]);
  assign t[74] = (x[16]);
  assign t[75] = (x[16]);
  assign t[76] = (x[19]);
  assign t[77] = (x[19]);
  assign t[78] = (x[22]);
  assign t[79] = (x[22]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[25]);
  assign t[81] = (x[25]);
  assign t[82] = (x[28]);
  assign t[83] = (x[28]);
  assign t[8] = ~(t[16]);
  assign t[9] = t[11] & t[17];
  assign y = (t[0]);
endmodule

module R2ind17(x, y);
 input [30:0] x;
 output y;

 wire [83:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[18] | t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = ~(t[22] & t[23]);
  assign t[14] = (t[24]);
  assign t[15] = (t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[9];
  assign t[27] = t[37] ^ x[12];
  assign t[28] = t[38] ^ x[15];
  assign t[29] = t[39] ^ x[18];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[21];
  assign t[31] = t[41] ^ x[24];
  assign t[32] = t[42] ^ x[27];
  assign t[33] = t[43] ^ x[30];
  assign t[34] = (t[44] & ~t[45]);
  assign t[35] = (t[46] & ~t[47]);
  assign t[36] = (t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[51]);
  assign t[38] = (t[52] & ~t[53]);
  assign t[39] = (t[54] & ~t[55]);
  assign t[3] = t[15] & t[5];
  assign t[40] = (t[56] & ~t[57]);
  assign t[41] = (t[58] & ~t[59]);
  assign t[42] = (t[60] & ~t[61]);
  assign t[43] = (t[62] & ~t[63]);
  assign t[44] = t[64] ^ x[2];
  assign t[45] = t[65] ^ x[1];
  assign t[46] = t[66] ^ x[5];
  assign t[47] = t[67] ^ x[4];
  assign t[48] = t[68] ^ x[9];
  assign t[49] = t[69] ^ x[8];
  assign t[4] = ~(x[6]);
  assign t[50] = t[70] ^ x[12];
  assign t[51] = t[71] ^ x[11];
  assign t[52] = t[72] ^ x[15];
  assign t[53] = t[73] ^ x[14];
  assign t[54] = t[74] ^ x[18];
  assign t[55] = t[75] ^ x[17];
  assign t[56] = t[76] ^ x[21];
  assign t[57] = t[77] ^ x[20];
  assign t[58] = t[78] ^ x[24];
  assign t[59] = t[79] ^ x[23];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = t[80] ^ x[27];
  assign t[61] = t[81] ^ x[26];
  assign t[62] = t[82] ^ x[30];
  assign t[63] = t[83] ^ x[29];
  assign t[64] = (x[0]);
  assign t[65] = (x[0]);
  assign t[66] = (x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[7]);
  assign t[69] = (x[7]);
  assign t[6] = ~(t[8] & t[9]);
  assign t[70] = (x[10]);
  assign t[71] = (x[10]);
  assign t[72] = (x[13]);
  assign t[73] = (x[13]);
  assign t[74] = (x[16]);
  assign t[75] = (x[16]);
  assign t[76] = (x[19]);
  assign t[77] = (x[19]);
  assign t[78] = (x[22]);
  assign t[79] = (x[22]);
  assign t[7] = ~(t[10]);
  assign t[80] = (x[25]);
  assign t[81] = (x[25]);
  assign t[82] = (x[28]);
  assign t[83] = (x[28]);
  assign t[8] = ~(t[16]);
  assign t[9] = t[11] & t[17];
  assign y = (t[0]);
endmodule

module R2ind18(x, y);
 input [27:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = ~(t[18] & t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[13] ^ t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = t[31] ^ x[2];
  assign t[23] = t[32] ^ x[6];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[15];
  assign t[27] = t[36] ^ x[18];
  assign t[28] = t[37] ^ x[21];
  assign t[29] = t[38] ^ x[24];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[27];
  assign t[31] = (t[40] & ~t[41]);
  assign t[32] = (t[42] & ~t[43]);
  assign t[33] = (t[44] & ~t[45]);
  assign t[34] = (t[46] & ~t[47]);
  assign t[35] = (t[48] & ~t[49]);
  assign t[36] = (t[50] & ~t[51]);
  assign t[37] = (t[52] & ~t[53]);
  assign t[38] = (t[54] & ~t[55]);
  assign t[39] = (t[56] & ~t[57]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[58] ^ x[2];
  assign t[41] = t[59] ^ x[1];
  assign t[42] = t[60] ^ x[6];
  assign t[43] = t[61] ^ x[5];
  assign t[44] = t[62] ^ x[9];
  assign t[45] = t[63] ^ x[8];
  assign t[46] = t[64] ^ x[12];
  assign t[47] = t[65] ^ x[11];
  assign t[48] = t[66] ^ x[15];
  assign t[49] = t[67] ^ x[14];
  assign t[4] = ~(x[3]);
  assign t[50] = t[68] ^ x[18];
  assign t[51] = t[69] ^ x[17];
  assign t[52] = t[70] ^ x[21];
  assign t[53] = t[71] ^ x[20];
  assign t[54] = t[72] ^ x[24];
  assign t[55] = t[73] ^ x[23];
  assign t[56] = t[74] ^ x[27];
  assign t[57] = t[75] ^ x[26];
  assign t[58] = (x[0]);
  assign t[59] = (x[0]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4]);
  assign t[61] = (x[4]);
  assign t[62] = (x[7]);
  assign t[63] = (x[7]);
  assign t[64] = (x[10]);
  assign t[65] = (x[10]);
  assign t[66] = (x[13]);
  assign t[67] = (x[13]);
  assign t[68] = (x[16]);
  assign t[69] = (x[16]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[19]);
  assign t[71] = (x[19]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[74] = (x[25]);
  assign t[75] = (x[25]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[10] & t[15];
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind19(x, y);
 input [27:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[16] | t[17]);
  assign t[11] = ~(t[18] & t[19]);
  assign t[12] = ~(t[20] & t[21]);
  assign t[13] = (t[22]);
  assign t[14] = (t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[13] ^ t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = t[31] ^ x[2];
  assign t[23] = t[32] ^ x[6];
  assign t[24] = t[33] ^ x[9];
  assign t[25] = t[34] ^ x[12];
  assign t[26] = t[35] ^ x[15];
  assign t[27] = t[36] ^ x[18];
  assign t[28] = t[37] ^ x[21];
  assign t[29] = t[38] ^ x[24];
  assign t[2] = ~(t[4]);
  assign t[30] = t[39] ^ x[27];
  assign t[31] = (t[40] & ~t[41]);
  assign t[32] = (t[42] & ~t[43]);
  assign t[33] = (t[44] & ~t[45]);
  assign t[34] = (t[46] & ~t[47]);
  assign t[35] = (t[48] & ~t[49]);
  assign t[36] = (t[50] & ~t[51]);
  assign t[37] = (t[52] & ~t[53]);
  assign t[38] = (t[54] & ~t[55]);
  assign t[39] = (t[56] & ~t[57]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[58] ^ x[2];
  assign t[41] = t[59] ^ x[1];
  assign t[42] = t[60] ^ x[6];
  assign t[43] = t[61] ^ x[5];
  assign t[44] = t[62] ^ x[9];
  assign t[45] = t[63] ^ x[8];
  assign t[46] = t[64] ^ x[12];
  assign t[47] = t[65] ^ x[11];
  assign t[48] = t[66] ^ x[15];
  assign t[49] = t[67] ^ x[14];
  assign t[4] = ~(x[3]);
  assign t[50] = t[68] ^ x[18];
  assign t[51] = t[69] ^ x[17];
  assign t[52] = t[70] ^ x[21];
  assign t[53] = t[71] ^ x[20];
  assign t[54] = t[72] ^ x[24];
  assign t[55] = t[73] ^ x[23];
  assign t[56] = t[74] ^ x[27];
  assign t[57] = t[75] ^ x[26];
  assign t[58] = (x[0]);
  assign t[59] = (x[0]);
  assign t[5] = ~(t[7] & t[8]);
  assign t[60] = (x[4]);
  assign t[61] = (x[4]);
  assign t[62] = (x[7]);
  assign t[63] = (x[7]);
  assign t[64] = (x[10]);
  assign t[65] = (x[10]);
  assign t[66] = (x[13]);
  assign t[67] = (x[13]);
  assign t[68] = (x[16]);
  assign t[69] = (x[16]);
  assign t[6] = ~(t[9]);
  assign t[70] = (x[19]);
  assign t[71] = (x[19]);
  assign t[72] = (x[22]);
  assign t[73] = (x[22]);
  assign t[74] = (x[25]);
  assign t[75] = (x[25]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[10] & t[15];
  assign t[9] = ~(t[11] | t[12]);
  assign y = (t[0]);
endmodule

module R2ind20(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[34]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[21]);
  assign t[12] = t[14] & t[22];
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[23] | t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = t[3] ^ t[17];
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = t[41] ^ x[2];
  assign t[2] = ~(t[4]);
  assign t[30] = t[42] ^ x[6];
  assign t[31] = t[43] ^ x[9];
  assign t[32] = t[44] ^ x[12];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[18];
  assign t[35] = t[47] ^ x[21];
  assign t[36] = t[48] ^ x[24];
  assign t[37] = t[49] ^ x[27];
  assign t[38] = t[50] ^ x[30];
  assign t[39] = t[51] ^ x[33];
  assign t[3] = t[5] | t[6];
  assign t[40] = t[52] ^ x[36];
  assign t[41] = (t[53] & ~t[54]);
  assign t[42] = (t[55] & ~t[56]);
  assign t[43] = (t[57] & ~t[58]);
  assign t[44] = (t[59] & ~t[60]);
  assign t[45] = (t[61] & ~t[62]);
  assign t[46] = (t[63] & ~t[64]);
  assign t[47] = (t[65] & ~t[66]);
  assign t[48] = (t[67] & ~t[68]);
  assign t[49] = (t[69] & ~t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = (t[71] & ~t[72]);
  assign t[51] = (t[73] & ~t[74]);
  assign t[52] = (t[75] & ~t[76]);
  assign t[53] = t[77] ^ x[2];
  assign t[54] = t[78] ^ x[1];
  assign t[55] = t[79] ^ x[6];
  assign t[56] = t[80] ^ x[5];
  assign t[57] = t[81] ^ x[9];
  assign t[58] = t[82] ^ x[8];
  assign t[59] = t[83] ^ x[12];
  assign t[5] = ~(t[18]);
  assign t[60] = t[84] ^ x[11];
  assign t[61] = t[85] ^ x[15];
  assign t[62] = t[86] ^ x[14];
  assign t[63] = t[87] ^ x[18];
  assign t[64] = t[88] ^ x[17];
  assign t[65] = t[89] ^ x[21];
  assign t[66] = t[90] ^ x[20];
  assign t[67] = t[91] ^ x[24];
  assign t[68] = t[92] ^ x[23];
  assign t[69] = t[93] ^ x[27];
  assign t[6] = ~(t[7] & t[19]);
  assign t[70] = t[94] ^ x[26];
  assign t[71] = t[95] ^ x[30];
  assign t[72] = t[96] ^ x[29];
  assign t[73] = t[97] ^ x[33];
  assign t[74] = t[98] ^ x[32];
  assign t[75] = t[99] ^ x[36];
  assign t[76] = t[100] ^ x[35];
  assign t[77] = (x[0]);
  assign t[78] = (x[0]);
  assign t[79] = (x[4]);
  assign t[7] = t[20] & t[8];
  assign t[80] = (x[4]);
  assign t[81] = (x[7]);
  assign t[82] = (x[7]);
  assign t[83] = (x[10]);
  assign t[84] = (x[10]);
  assign t[85] = (x[13]);
  assign t[86] = (x[13]);
  assign t[87] = (x[16]);
  assign t[88] = (x[16]);
  assign t[89] = (x[19]);
  assign t[8] = ~(t[9] | t[10]);
  assign t[90] = (x[19]);
  assign t[91] = (x[22]);
  assign t[92] = (x[22]);
  assign t[93] = (x[25]);
  assign t[94] = (x[25]);
  assign t[95] = (x[28]);
  assign t[96] = (x[28]);
  assign t[97] = (x[31]);
  assign t[98] = (x[31]);
  assign t[99] = (x[34]);
  assign t[9] = ~(t[11] & t[12]);
  assign y = (t[0]);
endmodule

module R2ind21(x, y);
 input [36:0] x;
 output y;

 wire [100:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[100] = (x[34]);
  assign t[10] = ~(t[13]);
  assign t[11] = ~(t[21]);
  assign t[12] = t[14] & t[22];
  assign t[13] = ~(t[15] | t[16]);
  assign t[14] = ~(t[23] | t[24]);
  assign t[15] = ~(t[25] & t[26]);
  assign t[16] = ~(t[27] & t[28]);
  assign t[17] = (t[29]);
  assign t[18] = (t[30]);
  assign t[19] = (t[31]);
  assign t[1] = t[3] ^ t[17];
  assign t[20] = (t[32]);
  assign t[21] = (t[33]);
  assign t[22] = (t[34]);
  assign t[23] = (t[35]);
  assign t[24] = (t[36]);
  assign t[25] = (t[37]);
  assign t[26] = (t[38]);
  assign t[27] = (t[39]);
  assign t[28] = (t[40]);
  assign t[29] = t[41] ^ x[2];
  assign t[2] = ~(t[4]);
  assign t[30] = t[42] ^ x[6];
  assign t[31] = t[43] ^ x[9];
  assign t[32] = t[44] ^ x[12];
  assign t[33] = t[45] ^ x[15];
  assign t[34] = t[46] ^ x[18];
  assign t[35] = t[47] ^ x[21];
  assign t[36] = t[48] ^ x[24];
  assign t[37] = t[49] ^ x[27];
  assign t[38] = t[50] ^ x[30];
  assign t[39] = t[51] ^ x[33];
  assign t[3] = t[5] | t[6];
  assign t[40] = t[52] ^ x[36];
  assign t[41] = (t[53] & ~t[54]);
  assign t[42] = (t[55] & ~t[56]);
  assign t[43] = (t[57] & ~t[58]);
  assign t[44] = (t[59] & ~t[60]);
  assign t[45] = (t[61] & ~t[62]);
  assign t[46] = (t[63] & ~t[64]);
  assign t[47] = (t[65] & ~t[66]);
  assign t[48] = (t[67] & ~t[68]);
  assign t[49] = (t[69] & ~t[70]);
  assign t[4] = ~(x[3]);
  assign t[50] = (t[71] & ~t[72]);
  assign t[51] = (t[73] & ~t[74]);
  assign t[52] = (t[75] & ~t[76]);
  assign t[53] = t[77] ^ x[2];
  assign t[54] = t[78] ^ x[1];
  assign t[55] = t[79] ^ x[6];
  assign t[56] = t[80] ^ x[5];
  assign t[57] = t[81] ^ x[9];
  assign t[58] = t[82] ^ x[8];
  assign t[59] = t[83] ^ x[12];
  assign t[5] = ~(t[18]);
  assign t[60] = t[84] ^ x[11];
  assign t[61] = t[85] ^ x[15];
  assign t[62] = t[86] ^ x[14];
  assign t[63] = t[87] ^ x[18];
  assign t[64] = t[88] ^ x[17];
  assign t[65] = t[89] ^ x[21];
  assign t[66] = t[90] ^ x[20];
  assign t[67] = t[91] ^ x[24];
  assign t[68] = t[92] ^ x[23];
  assign t[69] = t[93] ^ x[27];
  assign t[6] = ~(t[7] & t[19]);
  assign t[70] = t[94] ^ x[26];
  assign t[71] = t[95] ^ x[30];
  assign t[72] = t[96] ^ x[29];
  assign t[73] = t[97] ^ x[33];
  assign t[74] = t[98] ^ x[32];
  assign t[75] = t[99] ^ x[36];
  assign t[76] = t[100] ^ x[35];
  assign t[77] = (x[0]);
  assign t[78] = (x[0]);
  assign t[79] = (x[4]);
  assign t[7] = t[20] & t[8];
  assign t[80] = (x[4]);
  assign t[81] = (x[7]);
  assign t[82] = (x[7]);
  assign t[83] = (x[10]);
  assign t[84] = (x[10]);
  assign t[85] = (x[13]);
  assign t[86] = (x[13]);
  assign t[87] = (x[16]);
  assign t[88] = (x[16]);
  assign t[89] = (x[19]);
  assign t[8] = ~(t[9] | t[10]);
  assign t[90] = (x[19]);
  assign t[91] = (x[22]);
  assign t[92] = (x[22]);
  assign t[93] = (x[25]);
  assign t[94] = (x[25]);
  assign t[95] = (x[28]);
  assign t[96] = (x[28]);
  assign t[97] = (x[31]);
  assign t[98] = (x[31]);
  assign t[99] = (x[34]);
  assign t[9] = ~(t[11] & t[12]);
  assign y = (t[0]);
endmodule

module R2ind22(x, y);
 input [26:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[20]);
  assign t[13] = t[14] & t[21];
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[17];
  assign t[2] = t[15] ^ t[4];
  assign t[30] = t[39] ^ x[20];
  assign t[31] = t[40] ^ x[23];
  assign t[32] = t[41] ^ x[26];
  assign t[33] = (t[42] & ~t[43]);
  assign t[34] = (t[44] & ~t[45]);
  assign t[35] = (t[46] & ~t[47]);
  assign t[36] = (t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[51]);
  assign t[38] = (t[52] & ~t[53]);
  assign t[39] = (t[54] & ~t[55]);
  assign t[3] = ~(t[16]);
  assign t[40] = (t[56] & ~t[57]);
  assign t[41] = (t[58] & ~t[59]);
  assign t[42] = t[60] ^ x[2];
  assign t[43] = t[61] ^ x[1];
  assign t[44] = t[62] ^ x[5];
  assign t[45] = t[63] ^ x[4];
  assign t[46] = t[64] ^ x[8];
  assign t[47] = t[65] ^ x[7];
  assign t[48] = t[66] ^ x[11];
  assign t[49] = t[67] ^ x[10];
  assign t[4] = ~(t[5] & t[17]);
  assign t[50] = t[68] ^ x[14];
  assign t[51] = t[69] ^ x[13];
  assign t[52] = t[70] ^ x[17];
  assign t[53] = t[71] ^ x[16];
  assign t[54] = t[72] ^ x[20];
  assign t[55] = t[73] ^ x[19];
  assign t[56] = t[74] ^ x[23];
  assign t[57] = t[75] ^ x[22];
  assign t[58] = t[76] ^ x[26];
  assign t[59] = t[77] ^ x[25];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[0]);
  assign t[61] = (x[0]);
  assign t[62] = (x[3]);
  assign t[63] = (x[3]);
  assign t[64] = (x[6]);
  assign t[65] = (x[6]);
  assign t[66] = (x[9]);
  assign t[67] = (x[9]);
  assign t[68] = (x[12]);
  assign t[69] = (x[12]);
  assign t[6] = ~(t[18]);
  assign t[70] = (x[15]);
  assign t[71] = (x[15]);
  assign t[72] = (x[18]);
  assign t[73] = (x[18]);
  assign t[74] = (x[21]);
  assign t[75] = (x[21]);
  assign t[76] = (x[24]);
  assign t[77] = (x[24]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[19] | t[10]);
  assign y = (t[0]);
endmodule

module R2ind23(x, y);
 input [26:0] x;
 output y;

 wire [77:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11]);
  assign t[11] = ~(t[12] & t[13]);
  assign t[12] = ~(t[20]);
  assign t[13] = t[14] & t[21];
  assign t[14] = ~(t[22] | t[23]);
  assign t[15] = (t[24]);
  assign t[16] = (t[25]);
  assign t[17] = (t[26]);
  assign t[18] = (t[27]);
  assign t[19] = (t[28]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[29]);
  assign t[21] = (t[30]);
  assign t[22] = (t[31]);
  assign t[23] = (t[32]);
  assign t[24] = t[33] ^ x[2];
  assign t[25] = t[34] ^ x[5];
  assign t[26] = t[35] ^ x[8];
  assign t[27] = t[36] ^ x[11];
  assign t[28] = t[37] ^ x[14];
  assign t[29] = t[38] ^ x[17];
  assign t[2] = t[15] ^ t[4];
  assign t[30] = t[39] ^ x[20];
  assign t[31] = t[40] ^ x[23];
  assign t[32] = t[41] ^ x[26];
  assign t[33] = (t[42] & ~t[43]);
  assign t[34] = (t[44] & ~t[45]);
  assign t[35] = (t[46] & ~t[47]);
  assign t[36] = (t[48] & ~t[49]);
  assign t[37] = (t[50] & ~t[51]);
  assign t[38] = (t[52] & ~t[53]);
  assign t[39] = (t[54] & ~t[55]);
  assign t[3] = ~(t[16]);
  assign t[40] = (t[56] & ~t[57]);
  assign t[41] = (t[58] & ~t[59]);
  assign t[42] = t[60] ^ x[2];
  assign t[43] = t[61] ^ x[1];
  assign t[44] = t[62] ^ x[5];
  assign t[45] = t[63] ^ x[4];
  assign t[46] = t[64] ^ x[8];
  assign t[47] = t[65] ^ x[7];
  assign t[48] = t[66] ^ x[11];
  assign t[49] = t[67] ^ x[10];
  assign t[4] = ~(t[5] & t[17]);
  assign t[50] = t[68] ^ x[14];
  assign t[51] = t[69] ^ x[13];
  assign t[52] = t[70] ^ x[17];
  assign t[53] = t[71] ^ x[16];
  assign t[54] = t[72] ^ x[20];
  assign t[55] = t[73] ^ x[19];
  assign t[56] = t[74] ^ x[23];
  assign t[57] = t[75] ^ x[22];
  assign t[58] = t[76] ^ x[26];
  assign t[59] = t[77] ^ x[25];
  assign t[5] = ~(t[6] | t[7]);
  assign t[60] = (x[0]);
  assign t[61] = (x[0]);
  assign t[62] = (x[3]);
  assign t[63] = (x[3]);
  assign t[64] = (x[6]);
  assign t[65] = (x[6]);
  assign t[66] = (x[9]);
  assign t[67] = (x[9]);
  assign t[68] = (x[12]);
  assign t[69] = (x[12]);
  assign t[6] = ~(t[18]);
  assign t[70] = (x[15]);
  assign t[71] = (x[15]);
  assign t[72] = (x[18]);
  assign t[73] = (x[18]);
  assign t[74] = (x[21]);
  assign t[75] = (x[21]);
  assign t[76] = (x[24]);
  assign t[77] = (x[24]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(t[19] | t[10]);
  assign y = (t[0]);
endmodule

module R2ind24(x, y);
 input [29:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11]);
  assign t[11] = ~(t[22] | t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[23]);
  assign t[15] = t[16] & t[24];
  assign t[16] = ~(t[25] | t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[17] ^ t[3]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = t[37] ^ x[2];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[20];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[29];
  assign t[37] = (t[47] & ~t[48]);
  assign t[38] = (t[49] & ~t[50]);
  assign t[39] = (t[51] & ~t[52]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = (t[53] & ~t[54]);
  assign t[41] = (t[55] & ~t[56]);
  assign t[42] = (t[57] & ~t[58]);
  assign t[43] = (t[59] & ~t[60]);
  assign t[44] = (t[61] & ~t[62]);
  assign t[45] = (t[63] & ~t[64]);
  assign t[46] = (t[65] & ~t[66]);
  assign t[47] = t[67] ^ x[2];
  assign t[48] = t[68] ^ x[1];
  assign t[49] = t[69] ^ x[5];
  assign t[4] = ~(t[18]);
  assign t[50] = t[70] ^ x[4];
  assign t[51] = t[71] ^ x[8];
  assign t[52] = t[72] ^ x[7];
  assign t[53] = t[73] ^ x[11];
  assign t[54] = t[74] ^ x[10];
  assign t[55] = t[75] ^ x[14];
  assign t[56] = t[76] ^ x[13];
  assign t[57] = t[77] ^ x[17];
  assign t[58] = t[78] ^ x[16];
  assign t[59] = t[79] ^ x[20];
  assign t[5] = ~(t[19]);
  assign t[60] = t[80] ^ x[19];
  assign t[61] = t[81] ^ x[23];
  assign t[62] = t[82] ^ x[22];
  assign t[63] = t[83] ^ x[26];
  assign t[64] = t[84] ^ x[25];
  assign t[65] = t[85] ^ x[29];
  assign t[66] = t[86] ^ x[28];
  assign t[67] = (x[0]);
  assign t[68] = (x[0]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[7] & t[20]);
  assign t[70] = (x[3]);
  assign t[71] = (x[6]);
  assign t[72] = (x[6]);
  assign t[73] = (x[9]);
  assign t[74] = (x[9]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[15]);
  assign t[78] = (x[15]);
  assign t[79] = (x[18]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21]);
  assign t[82] = (x[21]);
  assign t[83] = (x[24]);
  assign t[84] = (x[24]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = ~(t[21]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind25(x, y);
 input [29:0] x;
 output y;

 wire [86:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11]);
  assign t[11] = ~(t[22] | t[12]);
  assign t[12] = ~(t[13]);
  assign t[13] = ~(t[14] & t[15]);
  assign t[14] = ~(t[23]);
  assign t[15] = t[16] & t[24];
  assign t[16] = ~(t[25] | t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = ~(t[17] ^ t[3]);
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = (t[36]);
  assign t[27] = t[37] ^ x[2];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[4]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[14];
  assign t[32] = t[42] ^ x[17];
  assign t[33] = t[43] ^ x[20];
  assign t[34] = t[44] ^ x[23];
  assign t[35] = t[45] ^ x[26];
  assign t[36] = t[46] ^ x[29];
  assign t[37] = (t[47] & ~t[48]);
  assign t[38] = (t[49] & ~t[50]);
  assign t[39] = (t[51] & ~t[52]);
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = (t[53] & ~t[54]);
  assign t[41] = (t[55] & ~t[56]);
  assign t[42] = (t[57] & ~t[58]);
  assign t[43] = (t[59] & ~t[60]);
  assign t[44] = (t[61] & ~t[62]);
  assign t[45] = (t[63] & ~t[64]);
  assign t[46] = (t[65] & ~t[66]);
  assign t[47] = t[67] ^ x[2];
  assign t[48] = t[68] ^ x[1];
  assign t[49] = t[69] ^ x[5];
  assign t[4] = ~(t[18]);
  assign t[50] = t[70] ^ x[4];
  assign t[51] = t[71] ^ x[8];
  assign t[52] = t[72] ^ x[7];
  assign t[53] = t[73] ^ x[11];
  assign t[54] = t[74] ^ x[10];
  assign t[55] = t[75] ^ x[14];
  assign t[56] = t[76] ^ x[13];
  assign t[57] = t[77] ^ x[17];
  assign t[58] = t[78] ^ x[16];
  assign t[59] = t[79] ^ x[20];
  assign t[5] = ~(t[19]);
  assign t[60] = t[80] ^ x[19];
  assign t[61] = t[81] ^ x[23];
  assign t[62] = t[82] ^ x[22];
  assign t[63] = t[83] ^ x[26];
  assign t[64] = t[84] ^ x[25];
  assign t[65] = t[85] ^ x[29];
  assign t[66] = t[86] ^ x[28];
  assign t[67] = (x[0]);
  assign t[68] = (x[0]);
  assign t[69] = (x[3]);
  assign t[6] = ~(t[7] & t[20]);
  assign t[70] = (x[3]);
  assign t[71] = (x[6]);
  assign t[72] = (x[6]);
  assign t[73] = (x[9]);
  assign t[74] = (x[9]);
  assign t[75] = (x[12]);
  assign t[76] = (x[12]);
  assign t[77] = (x[15]);
  assign t[78] = (x[15]);
  assign t[79] = (x[18]);
  assign t[7] = ~(t[8] | t[9]);
  assign t[80] = (x[18]);
  assign t[81] = (x[21]);
  assign t[82] = (x[21]);
  assign t[83] = (x[24]);
  assign t[84] = (x[24]);
  assign t[85] = (x[27]);
  assign t[86] = (x[27]);
  assign t[8] = ~(t[21]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind26(x, y);
 input [23:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[18]);
  assign t[12] = t[13] & t[19];
  assign t[13] = ~(t[20] | t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[14];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[20];
  assign t[29] = t[37] ^ x[23];
  assign t[2] = ~(t[4]);
  assign t[30] = (t[38] & ~t[39]);
  assign t[31] = (t[40] & ~t[41]);
  assign t[32] = (t[42] & ~t[43]);
  assign t[33] = (t[44] & ~t[45]);
  assign t[34] = (t[46] & ~t[47]);
  assign t[35] = (t[48] & ~t[49]);
  assign t[36] = (t[50] & ~t[51]);
  assign t[37] = (t[52] & ~t[53]);
  assign t[38] = t[54] ^ x[2];
  assign t[39] = t[55] ^ x[1];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[56] ^ x[5];
  assign t[41] = t[57] ^ x[4];
  assign t[42] = t[58] ^ x[8];
  assign t[43] = t[59] ^ x[7];
  assign t[44] = t[60] ^ x[11];
  assign t[45] = t[61] ^ x[10];
  assign t[46] = t[62] ^ x[14];
  assign t[47] = t[63] ^ x[13];
  assign t[48] = t[64] ^ x[17];
  assign t[49] = t[65] ^ x[16];
  assign t[4] = ~(t[15]);
  assign t[50] = t[66] ^ x[20];
  assign t[51] = t[67] ^ x[19];
  assign t[52] = t[68] ^ x[23];
  assign t[53] = t[69] ^ x[22];
  assign t[54] = (x[0]);
  assign t[55] = (x[0]);
  assign t[56] = (x[3]);
  assign t[57] = (x[3]);
  assign t[58] = (x[6]);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[16]);
  assign t[60] = (x[9]);
  assign t[61] = (x[9]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[15]);
  assign t[65] = (x[15]);
  assign t[66] = (x[18]);
  assign t[67] = (x[18]);
  assign t[68] = (x[21]);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[17] | t[9]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind27(x, y);
 input [23:0] x;
 output y;

 wire [69:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = ~(t[11] & t[12]);
  assign t[11] = ~(t[18]);
  assign t[12] = t[13] & t[19];
  assign t[13] = ~(t[20] | t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = ~(t[3] ^ t[14]);
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[5];
  assign t[24] = t[32] ^ x[8];
  assign t[25] = t[33] ^ x[11];
  assign t[26] = t[34] ^ x[14];
  assign t[27] = t[35] ^ x[17];
  assign t[28] = t[36] ^ x[20];
  assign t[29] = t[37] ^ x[23];
  assign t[2] = ~(t[4]);
  assign t[30] = (t[38] & ~t[39]);
  assign t[31] = (t[40] & ~t[41]);
  assign t[32] = (t[42] & ~t[43]);
  assign t[33] = (t[44] & ~t[45]);
  assign t[34] = (t[46] & ~t[47]);
  assign t[35] = (t[48] & ~t[49]);
  assign t[36] = (t[50] & ~t[51]);
  assign t[37] = (t[52] & ~t[53]);
  assign t[38] = t[54] ^ x[2];
  assign t[39] = t[55] ^ x[1];
  assign t[3] = ~(t[5] | t[6]);
  assign t[40] = t[56] ^ x[5];
  assign t[41] = t[57] ^ x[4];
  assign t[42] = t[58] ^ x[8];
  assign t[43] = t[59] ^ x[7];
  assign t[44] = t[60] ^ x[11];
  assign t[45] = t[61] ^ x[10];
  assign t[46] = t[62] ^ x[14];
  assign t[47] = t[63] ^ x[13];
  assign t[48] = t[64] ^ x[17];
  assign t[49] = t[65] ^ x[16];
  assign t[4] = ~(t[15]);
  assign t[50] = t[66] ^ x[20];
  assign t[51] = t[67] ^ x[19];
  assign t[52] = t[68] ^ x[23];
  assign t[53] = t[69] ^ x[22];
  assign t[54] = (x[0]);
  assign t[55] = (x[0]);
  assign t[56] = (x[3]);
  assign t[57] = (x[3]);
  assign t[58] = (x[6]);
  assign t[59] = (x[6]);
  assign t[5] = ~(t[16]);
  assign t[60] = (x[9]);
  assign t[61] = (x[9]);
  assign t[62] = (x[12]);
  assign t[63] = (x[12]);
  assign t[64] = (x[15]);
  assign t[65] = (x[15]);
  assign t[66] = (x[18]);
  assign t[67] = (x[18]);
  assign t[68] = (x[21]);
  assign t[69] = (x[21]);
  assign t[6] = ~(t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[17] | t[9]);
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind28(x, y);
 input [20:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[11] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = t[26] ^ x[2];
  assign t[1] = ~(t[3]);
  assign t[20] = t[27] ^ x[5];
  assign t[21] = t[28] ^ x[8];
  assign t[22] = t[29] ^ x[11];
  assign t[23] = t[30] ^ x[14];
  assign t[24] = t[31] ^ x[17];
  assign t[25] = t[32] ^ x[20];
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = (t[39] & ~t[40]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (t[41] & ~t[42]);
  assign t[31] = (t[43] & ~t[44]);
  assign t[32] = (t[45] & ~t[46]);
  assign t[33] = t[47] ^ x[2];
  assign t[34] = t[48] ^ x[1];
  assign t[35] = t[49] ^ x[5];
  assign t[36] = t[50] ^ x[4];
  assign t[37] = t[51] ^ x[8];
  assign t[38] = t[52] ^ x[7];
  assign t[39] = t[53] ^ x[11];
  assign t[3] = ~(t[12]);
  assign t[40] = t[54] ^ x[10];
  assign t[41] = t[55] ^ x[14];
  assign t[42] = t[56] ^ x[13];
  assign t[43] = t[57] ^ x[17];
  assign t[44] = t[58] ^ x[16];
  assign t[45] = t[59] ^ x[20];
  assign t[46] = t[60] ^ x[19];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = ~(t[13]);
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[55] = (x[12]);
  assign t[56] = (x[12]);
  assign t[57] = (x[15]);
  assign t[58] = (x[15]);
  assign t[59] = (x[18]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[18]);
  assign t[6] = ~(t[14] | t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind29(x, y);
 input [20:0] x;
 output y;

 wire [60:0] t;
  assign t[0] = ~(t[1] | t[2]);
  assign t[10] = t[11] & t[16];
  assign t[11] = ~(t[17] | t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = (t[22]);
  assign t[16] = (t[23]);
  assign t[17] = (t[24]);
  assign t[18] = (t[25]);
  assign t[19] = t[26] ^ x[2];
  assign t[1] = ~(t[3]);
  assign t[20] = t[27] ^ x[5];
  assign t[21] = t[28] ^ x[8];
  assign t[22] = t[29] ^ x[11];
  assign t[23] = t[30] ^ x[14];
  assign t[24] = t[31] ^ x[17];
  assign t[25] = t[32] ^ x[20];
  assign t[26] = (t[33] & ~t[34]);
  assign t[27] = (t[35] & ~t[36]);
  assign t[28] = (t[37] & ~t[38]);
  assign t[29] = (t[39] & ~t[40]);
  assign t[2] = t[4] ^ t[5];
  assign t[30] = (t[41] & ~t[42]);
  assign t[31] = (t[43] & ~t[44]);
  assign t[32] = (t[45] & ~t[46]);
  assign t[33] = t[47] ^ x[2];
  assign t[34] = t[48] ^ x[1];
  assign t[35] = t[49] ^ x[5];
  assign t[36] = t[50] ^ x[4];
  assign t[37] = t[51] ^ x[8];
  assign t[38] = t[52] ^ x[7];
  assign t[39] = t[53] ^ x[11];
  assign t[3] = ~(t[12]);
  assign t[40] = t[54] ^ x[10];
  assign t[41] = t[55] ^ x[14];
  assign t[42] = t[56] ^ x[13];
  assign t[43] = t[57] ^ x[17];
  assign t[44] = t[58] ^ x[16];
  assign t[45] = t[59] ^ x[20];
  assign t[46] = t[60] ^ x[19];
  assign t[47] = (x[0]);
  assign t[48] = (x[0]);
  assign t[49] = (x[3]);
  assign t[4] = ~(t[13]);
  assign t[50] = (x[3]);
  assign t[51] = (x[6]);
  assign t[52] = (x[6]);
  assign t[53] = (x[9]);
  assign t[54] = (x[9]);
  assign t[55] = (x[12]);
  assign t[56] = (x[12]);
  assign t[57] = (x[15]);
  assign t[58] = (x[15]);
  assign t[59] = (x[18]);
  assign t[5] = ~(t[6]);
  assign t[60] = (x[18]);
  assign t[6] = ~(t[14] | t[7]);
  assign t[7] = ~(t[8]);
  assign t[8] = ~(t[9] & t[10]);
  assign t[9] = ~(t[15]);
  assign y = (t[0]);
endmodule

module R2ind30(x, y);
 input [11:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[5] | t[1]);
  assign t[10] = t[14] ^ x[5];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[11];
  assign t[13] = (t[17] & ~t[18]);
  assign t[14] = (t[19] & ~t[20]);
  assign t[15] = (t[21] & ~t[22]);
  assign t[16] = (t[23] & ~t[24]);
  assign t[17] = t[25] ^ x[2];
  assign t[18] = t[26] ^ x[1];
  assign t[19] = t[27] ^ x[5];
  assign t[1] = ~(t[6] & t[2]);
  assign t[20] = t[28] ^ x[4];
  assign t[21] = t[29] ^ x[8];
  assign t[22] = t[30] ^ x[7];
  assign t[23] = t[31] ^ x[11];
  assign t[24] = t[32] ^ x[10];
  assign t[25] = (x[0]);
  assign t[26] = (x[0]);
  assign t[27] = (x[3]);
  assign t[28] = (x[3]);
  assign t[29] = (x[6]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = (x[6]);
  assign t[31] = (x[9]);
  assign t[32] = (x[9]);
  assign t[3] = ~(t[4]);
  assign t[4] = ~(t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind31(x, y);
 input [11:0] x;
 output y;

 wire [32:0] t;
  assign t[0] = ~(t[5] | t[1]);
  assign t[10] = t[14] ^ x[5];
  assign t[11] = t[15] ^ x[8];
  assign t[12] = t[16] ^ x[11];
  assign t[13] = (t[17] & ~t[18]);
  assign t[14] = (t[19] & ~t[20]);
  assign t[15] = (t[21] & ~t[22]);
  assign t[16] = (t[23] & ~t[24]);
  assign t[17] = t[25] ^ x[2];
  assign t[18] = t[26] ^ x[1];
  assign t[19] = t[27] ^ x[5];
  assign t[1] = ~(t[6] & t[2]);
  assign t[20] = t[28] ^ x[4];
  assign t[21] = t[29] ^ x[8];
  assign t[22] = t[30] ^ x[7];
  assign t[23] = t[31] ^ x[11];
  assign t[24] = t[32] ^ x[10];
  assign t[25] = (x[0]);
  assign t[26] = (x[0]);
  assign t[27] = (x[3]);
  assign t[28] = (x[3]);
  assign t[29] = (x[6]);
  assign t[2] = ~(t[7] | t[3]);
  assign t[30] = (x[6]);
  assign t[31] = (x[9]);
  assign t[32] = (x[9]);
  assign t[3] = ~(t[4]);
  assign t[4] = ~(t[8]);
  assign t[5] = (t[9]);
  assign t[6] = (t[10]);
  assign t[7] = (t[11]);
  assign t[8] = (t[12]);
  assign t[9] = t[13] ^ x[2];
  assign y = (t[0]);
endmodule

module R2ind32(x, y);
 input [12:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[3];
  assign t[14] = t[18] ^ x[6];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[12];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[3];
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[6];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[9];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = (x[1]);
  assign t[2] = ~(x[0]);
  assign t[30] = (x[1]);
  assign t[31] = (x[4]);
  assign t[32] = (x[4]);
  assign t[33] = (x[7]);
  assign t[34] = (x[7]);
  assign t[35] = (x[10]);
  assign t[36] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind33(x, y);
 input [12:0] x;
 output y;

 wire [36:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = t[17] ^ x[3];
  assign t[14] = t[18] ^ x[6];
  assign t[15] = t[19] ^ x[9];
  assign t[16] = t[20] ^ x[12];
  assign t[17] = (t[21] & ~t[22]);
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = ~(t[3]);
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = t[29] ^ x[3];
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[6];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[9];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[12];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = (x[1]);
  assign t[2] = ~(x[0]);
  assign t[30] = (x[1]);
  assign t[31] = (x[4]);
  assign t[32] = (x[4]);
  assign t[33] = (x[7]);
  assign t[34] = (x[7]);
  assign t[35] = (x[10]);
  assign t[36] = (x[10]);
  assign t[3] = ~(t[4] | t[5]);
  assign t[4] = ~(t[6] & t[7]);
  assign t[5] = ~(t[9] & t[8]);
  assign t[6] = ~(t[10]);
  assign t[7] = ~(t[11]);
  assign t[8] = ~(t[12]);
  assign t[9] = (t[13]);
  assign y = (t[0]);
endmodule

module R2ind34(x, y);
 input [17:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = t[20] ^ x[2];
  assign t[15] = t[21] ^ x[5];
  assign t[16] = t[22] ^ x[8];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = ~(t[8] | t[3]);
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = (t[34] & ~t[35]);
  assign t[25] = (t[36] & ~t[37]);
  assign t[26] = t[38] ^ x[2];
  assign t[27] = t[39] ^ x[1];
  assign t[28] = t[40] ^ x[5];
  assign t[29] = t[41] ^ x[4];
  assign t[2] = ~(t[9]);
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[7];
  assign t[32] = t[44] ^ x[11];
  assign t[33] = t[45] ^ x[10];
  assign t[34] = t[46] ^ x[14];
  assign t[35] = t[47] ^ x[13];
  assign t[36] = t[48] ^ x[17];
  assign t[37] = t[49] ^ x[16];
  assign t[38] = (x[0]);
  assign t[39] = (x[0]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[3]);
  assign t[41] = (x[3]);
  assign t[42] = (x[6]);
  assign t[43] = (x[6]);
  assign t[44] = (x[9]);
  assign t[45] = (x[9]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[15]);
  assign t[49] = (x[15]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = t[7] & t[11];
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind35(x, y);
 input [17:0] x;
 output y;

 wire [49:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = t[20] ^ x[2];
  assign t[15] = t[21] ^ x[5];
  assign t[16] = t[22] ^ x[8];
  assign t[17] = t[23] ^ x[11];
  assign t[18] = t[24] ^ x[14];
  assign t[19] = t[25] ^ x[17];
  assign t[1] = ~(t[8] | t[3]);
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = (t[34] & ~t[35]);
  assign t[25] = (t[36] & ~t[37]);
  assign t[26] = t[38] ^ x[2];
  assign t[27] = t[39] ^ x[1];
  assign t[28] = t[40] ^ x[5];
  assign t[29] = t[41] ^ x[4];
  assign t[2] = ~(t[9]);
  assign t[30] = t[42] ^ x[8];
  assign t[31] = t[43] ^ x[7];
  assign t[32] = t[44] ^ x[11];
  assign t[33] = t[45] ^ x[10];
  assign t[34] = t[46] ^ x[14];
  assign t[35] = t[47] ^ x[13];
  assign t[36] = t[48] ^ x[17];
  assign t[37] = t[49] ^ x[16];
  assign t[38] = (x[0]);
  assign t[39] = (x[0]);
  assign t[3] = ~(t[4]);
  assign t[40] = (x[3]);
  assign t[41] = (x[3]);
  assign t[42] = (x[6]);
  assign t[43] = (x[6]);
  assign t[44] = (x[9]);
  assign t[45] = (x[9]);
  assign t[46] = (x[12]);
  assign t[47] = (x[12]);
  assign t[48] = (x[15]);
  assign t[49] = (x[15]);
  assign t[4] = ~(t[5] & t[6]);
  assign t[5] = ~(t[10]);
  assign t[6] = t[7] & t[11];
  assign t[7] = ~(t[12] | t[13]);
  assign t[8] = (t[14]);
  assign t[9] = (t[15]);
  assign y = (t[0]);
endmodule

module R2ind36(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind37(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind38(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind39(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind40(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind41(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind42(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind43(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind44(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind45(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind46(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind47(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind48(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind49(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind50(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind51(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind52(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind53(x, y);
 input [2:0] x;
 output y;

 wire [7:0] t;
  assign t[0] = ~(t[1]);
  assign t[1] = (t[2]);
  assign t[2] = t[3] ^ x[2];
  assign t[3] = (t[4] & ~t[5]);
  assign t[4] = t[6] ^ x[2];
  assign t[5] = t[7] ^ x[1];
  assign t[6] = (x[0]);
  assign t[7] = (x[0]);
  assign y = (t[0]);
endmodule

module R2ind54(x, y);
 input [31:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[20] ^ t[21];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[22]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[14] = ~(x[28]);
  assign t[15] = ~(t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = t[16] ? t[4] : t[3];
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = t[40] ^ x[15];
  assign t[31] = t[41] ^ x[18];
  assign t[32] = t[42] ^ x[21];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = t[44] ^ x[27];
  assign t[35] = t[45] ^ x[31];
  assign t[36] = (t[46] & ~t[47]);
  assign t[37] = (t[48] & ~t[49]);
  assign t[38] = (t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[53]);
  assign t[3] = ~(t[17]);
  assign t[40] = (t[54] & ~t[55]);
  assign t[41] = (t[56] & ~t[57]);
  assign t[42] = (t[58] & ~t[59]);
  assign t[43] = (t[60] & ~t[61]);
  assign t[44] = (t[62] & ~t[63]);
  assign t[45] = (t[64] & ~t[65]);
  assign t[46] = t[66] ^ x[2];
  assign t[47] = t[67] ^ x[1];
  assign t[48] = t[68] ^ x[5];
  assign t[49] = t[69] ^ x[4];
  assign t[4] = ~(t[18] & t[7]);
  assign t[50] = t[70] ^ x[8];
  assign t[51] = t[71] ^ x[7];
  assign t[52] = t[72] ^ x[11];
  assign t[53] = t[73] ^ x[10];
  assign t[54] = t[74] ^ x[15];
  assign t[55] = t[75] ^ x[14];
  assign t[56] = t[76] ^ x[18];
  assign t[57] = t[77] ^ x[17];
  assign t[58] = t[78] ^ x[21];
  assign t[59] = t[79] ^ x[20];
  assign t[5] = ~(t[18] | t[8]);
  assign t[60] = t[80] ^ x[24];
  assign t[61] = t[81] ^ x[23];
  assign t[62] = t[82] ^ x[27];
  assign t[63] = t[83] ^ x[26];
  assign t[64] = t[84] ^ x[31];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = (x[0]);
  assign t[67] = (x[0]);
  assign t[68] = (x[3]);
  assign t[69] = (x[3]);
  assign t[6] = t[19] ? t[10] : t[9];
  assign t[70] = (x[6]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[9]);
  assign t[74] = (x[13]);
  assign t[75] = (x[13]);
  assign t[76] = (x[16]);
  assign t[77] = (x[16]);
  assign t[78] = (x[19]);
  assign t[79] = (x[19]);
  assign t[7] = t[11] ? x[12] : t[17];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[25]);
  assign t[83] = (x[25]);
  assign t[84] = (x[29]);
  assign t[85] = (x[29]);
  assign t[8] = ~(t[16]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0]);
endmodule

module R2ind55(x, y);
 input [31:0] x;
 output y;

 wire [85:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[20] ^ t[21];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[22]);
  assign t[13] = ~(t[23] ^ t[24]);
  assign t[14] = ~(x[28]);
  assign t[15] = ~(t[25]);
  assign t[16] = (t[26]);
  assign t[17] = (t[27]);
  assign t[18] = (t[28]);
  assign t[19] = (t[29]);
  assign t[1] = t[16] ? t[4] : t[3];
  assign t[20] = (t[30]);
  assign t[21] = (t[31]);
  assign t[22] = (t[32]);
  assign t[23] = (t[33]);
  assign t[24] = (t[34]);
  assign t[25] = (t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = t[40] ^ x[15];
  assign t[31] = t[41] ^ x[18];
  assign t[32] = t[42] ^ x[21];
  assign t[33] = t[43] ^ x[24];
  assign t[34] = t[44] ^ x[27];
  assign t[35] = t[45] ^ x[31];
  assign t[36] = (t[46] & ~t[47]);
  assign t[37] = (t[48] & ~t[49]);
  assign t[38] = (t[50] & ~t[51]);
  assign t[39] = (t[52] & ~t[53]);
  assign t[3] = ~(t[17]);
  assign t[40] = (t[54] & ~t[55]);
  assign t[41] = (t[56] & ~t[57]);
  assign t[42] = (t[58] & ~t[59]);
  assign t[43] = (t[60] & ~t[61]);
  assign t[44] = (t[62] & ~t[63]);
  assign t[45] = (t[64] & ~t[65]);
  assign t[46] = t[66] ^ x[2];
  assign t[47] = t[67] ^ x[1];
  assign t[48] = t[68] ^ x[5];
  assign t[49] = t[69] ^ x[4];
  assign t[4] = ~(t[18] & t[7]);
  assign t[50] = t[70] ^ x[8];
  assign t[51] = t[71] ^ x[7];
  assign t[52] = t[72] ^ x[11];
  assign t[53] = t[73] ^ x[10];
  assign t[54] = t[74] ^ x[15];
  assign t[55] = t[75] ^ x[14];
  assign t[56] = t[76] ^ x[18];
  assign t[57] = t[77] ^ x[17];
  assign t[58] = t[78] ^ x[21];
  assign t[59] = t[79] ^ x[20];
  assign t[5] = ~(t[18] | t[8]);
  assign t[60] = t[80] ^ x[24];
  assign t[61] = t[81] ^ x[23];
  assign t[62] = t[82] ^ x[27];
  assign t[63] = t[83] ^ x[26];
  assign t[64] = t[84] ^ x[31];
  assign t[65] = t[85] ^ x[30];
  assign t[66] = (x[0]);
  assign t[67] = (x[0]);
  assign t[68] = (x[3]);
  assign t[69] = (x[3]);
  assign t[6] = t[19] ? t[10] : t[9];
  assign t[70] = (x[6]);
  assign t[71] = (x[6]);
  assign t[72] = (x[9]);
  assign t[73] = (x[9]);
  assign t[74] = (x[13]);
  assign t[75] = (x[13]);
  assign t[76] = (x[16]);
  assign t[77] = (x[16]);
  assign t[78] = (x[19]);
  assign t[79] = (x[19]);
  assign t[7] = t[11] ? x[12] : t[17];
  assign t[80] = (x[22]);
  assign t[81] = (x[22]);
  assign t[82] = (x[25]);
  assign t[83] = (x[25]);
  assign t[84] = (x[29]);
  assign t[85] = (x[29]);
  assign t[8] = ~(t[16]);
  assign t[9] = ~(t[12] ^ t[13]);
  assign y = (t[0]);
endmodule

module R2ind56(x, y);
 input [34:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[28] ^ t[29];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(x[22]);
  assign t[15] = ~(t[19] | t[17]);
  assign t[16] = t[30] ? t[20] : t[31];
  assign t[17] = ~(t[32]);
  assign t[18] = ~(t[30] ^ t[33]);
  assign t[19] = ~(t[30] | t[33]);
  assign t[1] = t[23] ? t[4] : t[3];
  assign t[20] = ~(t[31] & t[21]);
  assign t[21] = ~(t[22] & t[17]);
  assign t[22] = ~(t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = t[45] ^ x[2];
  assign t[35] = t[46] ^ x[5];
  assign t[36] = t[47] ^ x[8];
  assign t[37] = t[48] ^ x[11];
  assign t[38] = t[49] ^ x[14];
  assign t[39] = t[50] ^ x[18];
  assign t[3] = ~(t[24]);
  assign t[40] = t[51] ^ x[21];
  assign t[41] = t[52] ^ x[25];
  assign t[42] = t[53] ^ x[28];
  assign t[43] = t[54] ^ x[31];
  assign t[44] = t[55] ^ x[34];
  assign t[45] = (t[56] & ~t[57]);
  assign t[46] = (t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[61]);
  assign t[48] = (t[62] & ~t[63]);
  assign t[49] = (t[64] & ~t[65]);
  assign t[4] = ~(t[25] & t[7]);
  assign t[50] = (t[66] & ~t[67]);
  assign t[51] = (t[68] & ~t[69]);
  assign t[52] = (t[70] & ~t[71]);
  assign t[53] = (t[72] & ~t[73]);
  assign t[54] = (t[74] & ~t[75]);
  assign t[55] = (t[76] & ~t[77]);
  assign t[56] = t[78] ^ x[2];
  assign t[57] = t[79] ^ x[1];
  assign t[58] = t[80] ^ x[5];
  assign t[59] = t[81] ^ x[4];
  assign t[5] = ~(t[25] | t[8]);
  assign t[60] = t[82] ^ x[8];
  assign t[61] = t[83] ^ x[7];
  assign t[62] = t[84] ^ x[11];
  assign t[63] = t[85] ^ x[10];
  assign t[64] = t[86] ^ x[14];
  assign t[65] = t[87] ^ x[13];
  assign t[66] = t[88] ^ x[18];
  assign t[67] = t[89] ^ x[17];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[20];
  assign t[6] = t[26] ? t[10] : t[9];
  assign t[70] = t[92] ^ x[25];
  assign t[71] = t[93] ^ x[24];
  assign t[72] = t[94] ^ x[28];
  assign t[73] = t[95] ^ x[27];
  assign t[74] = t[96] ^ x[31];
  assign t[75] = t[97] ^ x[30];
  assign t[76] = t[98] ^ x[34];
  assign t[77] = t[99] ^ x[33];
  assign t[78] = (x[0]);
  assign t[79] = (x[0]);
  assign t[7] = t[11] ? x[15] : t[27];
  assign t[80] = (x[3]);
  assign t[81] = (x[3]);
  assign t[82] = (x[6]);
  assign t[83] = (x[6]);
  assign t[84] = (x[9]);
  assign t[85] = (x[9]);
  assign t[86] = (x[12]);
  assign t[87] = (x[12]);
  assign t[88] = (x[16]);
  assign t[89] = (x[16]);
  assign t[8] = ~(t[23]);
  assign t[90] = (x[19]);
  assign t[91] = (x[19]);
  assign t[92] = (x[23]);
  assign t[93] = (x[23]);
  assign t[94] = (x[26]);
  assign t[95] = (x[26]);
  assign t[96] = (x[29]);
  assign t[97] = (x[29]);
  assign t[98] = (x[32]);
  assign t[99] = (x[32]);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind57(x, y);
 input [34:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[28] ^ t[29];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] | t[16]);
  assign t[13] = ~(t[17] | t[18]);
  assign t[14] = ~(x[22]);
  assign t[15] = ~(t[19] | t[17]);
  assign t[16] = t[30] ? t[20] : t[31];
  assign t[17] = ~(t[32]);
  assign t[18] = ~(t[30] ^ t[33]);
  assign t[19] = ~(t[30] | t[33]);
  assign t[1] = t[23] ? t[4] : t[3];
  assign t[20] = ~(t[31] & t[21]);
  assign t[21] = ~(t[22] & t[17]);
  assign t[22] = ~(t[33]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = t[45] ^ x[2];
  assign t[35] = t[46] ^ x[5];
  assign t[36] = t[47] ^ x[8];
  assign t[37] = t[48] ^ x[11];
  assign t[38] = t[49] ^ x[14];
  assign t[39] = t[50] ^ x[18];
  assign t[3] = ~(t[24]);
  assign t[40] = t[51] ^ x[21];
  assign t[41] = t[52] ^ x[25];
  assign t[42] = t[53] ^ x[28];
  assign t[43] = t[54] ^ x[31];
  assign t[44] = t[55] ^ x[34];
  assign t[45] = (t[56] & ~t[57]);
  assign t[46] = (t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[61]);
  assign t[48] = (t[62] & ~t[63]);
  assign t[49] = (t[64] & ~t[65]);
  assign t[4] = ~(t[25] & t[7]);
  assign t[50] = (t[66] & ~t[67]);
  assign t[51] = (t[68] & ~t[69]);
  assign t[52] = (t[70] & ~t[71]);
  assign t[53] = (t[72] & ~t[73]);
  assign t[54] = (t[74] & ~t[75]);
  assign t[55] = (t[76] & ~t[77]);
  assign t[56] = t[78] ^ x[2];
  assign t[57] = t[79] ^ x[1];
  assign t[58] = t[80] ^ x[5];
  assign t[59] = t[81] ^ x[4];
  assign t[5] = ~(t[25] | t[8]);
  assign t[60] = t[82] ^ x[8];
  assign t[61] = t[83] ^ x[7];
  assign t[62] = t[84] ^ x[11];
  assign t[63] = t[85] ^ x[10];
  assign t[64] = t[86] ^ x[14];
  assign t[65] = t[87] ^ x[13];
  assign t[66] = t[88] ^ x[18];
  assign t[67] = t[89] ^ x[17];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[20];
  assign t[6] = t[26] ? t[10] : t[9];
  assign t[70] = t[92] ^ x[25];
  assign t[71] = t[93] ^ x[24];
  assign t[72] = t[94] ^ x[28];
  assign t[73] = t[95] ^ x[27];
  assign t[74] = t[96] ^ x[31];
  assign t[75] = t[97] ^ x[30];
  assign t[76] = t[98] ^ x[34];
  assign t[77] = t[99] ^ x[33];
  assign t[78] = (x[0]);
  assign t[79] = (x[0]);
  assign t[7] = t[11] ? x[15] : t[27];
  assign t[80] = (x[3]);
  assign t[81] = (x[3]);
  assign t[82] = (x[6]);
  assign t[83] = (x[6]);
  assign t[84] = (x[9]);
  assign t[85] = (x[9]);
  assign t[86] = (x[12]);
  assign t[87] = (x[12]);
  assign t[88] = (x[16]);
  assign t[89] = (x[16]);
  assign t[8] = ~(t[23]);
  assign t[90] = (x[19]);
  assign t[91] = (x[19]);
  assign t[92] = (x[23]);
  assign t[93] = (x[23]);
  assign t[94] = (x[26]);
  assign t[95] = (x[26]);
  assign t[96] = (x[29]);
  assign t[97] = (x[29]);
  assign t[98] = (x[32]);
  assign t[99] = (x[32]);
  assign t[9] = ~(t[12] | t[13]);
  assign y = (t[0]);
endmodule

module R2ind58(x, y);
 input [34:0] x;
 output y;

 wire [103:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[29]);
  assign t[101] = (x[29]);
  assign t[102] = (x[32]);
  assign t[103] = (x[32]);
  assign t[10] = t[32] ^ t[33];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(x[22]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[35] & t[20]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = t[36] ? t[16] : t[35];
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = t[27] ? t[4] : t[3];
  assign t[20] = ~(t[25] & t[22]);
  assign t[21] = ~(t[36] | t[37]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[36]);
  assign t[24] = ~(t[25] & t[26]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[35]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = (t[45]);
  assign t[35] = (t[46]);
  assign t[36] = (t[47]);
  assign t[37] = (t[48]);
  assign t[38] = t[49] ^ x[2];
  assign t[39] = t[50] ^ x[5];
  assign t[3] = ~(t[28]);
  assign t[40] = t[51] ^ x[8];
  assign t[41] = t[52] ^ x[11];
  assign t[42] = t[53] ^ x[14];
  assign t[43] = t[54] ^ x[18];
  assign t[44] = t[55] ^ x[21];
  assign t[45] = t[56] ^ x[25];
  assign t[46] = t[57] ^ x[28];
  assign t[47] = t[58] ^ x[31];
  assign t[48] = t[59] ^ x[34];
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = ~(t[29] & t[7]);
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = (t[78] & ~t[79]);
  assign t[59] = (t[80] & ~t[81]);
  assign t[5] = ~(t[29] | t[8]);
  assign t[60] = t[82] ^ x[2];
  assign t[61] = t[83] ^ x[1];
  assign t[62] = t[84] ^ x[5];
  assign t[63] = t[85] ^ x[4];
  assign t[64] = t[86] ^ x[8];
  assign t[65] = t[87] ^ x[7];
  assign t[66] = t[88] ^ x[11];
  assign t[67] = t[89] ^ x[10];
  assign t[68] = t[90] ^ x[14];
  assign t[69] = t[91] ^ x[13];
  assign t[6] = t[30] ? t[10] : t[9];
  assign t[70] = t[92] ^ x[18];
  assign t[71] = t[93] ^ x[17];
  assign t[72] = t[94] ^ x[21];
  assign t[73] = t[95] ^ x[20];
  assign t[74] = t[96] ^ x[25];
  assign t[75] = t[97] ^ x[24];
  assign t[76] = t[98] ^ x[28];
  assign t[77] = t[99] ^ x[27];
  assign t[78] = t[100] ^ x[31];
  assign t[79] = t[101] ^ x[30];
  assign t[7] = t[11] ? x[15] : t[31];
  assign t[80] = t[102] ^ x[34];
  assign t[81] = t[103] ^ x[33];
  assign t[82] = (x[0]);
  assign t[83] = (x[0]);
  assign t[84] = (x[3]);
  assign t[85] = (x[3]);
  assign t[86] = (x[6]);
  assign t[87] = (x[6]);
  assign t[88] = (x[9]);
  assign t[89] = (x[9]);
  assign t[8] = ~(t[27]);
  assign t[90] = (x[12]);
  assign t[91] = (x[12]);
  assign t[92] = (x[16]);
  assign t[93] = (x[16]);
  assign t[94] = (x[19]);
  assign t[95] = (x[19]);
  assign t[96] = (x[23]);
  assign t[97] = (x[23]);
  assign t[98] = (x[26]);
  assign t[99] = (x[26]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind59(x, y);
 input [34:0] x;
 output y;

 wire [103:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[100] = (x[29]);
  assign t[101] = (x[29]);
  assign t[102] = (x[32]);
  assign t[103] = (x[32]);
  assign t[10] = t[32] ^ t[33];
  assign t[11] = ~(t[14]);
  assign t[12] = ~(t[15] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(x[22]);
  assign t[15] = ~(t[34] | t[19]);
  assign t[16] = ~(t[35] & t[20]);
  assign t[17] = ~(t[21] | t[22]);
  assign t[18] = t[36] ? t[16] : t[35];
  assign t[19] = ~(t[23] | t[24]);
  assign t[1] = t[27] ? t[4] : t[3];
  assign t[20] = ~(t[25] & t[22]);
  assign t[21] = ~(t[36] | t[37]);
  assign t[22] = ~(t[34]);
  assign t[23] = ~(t[36]);
  assign t[24] = ~(t[25] & t[26]);
  assign t[25] = ~(t[37]);
  assign t[26] = ~(t[35]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = (t[45]);
  assign t[35] = (t[46]);
  assign t[36] = (t[47]);
  assign t[37] = (t[48]);
  assign t[38] = t[49] ^ x[2];
  assign t[39] = t[50] ^ x[5];
  assign t[3] = ~(t[28]);
  assign t[40] = t[51] ^ x[8];
  assign t[41] = t[52] ^ x[11];
  assign t[42] = t[53] ^ x[14];
  assign t[43] = t[54] ^ x[18];
  assign t[44] = t[55] ^ x[21];
  assign t[45] = t[56] ^ x[25];
  assign t[46] = t[57] ^ x[28];
  assign t[47] = t[58] ^ x[31];
  assign t[48] = t[59] ^ x[34];
  assign t[49] = (t[60] & ~t[61]);
  assign t[4] = ~(t[29] & t[7]);
  assign t[50] = (t[62] & ~t[63]);
  assign t[51] = (t[64] & ~t[65]);
  assign t[52] = (t[66] & ~t[67]);
  assign t[53] = (t[68] & ~t[69]);
  assign t[54] = (t[70] & ~t[71]);
  assign t[55] = (t[72] & ~t[73]);
  assign t[56] = (t[74] & ~t[75]);
  assign t[57] = (t[76] & ~t[77]);
  assign t[58] = (t[78] & ~t[79]);
  assign t[59] = (t[80] & ~t[81]);
  assign t[5] = ~(t[29] | t[8]);
  assign t[60] = t[82] ^ x[2];
  assign t[61] = t[83] ^ x[1];
  assign t[62] = t[84] ^ x[5];
  assign t[63] = t[85] ^ x[4];
  assign t[64] = t[86] ^ x[8];
  assign t[65] = t[87] ^ x[7];
  assign t[66] = t[88] ^ x[11];
  assign t[67] = t[89] ^ x[10];
  assign t[68] = t[90] ^ x[14];
  assign t[69] = t[91] ^ x[13];
  assign t[6] = t[30] ? t[10] : t[9];
  assign t[70] = t[92] ^ x[18];
  assign t[71] = t[93] ^ x[17];
  assign t[72] = t[94] ^ x[21];
  assign t[73] = t[95] ^ x[20];
  assign t[74] = t[96] ^ x[25];
  assign t[75] = t[97] ^ x[24];
  assign t[76] = t[98] ^ x[28];
  assign t[77] = t[99] ^ x[27];
  assign t[78] = t[100] ^ x[31];
  assign t[79] = t[101] ^ x[30];
  assign t[7] = t[11] ? x[15] : t[31];
  assign t[80] = t[102] ^ x[34];
  assign t[81] = t[103] ^ x[33];
  assign t[82] = (x[0]);
  assign t[83] = (x[0]);
  assign t[84] = (x[3]);
  assign t[85] = (x[3]);
  assign t[86] = (x[6]);
  assign t[87] = (x[6]);
  assign t[88] = (x[9]);
  assign t[89] = (x[9]);
  assign t[8] = ~(t[27]);
  assign t[90] = (x[12]);
  assign t[91] = (x[12]);
  assign t[92] = (x[16]);
  assign t[93] = (x[16]);
  assign t[94] = (x[19]);
  assign t[95] = (x[19]);
  assign t[96] = (x[23]);
  assign t[97] = (x[23]);
  assign t[98] = (x[26]);
  assign t[99] = (x[26]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind60(x, y);
 input [34:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[28] ^ t[29];
  assign t[11] = ~(t[14]);
  assign t[12] = t[30] ? t[16] : t[15];
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(x[25]);
  assign t[15] = ~(t[31] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[30] | t[32]);
  assign t[18] = ~(t[31]);
  assign t[19] = ~(t[22] & t[20]);
  assign t[1] = t[23] ? t[4] : t[3];
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[22] & t[18]);
  assign t[22] = ~(t[32]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = t[45] ^ x[2];
  assign t[35] = t[46] ^ x[5];
  assign t[36] = t[47] ^ x[8];
  assign t[37] = t[48] ^ x[11];
  assign t[38] = t[49] ^ x[14];
  assign t[39] = t[50] ^ x[18];
  assign t[3] = ~(t[24]);
  assign t[40] = t[51] ^ x[21];
  assign t[41] = t[52] ^ x[24];
  assign t[42] = t[53] ^ x[28];
  assign t[43] = t[54] ^ x[31];
  assign t[44] = t[55] ^ x[34];
  assign t[45] = (t[56] & ~t[57]);
  assign t[46] = (t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[61]);
  assign t[48] = (t[62] & ~t[63]);
  assign t[49] = (t[64] & ~t[65]);
  assign t[4] = ~(t[25] & t[7]);
  assign t[50] = (t[66] & ~t[67]);
  assign t[51] = (t[68] & ~t[69]);
  assign t[52] = (t[70] & ~t[71]);
  assign t[53] = (t[72] & ~t[73]);
  assign t[54] = (t[74] & ~t[75]);
  assign t[55] = (t[76] & ~t[77]);
  assign t[56] = t[78] ^ x[2];
  assign t[57] = t[79] ^ x[1];
  assign t[58] = t[80] ^ x[5];
  assign t[59] = t[81] ^ x[4];
  assign t[5] = ~(t[25] | t[8]);
  assign t[60] = t[82] ^ x[8];
  assign t[61] = t[83] ^ x[7];
  assign t[62] = t[84] ^ x[11];
  assign t[63] = t[85] ^ x[10];
  assign t[64] = t[86] ^ x[14];
  assign t[65] = t[87] ^ x[13];
  assign t[66] = t[88] ^ x[18];
  assign t[67] = t[89] ^ x[17];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[20];
  assign t[6] = t[26] ? t[10] : t[9];
  assign t[70] = t[92] ^ x[24];
  assign t[71] = t[93] ^ x[23];
  assign t[72] = t[94] ^ x[28];
  assign t[73] = t[95] ^ x[27];
  assign t[74] = t[96] ^ x[31];
  assign t[75] = t[97] ^ x[30];
  assign t[76] = t[98] ^ x[34];
  assign t[77] = t[99] ^ x[33];
  assign t[78] = (x[0]);
  assign t[79] = (x[0]);
  assign t[7] = t[11] ? x[15] : t[27];
  assign t[80] = (x[3]);
  assign t[81] = (x[3]);
  assign t[82] = (x[6]);
  assign t[83] = (x[6]);
  assign t[84] = (x[9]);
  assign t[85] = (x[9]);
  assign t[86] = (x[12]);
  assign t[87] = (x[12]);
  assign t[88] = (x[16]);
  assign t[89] = (x[16]);
  assign t[8] = ~(t[23]);
  assign t[90] = (x[19]);
  assign t[91] = (x[19]);
  assign t[92] = (x[22]);
  assign t[93] = (x[22]);
  assign t[94] = (x[26]);
  assign t[95] = (x[26]);
  assign t[96] = (x[29]);
  assign t[97] = (x[29]);
  assign t[98] = (x[32]);
  assign t[99] = (x[32]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind61(x, y);
 input [34:0] x;
 output y;

 wire [99:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[28] ^ t[29];
  assign t[11] = ~(t[14]);
  assign t[12] = t[30] ? t[16] : t[15];
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(x[25]);
  assign t[15] = ~(t[31] & t[19]);
  assign t[16] = ~(t[20] & t[21]);
  assign t[17] = ~(t[30] | t[32]);
  assign t[18] = ~(t[31]);
  assign t[19] = ~(t[22] & t[20]);
  assign t[1] = t[23] ? t[4] : t[3];
  assign t[20] = ~(t[33]);
  assign t[21] = ~(t[22] & t[18]);
  assign t[22] = ~(t[32]);
  assign t[23] = (t[34]);
  assign t[24] = (t[35]);
  assign t[25] = (t[36]);
  assign t[26] = (t[37]);
  assign t[27] = (t[38]);
  assign t[28] = (t[39]);
  assign t[29] = (t[40]);
  assign t[2] = ~(t[5] & t[6]);
  assign t[30] = (t[41]);
  assign t[31] = (t[42]);
  assign t[32] = (t[43]);
  assign t[33] = (t[44]);
  assign t[34] = t[45] ^ x[2];
  assign t[35] = t[46] ^ x[5];
  assign t[36] = t[47] ^ x[8];
  assign t[37] = t[48] ^ x[11];
  assign t[38] = t[49] ^ x[14];
  assign t[39] = t[50] ^ x[18];
  assign t[3] = ~(t[24]);
  assign t[40] = t[51] ^ x[21];
  assign t[41] = t[52] ^ x[24];
  assign t[42] = t[53] ^ x[28];
  assign t[43] = t[54] ^ x[31];
  assign t[44] = t[55] ^ x[34];
  assign t[45] = (t[56] & ~t[57]);
  assign t[46] = (t[58] & ~t[59]);
  assign t[47] = (t[60] & ~t[61]);
  assign t[48] = (t[62] & ~t[63]);
  assign t[49] = (t[64] & ~t[65]);
  assign t[4] = ~(t[25] & t[7]);
  assign t[50] = (t[66] & ~t[67]);
  assign t[51] = (t[68] & ~t[69]);
  assign t[52] = (t[70] & ~t[71]);
  assign t[53] = (t[72] & ~t[73]);
  assign t[54] = (t[74] & ~t[75]);
  assign t[55] = (t[76] & ~t[77]);
  assign t[56] = t[78] ^ x[2];
  assign t[57] = t[79] ^ x[1];
  assign t[58] = t[80] ^ x[5];
  assign t[59] = t[81] ^ x[4];
  assign t[5] = ~(t[25] | t[8]);
  assign t[60] = t[82] ^ x[8];
  assign t[61] = t[83] ^ x[7];
  assign t[62] = t[84] ^ x[11];
  assign t[63] = t[85] ^ x[10];
  assign t[64] = t[86] ^ x[14];
  assign t[65] = t[87] ^ x[13];
  assign t[66] = t[88] ^ x[18];
  assign t[67] = t[89] ^ x[17];
  assign t[68] = t[90] ^ x[21];
  assign t[69] = t[91] ^ x[20];
  assign t[6] = t[26] ? t[10] : t[9];
  assign t[70] = t[92] ^ x[24];
  assign t[71] = t[93] ^ x[23];
  assign t[72] = t[94] ^ x[28];
  assign t[73] = t[95] ^ x[27];
  assign t[74] = t[96] ^ x[31];
  assign t[75] = t[97] ^ x[30];
  assign t[76] = t[98] ^ x[34];
  assign t[77] = t[99] ^ x[33];
  assign t[78] = (x[0]);
  assign t[79] = (x[0]);
  assign t[7] = t[11] ? x[15] : t[27];
  assign t[80] = (x[3]);
  assign t[81] = (x[3]);
  assign t[82] = (x[6]);
  assign t[83] = (x[6]);
  assign t[84] = (x[9]);
  assign t[85] = (x[9]);
  assign t[86] = (x[12]);
  assign t[87] = (x[12]);
  assign t[88] = (x[16]);
  assign t[89] = (x[16]);
  assign t[8] = ~(t[23]);
  assign t[90] = (x[19]);
  assign t[91] = (x[19]);
  assign t[92] = (x[22]);
  assign t[93] = (x[22]);
  assign t[94] = (x[26]);
  assign t[95] = (x[26]);
  assign t[96] = (x[29]);
  assign t[97] = (x[29]);
  assign t[98] = (x[32]);
  assign t[99] = (x[32]);
  assign t[9] = ~(t[12] & t[13]);
  assign y = (t[0]);
endmodule

module R2ind62(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind63(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind64(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind65(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind66(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind67(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind68(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind69(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind70(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind71(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind72(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind73(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind74(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind75(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind76(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind77(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind78(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind79(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind80(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind81(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind82(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind83(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind84(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind85(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind86(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind87(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind88(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind89(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind90(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind91(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind92(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind93(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind94(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind95(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind96(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind97(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind98(x, y);
 input [13:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = t[22] ^ x[11];
  assign t[19] = (t[23] & ~t[24]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[1];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[4];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[7];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[38] ^ x[10];
  assign t[31] = (x[0]);
  assign t[32] = (x[0]);
  assign t[33] = (x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6]);
  assign t[36] = (x[6]);
  assign t[37] = (x[9]);
  assign t[38] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[12] : t[12];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind99(x, y);
 input [13:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = t[22] ^ x[11];
  assign t[19] = (t[23] & ~t[24]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[1];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[4];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[7];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[38] ^ x[10];
  assign t[31] = (x[0]);
  assign t[32] = (x[0]);
  assign t[33] = (x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6]);
  assign t[36] = (x[6]);
  assign t[37] = (x[9]);
  assign t[38] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[12] : t[12];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind100(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind101(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind102(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind103(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind104(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind105(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind106(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind107(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind108(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind109(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind110(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind111(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind112(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind113(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind114(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind115(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind116(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind117(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind118(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind119(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind120(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind121(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind122(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind123(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind124(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind125(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind126(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind127(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind128(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind129(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind130(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind131(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind132(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind133(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind134(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind135(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind136(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind137(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind138(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind139(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind140(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind141(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind142(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind143(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind144(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind145(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind146(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind147(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind148(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind149(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind150(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind151(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind152(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind153(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind154(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind155(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind156(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind157(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind158(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind159(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind160(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind161(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind162(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind163(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind164(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind165(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind166(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind167(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind168(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind169(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind170(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind171(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind172(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind173(x, y);
 input [19:0] x;
 output y;

 wire [51:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[16]);
  assign t[11] = (t[17]);
  assign t[12] = (t[18]);
  assign t[13] = (t[19]);
  assign t[14] = (t[20]);
  assign t[15] = (t[21]);
  assign t[16] = t[22] ^ x[2];
  assign t[17] = t[23] ^ x[5];
  assign t[18] = t[24] ^ x[8];
  assign t[19] = t[25] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[26] ^ x[16];
  assign t[21] = t[27] ^ x[19];
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = (t[36] & ~t[37]);
  assign t[27] = (t[38] & ~t[39]);
  assign t[28] = t[40] ^ x[2];
  assign t[29] = t[41] ^ x[1];
  assign t[2] = ~(t[6] & t[10]);
  assign t[30] = t[42] ^ x[5];
  assign t[31] = t[43] ^ x[4];
  assign t[32] = t[44] ^ x[8];
  assign t[33] = t[45] ^ x[7];
  assign t[34] = t[46] ^ x[11];
  assign t[35] = t[47] ^ x[10];
  assign t[36] = t[48] ^ x[16];
  assign t[37] = t[49] ^ x[15];
  assign t[38] = t[50] ^ x[19];
  assign t[39] = t[51] ^ x[18];
  assign t[3] = ~(t[7]);
  assign t[40] = (x[0]);
  assign t[41] = (x[0]);
  assign t[42] = (x[3]);
  assign t[43] = (x[3]);
  assign t[44] = (x[6]);
  assign t[45] = (x[6]);
  assign t[46] = (x[9]);
  assign t[47] = (x[9]);
  assign t[48] = (x[14]);
  assign t[49] = (x[14]);
  assign t[4] = ~(t[11]);
  assign t[50] = (x[17]);
  assign t[51] = (x[17]);
  assign t[5] = ~(t[12] & t[8]);
  assign t[6] = ~(t[12] | t[7]);
  assign t[7] = ~(t[13]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = t[14] ^ t[15];
  assign y = (t[0]);
endmodule

module R2ind174(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind175(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind176(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind177(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind178(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind179(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind180(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind181(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind182(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind183(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind184(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind185(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind186(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind187(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind188(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind189(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind190(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind191(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind192(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind193(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind194(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind195(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind196(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind197(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind198(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind199(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind200(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind201(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind202(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind203(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind204(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind205(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind206(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind207(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind208(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind209(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind210(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind211(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind212(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind213(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind214(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind215(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind216(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[2];
  assign t[15] = t[19] ^ x[5];
  assign t[16] = t[20] ^ x[8];
  assign t[17] = t[21] ^ x[11];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[1];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[4];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[7];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = (x[0]);
  assign t[31] = (x[0]);
  assign t[32] = (x[3]);
  assign t[33] = (x[3]);
  assign t[34] = (x[6]);
  assign t[35] = (x[6]);
  assign t[36] = (x[9]);
  assign t[37] = (x[9]);
  assign t[3] = ~(t[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[12] : t[12];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[13]);
  assign y = (t[0]);
endmodule

module R2ind217(x, y);
 input [13:0] x;
 output y;

 wire [37:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[14]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = t[18] ^ x[2];
  assign t[15] = t[19] ^ x[5];
  assign t[16] = t[20] ^ x[8];
  assign t[17] = t[21] ^ x[11];
  assign t[18] = (t[22] & ~t[23]);
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = t[30] ^ x[2];
  assign t[23] = t[31] ^ x[1];
  assign t[24] = t[32] ^ x[5];
  assign t[25] = t[33] ^ x[4];
  assign t[26] = t[34] ^ x[8];
  assign t[27] = t[35] ^ x[7];
  assign t[28] = t[36] ^ x[11];
  assign t[29] = t[37] ^ x[10];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = (x[0]);
  assign t[31] = (x[0]);
  assign t[32] = (x[3]);
  assign t[33] = (x[3]);
  assign t[34] = (x[6]);
  assign t[35] = (x[6]);
  assign t[36] = (x[9]);
  assign t[37] = (x[9]);
  assign t[3] = ~(t[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[12] : t[12];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[13]);
  assign y = (t[0]);
endmodule

module R2ind218(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind219(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind220(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind221(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind222(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind223(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind224(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind225(x, y);
 input [16:0] x;
 output y;

 wire [44:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = t[20] ^ x[2];
  assign t[16] = t[21] ^ x[5];
  assign t[17] = t[22] ^ x[8];
  assign t[18] = t[23] ^ x[11];
  assign t[19] = t[24] ^ x[14];
  assign t[1] = t[10] ? t[4] : t[3];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = t[35] ^ x[2];
  assign t[26] = t[36] ^ x[1];
  assign t[27] = t[37] ^ x[5];
  assign t[28] = t[38] ^ x[4];
  assign t[29] = t[39] ^ x[8];
  assign t[2] = ~(t[5] & t[11]);
  assign t[30] = t[40] ^ x[7];
  assign t[31] = t[41] ^ x[11];
  assign t[32] = t[42] ^ x[10];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = t[44] ^ x[13];
  assign t[35] = (x[0]);
  assign t[36] = (x[0]);
  assign t[37] = (x[3]);
  assign t[38] = (x[3]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[12]);
  assign t[40] = (x[6]);
  assign t[41] = (x[9]);
  assign t[42] = (x[9]);
  assign t[43] = (x[12]);
  assign t[44] = (x[12]);
  assign t[4] = ~(t[13] & t[6]);
  assign t[5] = ~(t[13] | t[7]);
  assign t[6] = t[8] ? x[15] : t[14];
  assign t[7] = ~(t[10]);
  assign t[8] = ~(t[9]);
  assign t[9] = ~(x[16]);
  assign y = (t[0]);
endmodule

module R2ind226(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind227(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind228(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind229(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind230(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind231(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind232(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind233(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind234(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind235(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind236(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind237(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind238(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind239(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind240(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind241(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind242(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind243(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind244(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind245(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind246(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind247(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind248(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind249(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind250(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind251(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind252(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind253(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind254(x, y);
 input [13:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = t[22] ^ x[11];
  assign t[19] = (t[23] & ~t[24]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[1];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[4];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[7];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[38] ^ x[10];
  assign t[31] = (x[0]);
  assign t[32] = (x[0]);
  assign t[33] = (x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6]);
  assign t[36] = (x[6]);
  assign t[37] = (x[9]);
  assign t[38] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[12] : t[12];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind255(x, y);
 input [13:0] x;
 output y;

 wire [38:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[13]);
  assign t[11] = (t[15]);
  assign t[12] = (t[16]);
  assign t[13] = (t[17]);
  assign t[14] = (t[18]);
  assign t[15] = t[19] ^ x[2];
  assign t[16] = t[20] ^ x[5];
  assign t[17] = t[21] ^ x[8];
  assign t[18] = t[22] ^ x[11];
  assign t[19] = (t[23] & ~t[24]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[25] & ~t[26]);
  assign t[21] = (t[27] & ~t[28]);
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = t[31] ^ x[2];
  assign t[24] = t[32] ^ x[1];
  assign t[25] = t[33] ^ x[5];
  assign t[26] = t[34] ^ x[4];
  assign t[27] = t[35] ^ x[8];
  assign t[28] = t[36] ^ x[7];
  assign t[29] = t[37] ^ x[11];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[38] ^ x[10];
  assign t[31] = (x[0]);
  assign t[32] = (x[0]);
  assign t[33] = (x[3]);
  assign t[34] = (x[3]);
  assign t[35] = (x[6]);
  assign t[36] = (x[6]);
  assign t[37] = (x[9]);
  assign t[38] = (x[9]);
  assign t[3] = ~(t[7]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[12] : t[12];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind256(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind257(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind258(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind259(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind260(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind261(x, y);
 input [16:0] x;
 output y;

 wire [45:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(x[16]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = (t[19]);
  assign t[15] = (t[20]);
  assign t[16] = t[21] ^ x[2];
  assign t[17] = t[22] ^ x[5];
  assign t[18] = t[23] ^ x[8];
  assign t[19] = t[24] ^ x[11];
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = t[25] ^ x[14];
  assign t[21] = (t[26] & ~t[27]);
  assign t[22] = (t[28] & ~t[29]);
  assign t[23] = (t[30] & ~t[31]);
  assign t[24] = (t[32] & ~t[33]);
  assign t[25] = (t[34] & ~t[35]);
  assign t[26] = t[36] ^ x[2];
  assign t[27] = t[37] ^ x[1];
  assign t[28] = t[38] ^ x[5];
  assign t[29] = t[39] ^ x[4];
  assign t[2] = ~(t[6] & t[11]);
  assign t[30] = t[40] ^ x[8];
  assign t[31] = t[41] ^ x[7];
  assign t[32] = t[42] ^ x[11];
  assign t[33] = t[43] ^ x[10];
  assign t[34] = t[44] ^ x[14];
  assign t[35] = t[45] ^ x[13];
  assign t[36] = (x[0]);
  assign t[37] = (x[0]);
  assign t[38] = (x[3]);
  assign t[39] = (x[3]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[6]);
  assign t[41] = (x[6]);
  assign t[42] = (x[9]);
  assign t[43] = (x[9]);
  assign t[44] = (x[12]);
  assign t[45] = (x[12]);
  assign t[4] = ~(t[12]);
  assign t[5] = ~(t[13] & t[8]);
  assign t[6] = ~(t[13] | t[7]);
  assign t[7] = ~(t[14]);
  assign t[8] = t[9] ? x[15] : t[15];
  assign t[9] = ~(t[10]);
  assign y = (t[0]);
endmodule

module R2ind262(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind263(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind264(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind265(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind266(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind267(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind268(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind269(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind270(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind271(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind272(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind273(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind274(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind275(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind276(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind277(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind278(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind279(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind280(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind281(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind282(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind283(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind284(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind285(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind286(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind287(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind288(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind289(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind290(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind291(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind292(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind293(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind294(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind295(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind296(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind297(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind298(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind299(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind300(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind301(x, y);
 input [16:0] x;
 output y;

 wire [42:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = t[18] ^ x[2];
  assign t[14] = t[19] ^ x[5];
  assign t[15] = t[20] ^ x[8];
  assign t[16] = t[21] ^ x[11];
  assign t[17] = t[22] ^ x[15];
  assign t[18] = (t[23] & ~t[24]);
  assign t[19] = (t[25] & ~t[26]);
  assign t[1] = t[8] ? t[4] : t[3];
  assign t[20] = (t[27] & ~t[28]);
  assign t[21] = (t[29] & ~t[30]);
  assign t[22] = (t[31] & ~t[32]);
  assign t[23] = t[33] ^ x[2];
  assign t[24] = t[34] ^ x[1];
  assign t[25] = t[35] ^ x[5];
  assign t[26] = t[36] ^ x[4];
  assign t[27] = t[37] ^ x[8];
  assign t[28] = t[38] ^ x[7];
  assign t[29] = t[39] ^ x[11];
  assign t[2] = ~(t[5] & t[9]);
  assign t[30] = t[40] ^ x[10];
  assign t[31] = t[41] ^ x[15];
  assign t[32] = t[42] ^ x[14];
  assign t[33] = (x[0]);
  assign t[34] = (x[0]);
  assign t[35] = (x[3]);
  assign t[36] = (x[3]);
  assign t[37] = (x[6]);
  assign t[38] = (x[6]);
  assign t[39] = (x[9]);
  assign t[3] = ~(t[10]);
  assign t[40] = (x[9]);
  assign t[41] = (x[13]);
  assign t[42] = (x[13]);
  assign t[4] = ~(t[11] & t[6]);
  assign t[5] = ~(t[11] | t[7]);
  assign t[6] = x[12] ? x[16] : t[12];
  assign t[7] = ~(t[8]);
  assign t[8] = (t[13]);
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind302(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind303(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind304(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind305(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind306(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind307(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind308(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind309(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind310(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind311(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind312(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind313(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind314(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind315(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind316(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind317(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind318(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind319(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind320(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind321(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind322(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind323(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind324(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind325(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind326(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind327(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind328(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind329(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind330(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind331(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind332(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind333(x, y);
 input [16:0] x;
 output y;

 wire [43:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = (t[15]);
  assign t[11] = (t[16]);
  assign t[12] = (t[17]);
  assign t[13] = (t[18]);
  assign t[14] = t[19] ^ x[2];
  assign t[15] = t[20] ^ x[5];
  assign t[16] = t[21] ^ x[8];
  assign t[17] = t[22] ^ x[11];
  assign t[18] = t[23] ^ x[15];
  assign t[19] = (t[24] & ~t[25]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[26] & ~t[27]);
  assign t[21] = (t[28] & ~t[29]);
  assign t[22] = (t[30] & ~t[31]);
  assign t[23] = (t[32] & ~t[33]);
  assign t[24] = t[34] ^ x[2];
  assign t[25] = t[35] ^ x[1];
  assign t[26] = t[36] ^ x[5];
  assign t[27] = t[37] ^ x[4];
  assign t[28] = t[38] ^ x[8];
  assign t[29] = t[39] ^ x[7];
  assign t[2] = ~(t[6] & t[9]);
  assign t[30] = t[40] ^ x[11];
  assign t[31] = t[41] ^ x[10];
  assign t[32] = t[42] ^ x[15];
  assign t[33] = t[43] ^ x[14];
  assign t[34] = (x[0]);
  assign t[35] = (x[0]);
  assign t[36] = (x[3]);
  assign t[37] = (x[3]);
  assign t[38] = (x[6]);
  assign t[39] = (x[6]);
  assign t[3] = ~(t[7]);
  assign t[40] = (x[9]);
  assign t[41] = (x[9]);
  assign t[42] = (x[13]);
  assign t[43] = (x[13]);
  assign t[4] = ~(t[10]);
  assign t[5] = ~(t[11] & t[8]);
  assign t[6] = ~(t[11] | t[7]);
  assign t[7] = ~(t[12]);
  assign t[8] = x[12] ? x[16] : t[13];
  assign t[9] = (t[14]);
  assign y = (t[0]);
endmodule

module R2ind334(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[24] ? t[13] : t[12];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[25] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[24] | t[26]);
  assign t[15] = ~(t[25]);
  assign t[16] = ~(t[19] & t[17]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[19] & t[15]);
  assign t[19] = ~(t[26]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = t[36] ^ x[2];
  assign t[29] = t[37] ^ x[5];
  assign t[2] = ~(t[6] & t[20]);
  assign t[30] = t[38] ^ x[8];
  assign t[31] = t[39] ^ x[11];
  assign t[32] = t[40] ^ x[16];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[45]);
  assign t[37] = (t[46] & ~t[47]);
  assign t[38] = (t[48] & ~t[49]);
  assign t[39] = (t[50] & ~t[51]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[1];
  assign t[46] = t[62] ^ x[5];
  assign t[47] = t[63] ^ x[4];
  assign t[48] = t[64] ^ x[8];
  assign t[49] = t[65] ^ x[7];
  assign t[4] = ~(t[21]);
  assign t[50] = t[66] ^ x[11];
  assign t[51] = t[67] ^ x[10];
  assign t[52] = t[68] ^ x[16];
  assign t[53] = t[69] ^ x[15];
  assign t[54] = t[70] ^ x[19];
  assign t[55] = t[71] ^ x[18];
  assign t[56] = t[72] ^ x[22];
  assign t[57] = t[73] ^ x[21];
  assign t[58] = t[74] ^ x[25];
  assign t[59] = t[75] ^ x[24];
  assign t[5] = ~(t[22] & t[8]);
  assign t[60] = (x[0]);
  assign t[61] = (x[0]);
  assign t[62] = (x[3]);
  assign t[63] = (x[3]);
  assign t[64] = (x[6]);
  assign t[65] = (x[6]);
  assign t[66] = (x[9]);
  assign t[67] = (x[9]);
  assign t[68] = (x[14]);
  assign t[69] = (x[14]);
  assign t[6] = ~(t[22] | t[7]);
  assign t[70] = (x[17]);
  assign t[71] = (x[17]);
  assign t[72] = (x[20]);
  assign t[73] = (x[20]);
  assign t[74] = (x[23]);
  assign t[75] = (x[23]);
  assign t[7] = ~(t[23]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind335(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = t[24] ? t[13] : t[12];
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[25] & t[16]);
  assign t[13] = ~(t[17] & t[18]);
  assign t[14] = ~(t[24] | t[26]);
  assign t[15] = ~(t[25]);
  assign t[16] = ~(t[19] & t[17]);
  assign t[17] = ~(t[27]);
  assign t[18] = ~(t[19] & t[15]);
  assign t[19] = ~(t[26]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = t[36] ^ x[2];
  assign t[29] = t[37] ^ x[5];
  assign t[2] = ~(t[6] & t[20]);
  assign t[30] = t[38] ^ x[8];
  assign t[31] = t[39] ^ x[11];
  assign t[32] = t[40] ^ x[16];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[45]);
  assign t[37] = (t[46] & ~t[47]);
  assign t[38] = (t[48] & ~t[49]);
  assign t[39] = (t[50] & ~t[51]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[1];
  assign t[46] = t[62] ^ x[5];
  assign t[47] = t[63] ^ x[4];
  assign t[48] = t[64] ^ x[8];
  assign t[49] = t[65] ^ x[7];
  assign t[4] = ~(t[21]);
  assign t[50] = t[66] ^ x[11];
  assign t[51] = t[67] ^ x[10];
  assign t[52] = t[68] ^ x[16];
  assign t[53] = t[69] ^ x[15];
  assign t[54] = t[70] ^ x[19];
  assign t[55] = t[71] ^ x[18];
  assign t[56] = t[72] ^ x[22];
  assign t[57] = t[73] ^ x[21];
  assign t[58] = t[74] ^ x[25];
  assign t[59] = t[75] ^ x[24];
  assign t[5] = ~(t[22] & t[8]);
  assign t[60] = (x[0]);
  assign t[61] = (x[0]);
  assign t[62] = (x[3]);
  assign t[63] = (x[3]);
  assign t[64] = (x[6]);
  assign t[65] = (x[6]);
  assign t[66] = (x[9]);
  assign t[67] = (x[9]);
  assign t[68] = (x[14]);
  assign t[69] = (x[14]);
  assign t[6] = ~(t[22] | t[7]);
  assign t[70] = (x[17]);
  assign t[71] = (x[17]);
  assign t[72] = (x[20]);
  assign t[73] = (x[20]);
  assign t[74] = (x[23]);
  assign t[75] = (x[23]);
  assign t[7] = ~(t[23]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind336(x, y);
 input [25:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[28] | t[16]);
  assign t[13] = ~(t[29] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = t[30] ? t[13] : t[29];
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[22] & t[19]);
  assign t[18] = ~(t[30] | t[31]);
  assign t[19] = ~(t[28]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[29]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[6] & t[24]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[5];
  assign t[34] = t[42] ^ x[8];
  assign t[35] = t[43] ^ x[11];
  assign t[36] = t[44] ^ x[16];
  assign t[37] = t[45] ^ x[19];
  assign t[38] = t[46] ^ x[22];
  assign t[39] = t[47] ^ x[25];
  assign t[3] = ~(t[7]);
  assign t[40] = (t[48] & ~t[49]);
  assign t[41] = (t[50] & ~t[51]);
  assign t[42] = (t[52] & ~t[53]);
  assign t[43] = (t[54] & ~t[55]);
  assign t[44] = (t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[59]);
  assign t[46] = (t[60] & ~t[61]);
  assign t[47] = (t[62] & ~t[63]);
  assign t[48] = t[64] ^ x[2];
  assign t[49] = t[65] ^ x[1];
  assign t[4] = ~(t[25]);
  assign t[50] = t[66] ^ x[5];
  assign t[51] = t[67] ^ x[4];
  assign t[52] = t[68] ^ x[8];
  assign t[53] = t[69] ^ x[7];
  assign t[54] = t[70] ^ x[11];
  assign t[55] = t[71] ^ x[10];
  assign t[56] = t[72] ^ x[16];
  assign t[57] = t[73] ^ x[15];
  assign t[58] = t[74] ^ x[19];
  assign t[59] = t[75] ^ x[18];
  assign t[5] = ~(t[26] & t[8]);
  assign t[60] = t[76] ^ x[22];
  assign t[61] = t[77] ^ x[21];
  assign t[62] = t[78] ^ x[25];
  assign t[63] = t[79] ^ x[24];
  assign t[64] = (x[0]);
  assign t[65] = (x[0]);
  assign t[66] = (x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[26] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[14]);
  assign t[73] = (x[14]);
  assign t[74] = (x[17]);
  assign t[75] = (x[17]);
  assign t[76] = (x[20]);
  assign t[77] = (x[20]);
  assign t[78] = (x[23]);
  assign t[79] = (x[23]);
  assign t[7] = ~(t[27]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind337(x, y);
 input [25:0] x;
 output y;

 wire [79:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] & t[13]);
  assign t[11] = ~(t[14] & t[15]);
  assign t[12] = ~(t[28] | t[16]);
  assign t[13] = ~(t[29] & t[17]);
  assign t[14] = ~(t[18] | t[19]);
  assign t[15] = t[30] ? t[13] : t[29];
  assign t[16] = ~(t[20] | t[21]);
  assign t[17] = ~(t[22] & t[19]);
  assign t[18] = ~(t[30] | t[31]);
  assign t[19] = ~(t[28]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = ~(t[30]);
  assign t[21] = ~(t[22] & t[23]);
  assign t[22] = ~(t[31]);
  assign t[23] = ~(t[29]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = (t[36]);
  assign t[29] = (t[37]);
  assign t[2] = ~(t[6] & t[24]);
  assign t[30] = (t[38]);
  assign t[31] = (t[39]);
  assign t[32] = t[40] ^ x[2];
  assign t[33] = t[41] ^ x[5];
  assign t[34] = t[42] ^ x[8];
  assign t[35] = t[43] ^ x[11];
  assign t[36] = t[44] ^ x[16];
  assign t[37] = t[45] ^ x[19];
  assign t[38] = t[46] ^ x[22];
  assign t[39] = t[47] ^ x[25];
  assign t[3] = ~(t[7]);
  assign t[40] = (t[48] & ~t[49]);
  assign t[41] = (t[50] & ~t[51]);
  assign t[42] = (t[52] & ~t[53]);
  assign t[43] = (t[54] & ~t[55]);
  assign t[44] = (t[56] & ~t[57]);
  assign t[45] = (t[58] & ~t[59]);
  assign t[46] = (t[60] & ~t[61]);
  assign t[47] = (t[62] & ~t[63]);
  assign t[48] = t[64] ^ x[2];
  assign t[49] = t[65] ^ x[1];
  assign t[4] = ~(t[25]);
  assign t[50] = t[66] ^ x[5];
  assign t[51] = t[67] ^ x[4];
  assign t[52] = t[68] ^ x[8];
  assign t[53] = t[69] ^ x[7];
  assign t[54] = t[70] ^ x[11];
  assign t[55] = t[71] ^ x[10];
  assign t[56] = t[72] ^ x[16];
  assign t[57] = t[73] ^ x[15];
  assign t[58] = t[74] ^ x[19];
  assign t[59] = t[75] ^ x[18];
  assign t[5] = ~(t[26] & t[8]);
  assign t[60] = t[76] ^ x[22];
  assign t[61] = t[77] ^ x[21];
  assign t[62] = t[78] ^ x[25];
  assign t[63] = t[79] ^ x[24];
  assign t[64] = (x[0]);
  assign t[65] = (x[0]);
  assign t[66] = (x[3]);
  assign t[67] = (x[3]);
  assign t[68] = (x[6]);
  assign t[69] = (x[6]);
  assign t[6] = ~(t[26] | t[7]);
  assign t[70] = (x[9]);
  assign t[71] = (x[9]);
  assign t[72] = (x[14]);
  assign t[73] = (x[14]);
  assign t[74] = (x[17]);
  assign t[75] = (x[17]);
  assign t[76] = (x[20]);
  assign t[77] = (x[20]);
  assign t[78] = (x[23]);
  assign t[79] = (x[23]);
  assign t[7] = ~(t[27]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = ~(t[10] & t[11]);
  assign y = (t[0]);
endmodule

module R2ind338(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[14]);
  assign t[13] = t[24] ? t[17] : t[25];
  assign t[14] = ~(t[26]);
  assign t[15] = ~(t[24] ^ t[27]);
  assign t[16] = ~(t[24] | t[27]);
  assign t[17] = ~(t[25] & t[18]);
  assign t[18] = ~(t[19] & t[14]);
  assign t[19] = ~(t[27]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = t[36] ^ x[2];
  assign t[29] = t[37] ^ x[5];
  assign t[2] = ~(t[6] & t[20]);
  assign t[30] = t[38] ^ x[8];
  assign t[31] = t[39] ^ x[11];
  assign t[32] = t[40] ^ x[16];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[45]);
  assign t[37] = (t[46] & ~t[47]);
  assign t[38] = (t[48] & ~t[49]);
  assign t[39] = (t[50] & ~t[51]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[1];
  assign t[46] = t[62] ^ x[5];
  assign t[47] = t[63] ^ x[4];
  assign t[48] = t[64] ^ x[8];
  assign t[49] = t[65] ^ x[7];
  assign t[4] = ~(t[21]);
  assign t[50] = t[66] ^ x[11];
  assign t[51] = t[67] ^ x[10];
  assign t[52] = t[68] ^ x[16];
  assign t[53] = t[69] ^ x[15];
  assign t[54] = t[70] ^ x[19];
  assign t[55] = t[71] ^ x[18];
  assign t[56] = t[72] ^ x[22];
  assign t[57] = t[73] ^ x[21];
  assign t[58] = t[74] ^ x[25];
  assign t[59] = t[75] ^ x[24];
  assign t[5] = ~(t[22] & t[8]);
  assign t[60] = (x[0]);
  assign t[61] = (x[0]);
  assign t[62] = (x[3]);
  assign t[63] = (x[3]);
  assign t[64] = (x[6]);
  assign t[65] = (x[6]);
  assign t[66] = (x[9]);
  assign t[67] = (x[9]);
  assign t[68] = (x[14]);
  assign t[69] = (x[14]);
  assign t[6] = ~(t[22] | t[7]);
  assign t[70] = (x[17]);
  assign t[71] = (x[17]);
  assign t[72] = (x[20]);
  assign t[73] = (x[20]);
  assign t[74] = (x[23]);
  assign t[75] = (x[23]);
  assign t[7] = ~(t[23]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = ~(t[10] | t[11]);
  assign y = (t[0]);
endmodule

module R2ind339(x, y);
 input [25:0] x;
 output y;

 wire [75:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] | t[13]);
  assign t[11] = ~(t[14] | t[15]);
  assign t[12] = ~(t[16] | t[14]);
  assign t[13] = t[24] ? t[17] : t[25];
  assign t[14] = ~(t[26]);
  assign t[15] = ~(t[24] ^ t[27]);
  assign t[16] = ~(t[24] | t[27]);
  assign t[17] = ~(t[25] & t[18]);
  assign t[18] = ~(t[19] & t[14]);
  assign t[19] = ~(t[27]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = (t[29]);
  assign t[22] = (t[30]);
  assign t[23] = (t[31]);
  assign t[24] = (t[32]);
  assign t[25] = (t[33]);
  assign t[26] = (t[34]);
  assign t[27] = (t[35]);
  assign t[28] = t[36] ^ x[2];
  assign t[29] = t[37] ^ x[5];
  assign t[2] = ~(t[6] & t[20]);
  assign t[30] = t[38] ^ x[8];
  assign t[31] = t[39] ^ x[11];
  assign t[32] = t[40] ^ x[16];
  assign t[33] = t[41] ^ x[19];
  assign t[34] = t[42] ^ x[22];
  assign t[35] = t[43] ^ x[25];
  assign t[36] = (t[44] & ~t[45]);
  assign t[37] = (t[46] & ~t[47]);
  assign t[38] = (t[48] & ~t[49]);
  assign t[39] = (t[50] & ~t[51]);
  assign t[3] = ~(t[7]);
  assign t[40] = (t[52] & ~t[53]);
  assign t[41] = (t[54] & ~t[55]);
  assign t[42] = (t[56] & ~t[57]);
  assign t[43] = (t[58] & ~t[59]);
  assign t[44] = t[60] ^ x[2];
  assign t[45] = t[61] ^ x[1];
  assign t[46] = t[62] ^ x[5];
  assign t[47] = t[63] ^ x[4];
  assign t[48] = t[64] ^ x[8];
  assign t[49] = t[65] ^ x[7];
  assign t[4] = ~(t[21]);
  assign t[50] = t[66] ^ x[11];
  assign t[51] = t[67] ^ x[10];
  assign t[52] = t[68] ^ x[16];
  assign t[53] = t[69] ^ x[15];
  assign t[54] = t[70] ^ x[19];
  assign t[55] = t[71] ^ x[18];
  assign t[56] = t[72] ^ x[22];
  assign t[57] = t[73] ^ x[21];
  assign t[58] = t[74] ^ x[25];
  assign t[59] = t[75] ^ x[24];
  assign t[5] = ~(t[22] & t[8]);
  assign t[60] = (x[0]);
  assign t[61] = (x[0]);
  assign t[62] = (x[3]);
  assign t[63] = (x[3]);
  assign t[64] = (x[6]);
  assign t[65] = (x[6]);
  assign t[66] = (x[9]);
  assign t[67] = (x[9]);
  assign t[68] = (x[14]);
  assign t[69] = (x[14]);
  assign t[6] = ~(t[22] | t[7]);
  assign t[70] = (x[17]);
  assign t[71] = (x[17]);
  assign t[72] = (x[20]);
  assign t[73] = (x[20]);
  assign t[74] = (x[23]);
  assign t[75] = (x[23]);
  assign t[7] = ~(t[23]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = ~(t[10] | t[11]);
  assign y = (t[0]);
endmodule

module R2ind340(x, y);
 input [25:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] | t[17]);
  assign t[11] = ~(t[18] ^ t[19]);
  assign t[12] = ~(t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = t[29] ^ x[2];
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[8];
  assign t[24] = t[32] ^ x[11];
  assign t[25] = t[33] ^ x[16];
  assign t[26] = t[34] ^ x[19];
  assign t[27] = t[35] ^ x[22];
  assign t[28] = t[36] ^ x[25];
  assign t[29] = (t[37] & ~t[38]);
  assign t[2] = ~(t[6] & t[13]);
  assign t[30] = (t[39] & ~t[40]);
  assign t[31] = (t[41] & ~t[42]);
  assign t[32] = (t[43] & ~t[44]);
  assign t[33] = (t[45] & ~t[46]);
  assign t[34] = (t[47] & ~t[48]);
  assign t[35] = (t[49] & ~t[50]);
  assign t[36] = (t[51] & ~t[52]);
  assign t[37] = t[53] ^ x[2];
  assign t[38] = t[54] ^ x[1];
  assign t[39] = t[55] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[56] ^ x[4];
  assign t[41] = t[57] ^ x[8];
  assign t[42] = t[58] ^ x[7];
  assign t[43] = t[59] ^ x[11];
  assign t[44] = t[60] ^ x[10];
  assign t[45] = t[61] ^ x[16];
  assign t[46] = t[62] ^ x[15];
  assign t[47] = t[63] ^ x[19];
  assign t[48] = t[64] ^ x[18];
  assign t[49] = t[65] ^ x[22];
  assign t[4] = ~(t[14]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[25];
  assign t[52] = t[68] ^ x[24];
  assign t[53] = (x[0]);
  assign t[54] = (x[0]);
  assign t[55] = (x[3]);
  assign t[56] = (x[3]);
  assign t[57] = (x[6]);
  assign t[58] = (x[6]);
  assign t[59] = (x[9]);
  assign t[5] = ~(t[15] & t[8]);
  assign t[60] = (x[9]);
  assign t[61] = (x[14]);
  assign t[62] = (x[14]);
  assign t[63] = (x[17]);
  assign t[64] = (x[17]);
  assign t[65] = (x[20]);
  assign t[66] = (x[20]);
  assign t[67] = (x[23]);
  assign t[68] = (x[23]);
  assign t[6] = ~(t[15] | t[7]);
  assign t[7] = ~(t[16]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = ~(t[10] ^ t[11]);
  assign y = (t[0]);
endmodule

module R2ind341(x, y);
 input [25:0] x;
 output y;

 wire [68:0] t;
  assign t[0] = ~(t[1] & t[2]);
  assign t[10] = ~(t[12] | t[17]);
  assign t[11] = ~(t[18] ^ t[19]);
  assign t[12] = ~(t[20]);
  assign t[13] = (t[21]);
  assign t[14] = (t[22]);
  assign t[15] = (t[23]);
  assign t[16] = (t[24]);
  assign t[17] = (t[25]);
  assign t[18] = (t[26]);
  assign t[19] = (t[27]);
  assign t[1] = t[3] ? t[5] : t[4];
  assign t[20] = (t[28]);
  assign t[21] = t[29] ^ x[2];
  assign t[22] = t[30] ^ x[5];
  assign t[23] = t[31] ^ x[8];
  assign t[24] = t[32] ^ x[11];
  assign t[25] = t[33] ^ x[16];
  assign t[26] = t[34] ^ x[19];
  assign t[27] = t[35] ^ x[22];
  assign t[28] = t[36] ^ x[25];
  assign t[29] = (t[37] & ~t[38]);
  assign t[2] = ~(t[6] & t[13]);
  assign t[30] = (t[39] & ~t[40]);
  assign t[31] = (t[41] & ~t[42]);
  assign t[32] = (t[43] & ~t[44]);
  assign t[33] = (t[45] & ~t[46]);
  assign t[34] = (t[47] & ~t[48]);
  assign t[35] = (t[49] & ~t[50]);
  assign t[36] = (t[51] & ~t[52]);
  assign t[37] = t[53] ^ x[2];
  assign t[38] = t[54] ^ x[1];
  assign t[39] = t[55] ^ x[5];
  assign t[3] = ~(t[7]);
  assign t[40] = t[56] ^ x[4];
  assign t[41] = t[57] ^ x[8];
  assign t[42] = t[58] ^ x[7];
  assign t[43] = t[59] ^ x[11];
  assign t[44] = t[60] ^ x[10];
  assign t[45] = t[61] ^ x[16];
  assign t[46] = t[62] ^ x[15];
  assign t[47] = t[63] ^ x[19];
  assign t[48] = t[64] ^ x[18];
  assign t[49] = t[65] ^ x[22];
  assign t[4] = ~(t[14]);
  assign t[50] = t[66] ^ x[21];
  assign t[51] = t[67] ^ x[25];
  assign t[52] = t[68] ^ x[24];
  assign t[53] = (x[0]);
  assign t[54] = (x[0]);
  assign t[55] = (x[3]);
  assign t[56] = (x[3]);
  assign t[57] = (x[6]);
  assign t[58] = (x[6]);
  assign t[59] = (x[9]);
  assign t[5] = ~(t[15] & t[8]);
  assign t[60] = (x[9]);
  assign t[61] = (x[14]);
  assign t[62] = (x[14]);
  assign t[63] = (x[17]);
  assign t[64] = (x[17]);
  assign t[65] = (x[20]);
  assign t[66] = (x[20]);
  assign t[67] = (x[23]);
  assign t[68] = (x[23]);
  assign t[6] = ~(t[15] | t[7]);
  assign t[7] = ~(t[16]);
  assign t[8] = x[12] ? x[13] : t[9];
  assign t[9] = ~(t[10] ^ t[11]);
  assign y = (t[0]);
endmodule

module R2ind342(x, y);
 input [20:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[2];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[8];
  assign t[18] = t[25] ^ x[11];
  assign t[19] = t[26] ^ x[14];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[17];
  assign t[21] = t[28] ^ x[20];
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = (t[35] & ~t[36]);
  assign t[26] = (t[37] & ~t[38]);
  assign t[27] = (t[39] & ~t[40]);
  assign t[28] = (t[41] & ~t[42]);
  assign t[29] = t[43] ^ x[2];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[1];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[4];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[7];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[10];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[13];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[16];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = (x[0]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[46] = (x[3]);
  assign t[47] = (x[6]);
  assign t[48] = (x[6]);
  assign t[49] = (x[9]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[9]);
  assign t[51] = (x[12]);
  assign t[52] = (x[12]);
  assign t[53] = (x[15]);
  assign t[54] = (x[15]);
  assign t[55] = (x[18]);
  assign t[56] = (x[18]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind343(x, y);
 input [20:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[2];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[8];
  assign t[18] = t[25] ^ x[11];
  assign t[19] = t[26] ^ x[14];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[17];
  assign t[21] = t[28] ^ x[20];
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = (t[35] & ~t[36]);
  assign t[26] = (t[37] & ~t[38]);
  assign t[27] = (t[39] & ~t[40]);
  assign t[28] = (t[41] & ~t[42]);
  assign t[29] = t[43] ^ x[2];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[1];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[4];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[7];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[10];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[13];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[16];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = (x[0]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[46] = (x[3]);
  assign t[47] = (x[6]);
  assign t[48] = (x[6]);
  assign t[49] = (x[9]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[9]);
  assign t[51] = (x[12]);
  assign t[52] = (x[12]);
  assign t[53] = (x[15]);
  assign t[54] = (x[15]);
  assign t[55] = (x[18]);
  assign t[56] = (x[18]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind344(x, y);
 input [20:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[2];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[8];
  assign t[18] = t[25] ^ x[11];
  assign t[19] = t[26] ^ x[14];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[17];
  assign t[21] = t[28] ^ x[20];
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = (t[35] & ~t[36]);
  assign t[26] = (t[37] & ~t[38]);
  assign t[27] = (t[39] & ~t[40]);
  assign t[28] = (t[41] & ~t[42]);
  assign t[29] = t[43] ^ x[2];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[1];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[4];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[7];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[10];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[13];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[16];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = (x[0]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[46] = (x[3]);
  assign t[47] = (x[6]);
  assign t[48] = (x[6]);
  assign t[49] = (x[9]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[9]);
  assign t[51] = (x[12]);
  assign t[52] = (x[12]);
  assign t[53] = (x[15]);
  assign t[54] = (x[15]);
  assign t[55] = (x[18]);
  assign t[56] = (x[18]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind345(x, y);
 input [20:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[2];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[8];
  assign t[18] = t[25] ^ x[11];
  assign t[19] = t[26] ^ x[14];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[17];
  assign t[21] = t[28] ^ x[20];
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = (t[35] & ~t[36]);
  assign t[26] = (t[37] & ~t[38]);
  assign t[27] = (t[39] & ~t[40]);
  assign t[28] = (t[41] & ~t[42]);
  assign t[29] = t[43] ^ x[2];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[1];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[4];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[7];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[10];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[13];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[16];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = (x[0]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[46] = (x[3]);
  assign t[47] = (x[6]);
  assign t[48] = (x[6]);
  assign t[49] = (x[9]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[9]);
  assign t[51] = (x[12]);
  assign t[52] = (x[12]);
  assign t[53] = (x[15]);
  assign t[54] = (x[15]);
  assign t[55] = (x[18]);
  assign t[56] = (x[18]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind346(x, y);
 input [20:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[2];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[8];
  assign t[18] = t[25] ^ x[11];
  assign t[19] = t[26] ^ x[14];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[17];
  assign t[21] = t[28] ^ x[20];
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = (t[35] & ~t[36]);
  assign t[26] = (t[37] & ~t[38]);
  assign t[27] = (t[39] & ~t[40]);
  assign t[28] = (t[41] & ~t[42]);
  assign t[29] = t[43] ^ x[2];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[1];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[4];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[7];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[10];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[13];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[16];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = (x[0]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[46] = (x[3]);
  assign t[47] = (x[6]);
  assign t[48] = (x[6]);
  assign t[49] = (x[9]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[9]);
  assign t[51] = (x[12]);
  assign t[52] = (x[12]);
  assign t[53] = (x[15]);
  assign t[54] = (x[15]);
  assign t[55] = (x[18]);
  assign t[56] = (x[18]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind347(x, y);
 input [20:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[2];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[8];
  assign t[18] = t[25] ^ x[11];
  assign t[19] = t[26] ^ x[14];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[17];
  assign t[21] = t[28] ^ x[20];
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = (t[35] & ~t[36]);
  assign t[26] = (t[37] & ~t[38]);
  assign t[27] = (t[39] & ~t[40]);
  assign t[28] = (t[41] & ~t[42]);
  assign t[29] = t[43] ^ x[2];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[1];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[4];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[7];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[10];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[13];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[16];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = (x[0]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[46] = (x[3]);
  assign t[47] = (x[6]);
  assign t[48] = (x[6]);
  assign t[49] = (x[9]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[9]);
  assign t[51] = (x[12]);
  assign t[52] = (x[12]);
  assign t[53] = (x[15]);
  assign t[54] = (x[15]);
  assign t[55] = (x[18]);
  assign t[56] = (x[18]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind348(x, y);
 input [20:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[2];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[8];
  assign t[18] = t[25] ^ x[11];
  assign t[19] = t[26] ^ x[14];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[17];
  assign t[21] = t[28] ^ x[20];
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = (t[35] & ~t[36]);
  assign t[26] = (t[37] & ~t[38]);
  assign t[27] = (t[39] & ~t[40]);
  assign t[28] = (t[41] & ~t[42]);
  assign t[29] = t[43] ^ x[2];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[1];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[4];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[7];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[10];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[13];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[16];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = (x[0]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[46] = (x[3]);
  assign t[47] = (x[6]);
  assign t[48] = (x[6]);
  assign t[49] = (x[9]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[9]);
  assign t[51] = (x[12]);
  assign t[52] = (x[12]);
  assign t[53] = (x[15]);
  assign t[54] = (x[15]);
  assign t[55] = (x[18]);
  assign t[56] = (x[18]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2ind349(x, y);
 input [20:0] x;
 output y;

 wire [56:0] t;
  assign t[0] = t[1] ? t[8] : t[2];
  assign t[10] = (t[17]);
  assign t[11] = (t[18]);
  assign t[12] = (t[19]);
  assign t[13] = (t[20]);
  assign t[14] = (t[21]);
  assign t[15] = t[22] ^ x[2];
  assign t[16] = t[23] ^ x[5];
  assign t[17] = t[24] ^ x[8];
  assign t[18] = t[25] ^ x[11];
  assign t[19] = t[26] ^ x[14];
  assign t[1] = ~(t[3] | t[4]);
  assign t[20] = t[27] ^ x[17];
  assign t[21] = t[28] ^ x[20];
  assign t[22] = (t[29] & ~t[30]);
  assign t[23] = (t[31] & ~t[32]);
  assign t[24] = (t[33] & ~t[34]);
  assign t[25] = (t[35] & ~t[36]);
  assign t[26] = (t[37] & ~t[38]);
  assign t[27] = (t[39] & ~t[40]);
  assign t[28] = (t[41] & ~t[42]);
  assign t[29] = t[43] ^ x[2];
  assign t[2] = t[9] ^ t[10];
  assign t[30] = t[44] ^ x[1];
  assign t[31] = t[45] ^ x[5];
  assign t[32] = t[46] ^ x[4];
  assign t[33] = t[47] ^ x[8];
  assign t[34] = t[48] ^ x[7];
  assign t[35] = t[49] ^ x[11];
  assign t[36] = t[50] ^ x[10];
  assign t[37] = t[51] ^ x[14];
  assign t[38] = t[52] ^ x[13];
  assign t[39] = t[53] ^ x[17];
  assign t[3] = ~(t[5] & t[6]);
  assign t[40] = t[54] ^ x[16];
  assign t[41] = t[55] ^ x[20];
  assign t[42] = t[56] ^ x[19];
  assign t[43] = (x[0]);
  assign t[44] = (x[0]);
  assign t[45] = (x[3]);
  assign t[46] = (x[3]);
  assign t[47] = (x[6]);
  assign t[48] = (x[6]);
  assign t[49] = (x[9]);
  assign t[4] = ~(t[11] & t[7]);
  assign t[50] = (x[9]);
  assign t[51] = (x[12]);
  assign t[52] = (x[12]);
  assign t[53] = (x[15]);
  assign t[54] = (x[15]);
  assign t[55] = (x[18]);
  assign t[56] = (x[18]);
  assign t[5] = ~(t[12]);
  assign t[6] = ~(t[13]);
  assign t[7] = ~(t[14]);
  assign t[8] = (t[15]);
  assign t[9] = (t[16]);
  assign y = (t[0]);
endmodule

module R2_ind(x, y);
 input [666:0] x;
 output [349:0] y;

  R2ind0 R2ind0_inst(.x({x[2], x[1], x[0]}), .y(y[0]));
  R2ind1 R2ind1_inst(.x({x[1], x[2], x[0]}), .y(y[1]));
  R2ind2 R2ind2_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[2]));
  R2ind3 R2ind3_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3]}), .y(y[3]));
  R2ind4 R2ind4_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30]}), .y(y[4]));
  R2ind5 R2ind5_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30]}), .y(y[5]));
  R2ind6 R2ind6_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[8], x[7], x[6], x[11], x[10], x[9], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[6]));
  R2ind7 R2ind7_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[8], x[7], x[6], x[11], x[10], x[9], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[30]}), .y(y[7]));
  R2ind8 R2ind8_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[30]}), .y(y[8]));
  R2ind9 R2ind9_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[17], x[16], x[15], x[14], x[13], x[12], x[11], x[10], x[9], x[8], x[7], x[6], x[5], x[4], x[3], x[30]}), .y(y[9]));
  R2ind10 R2ind10_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[5], x[4], x[3], x[14], x[13], x[12], x[30]}), .y(y[10]));
  R2ind11 R2ind11_inst(.x({x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6], x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[45], x[44], x[43], x[42], x[41], x[40], x[39], x[38], x[37], x[36], x[35], x[34], x[33], x[32], x[31], x[5], x[4], x[3], x[14], x[13], x[12], x[30]}), .y(y[11]));
  R2ind12 R2ind12_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[33], x[32], x[31], x[39], x[38], x[37], x[36], x[35], x[34], x[30], x[42], x[41], x[40]}), .y(y[12]));
  R2ind13 R2ind13_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[33], x[32], x[31], x[39], x[38], x[37], x[36], x[35], x[34], x[30], x[42], x[41], x[40]}), .y(y[13]));
  R2ind14 R2ind14_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[30], x[33], x[32], x[31], x[39], x[38], x[37]}), .y(y[14]));
  R2ind15 R2ind15_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[30], x[33], x[32], x[31], x[39], x[38], x[37]}), .y(y[15]));
  R2ind16 R2ind16_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[45], x[44], x[43], x[33], x[32], x[31]}), .y(y[16]));
  R2ind17 R2ind17_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[45], x[44], x[43], x[33], x[32], x[31]}), .y(y[17]));
  R2ind18 R2ind18_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[45], x[44], x[43]}), .y(y[18]));
  R2ind19 R2ind19_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[30], x[45], x[44], x[43]}), .y(y[19]));
  R2ind20 R2ind20_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[33], x[32], x[31], x[39], x[38], x[37], x[30], x[36], x[35], x[34]}), .y(y[20]));
  R2ind21 R2ind21_inst(.x({x[29], x[28], x[27], x[26], x[25], x[24], x[23], x[22], x[21], x[20], x[19], x[18], x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[45], x[44], x[43], x[33], x[32], x[31], x[39], x[38], x[37], x[30], x[36], x[35], x[34]}), .y(y[21]));
  R2ind22 R2ind22_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[26], x[25], x[24], x[29], x[28], x[27], x[48], x[47], x[46], x[20], x[19], x[18]}), .y(y[22]));
  R2ind23 R2ind23_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[26], x[25], x[24], x[29], x[28], x[27], x[48], x[47], x[46], x[20], x[19], x[18]}), .y(y[23]));
  R2ind24 R2ind24_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[26], x[25], x[24], x[29], x[28], x[27], x[20], x[19], x[18], x[48], x[47], x[46], x[23], x[22], x[21]}), .y(y[24]));
  R2ind25 R2ind25_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[26], x[25], x[24], x[29], x[28], x[27], x[20], x[19], x[18], x[48], x[47], x[46], x[23], x[22], x[21]}), .y(y[25]));
  R2ind26 R2ind26_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[26], x[25], x[24], x[48], x[47], x[46], x[29], x[28], x[27]}), .y(y[26]));
  R2ind27 R2ind27_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[26], x[25], x[24], x[48], x[47], x[46], x[29], x[28], x[27]}), .y(y[27]));
  R2ind28 R2ind28_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[26], x[25], x[24], x[48], x[47], x[46]}), .y(y[28]));
  R2ind29 R2ind29_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[5], x[4], x[3], x[26], x[25], x[24], x[48], x[47], x[46]}), .y(y[29]));
  R2ind30 R2ind30_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[30]));
  R2ind31 R2ind31_inst(.x({x[14], x[13], x[12], x[17], x[16], x[15], x[11], x[10], x[9], x[8], x[7], x[6]}), .y(y[31]));
  R2ind32 R2ind32_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[30]}), .y(y[32]));
  R2ind33 R2ind33_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[30]}), .y(y[33]));
  R2ind34 R2ind34_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[48], x[47], x[46], x[5], x[4], x[3]}), .y(y[34]));
  R2ind35 R2ind35_inst(.x({x[11], x[10], x[9], x[8], x[7], x[6], x[14], x[13], x[12], x[17], x[16], x[15], x[48], x[47], x[46], x[5], x[4], x[3]}), .y(y[35]));
  R2ind36 R2ind36_inst(.x({x[48], x[47], x[46]}), .y(y[36]));
  R2ind37 R2ind37_inst(.x({x[48], x[47], x[46]}), .y(y[37]));
  R2ind38 R2ind38_inst(.x({x[48], x[47], x[46]}), .y(y[38]));
  R2ind39 R2ind39_inst(.x({x[48], x[47], x[46]}), .y(y[39]));
  R2ind40 R2ind40_inst(.x({x[51], x[50], x[49]}), .y(y[40]));
  R2ind41 R2ind41_inst(.x({x[51], x[50], x[49]}), .y(y[41]));
  R2ind42 R2ind42_inst(.x({x[51], x[50], x[49]}), .y(y[42]));
  R2ind43 R2ind43_inst(.x({x[51], x[50], x[49]}), .y(y[43]));
  R2ind44 R2ind44_inst(.x({x[54], x[53], x[52]}), .y(y[44]));
  R2ind45 R2ind45_inst(.x({x[54], x[53], x[52]}), .y(y[45]));
  R2ind46 R2ind46_inst(.x({x[57], x[56], x[55]}), .y(y[46]));
  R2ind47 R2ind47_inst(.x({x[57], x[56], x[55]}), .y(y[47]));
  R2ind48 R2ind48_inst(.x({x[57], x[56], x[55]}), .y(y[48]));
  R2ind49 R2ind49_inst(.x({x[57], x[56], x[55]}), .y(y[49]));
  R2ind50 R2ind50_inst(.x({x[60], x[59], x[58]}), .y(y[50]));
  R2ind51 R2ind51_inst(.x({x[60], x[59], x[58]}), .y(y[51]));
  R2ind52 R2ind52_inst(.x({x[60], x[59], x[58]}), .y(y[52]));
  R2ind53 R2ind53_inst(.x({x[60], x[59], x[58]}), .y(y[53]));
  R2ind54 R2ind54_inst(.x({x[82], x[81], x[80], x[30], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[5], x[4], x[3], x[48], x[47], x[46], x[63], x[62], x[61], x[54], x[53], x[52]}), .y(y[54]));
  R2ind55 R2ind55_inst(.x({x[82], x[81], x[80], x[30], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[70], x[69], x[68], x[67], x[66], x[65], x[64], x[5], x[4], x[3], x[48], x[47], x[46], x[63], x[62], x[61], x[54], x[53], x[52]}), .y(y[55]));
  R2ind56 R2ind56_inst(.x({x[79], x[78], x[77], x[82], x[81], x[80], x[73], x[72], x[71], x[76], x[75], x[74], x[30], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[5], x[4], x[3], x[48], x[47], x[46], x[85], x[84], x[83], x[54], x[53], x[52]}), .y(y[56]));
  R2ind57 R2ind57_inst(.x({x[79], x[78], x[77], x[82], x[81], x[80], x[73], x[72], x[71], x[76], x[75], x[74], x[30], x[95], x[94], x[93], x[92], x[91], x[90], x[89], x[88], x[87], x[86], x[5], x[4], x[3], x[48], x[47], x[46], x[85], x[84], x[83], x[54], x[53], x[52]}), .y(y[57]));
  R2ind58 R2ind58_inst(.x({x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[82], x[81], x[80], x[30], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[5], x[4], x[3], x[48], x[47], x[46], x[98], x[97], x[96], x[54], x[53], x[52]}), .y(y[58]));
  R2ind59 R2ind59_inst(.x({x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[82], x[81], x[80], x[30], x[108], x[107], x[106], x[105], x[104], x[103], x[102], x[101], x[100], x[99], x[5], x[4], x[3], x[48], x[47], x[46], x[98], x[97], x[96], x[54], x[53], x[52]}), .y(y[59]));
  R2ind60 R2ind60_inst(.x({x[82], x[81], x[80], x[79], x[78], x[77], x[73], x[72], x[71], x[30], x[76], x[75], x[74], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[5], x[4], x[3], x[48], x[47], x[46], x[111], x[110], x[109], x[54], x[53], x[52]}), .y(y[60]));
  R2ind61 R2ind61_inst(.x({x[82], x[81], x[80], x[79], x[78], x[77], x[73], x[72], x[71], x[30], x[76], x[75], x[74], x[121], x[120], x[119], x[118], x[117], x[116], x[115], x[114], x[113], x[112], x[5], x[4], x[3], x[48], x[47], x[46], x[111], x[110], x[109], x[54], x[53], x[52]}), .y(y[61]));
  R2ind62 R2ind62_inst(.x({x[30], x[128], x[127], x[126], x[125], x[54], x[53], x[52], x[48], x[47], x[46], x[124], x[123], x[122], x[111], x[110], x[109]}), .y(y[62]));
  R2ind63 R2ind63_inst(.x({x[30], x[128], x[127], x[126], x[125], x[54], x[53], x[52], x[48], x[47], x[46], x[124], x[123], x[122], x[111], x[110], x[109]}), .y(y[63]));
  R2ind64 R2ind64_inst(.x({x[30], x[135], x[134], x[133], x[132], x[54], x[53], x[52], x[48], x[47], x[46], x[131], x[130], x[129], x[98], x[97], x[96]}), .y(y[64]));
  R2ind65 R2ind65_inst(.x({x[30], x[135], x[134], x[133], x[132], x[54], x[53], x[52], x[48], x[47], x[46], x[131], x[130], x[129], x[98], x[97], x[96]}), .y(y[65]));
  R2ind66 R2ind66_inst(.x({x[30], x[142], x[141], x[140], x[139], x[54], x[53], x[52], x[48], x[47], x[46], x[138], x[137], x[136], x[85], x[84], x[83]}), .y(y[66]));
  R2ind67 R2ind67_inst(.x({x[30], x[142], x[141], x[140], x[139], x[54], x[53], x[52], x[48], x[47], x[46], x[138], x[137], x[136], x[85], x[84], x[83]}), .y(y[67]));
  R2ind68 R2ind68_inst(.x({x[30], x[146], x[145], x[144], x[143], x[54], x[53], x[52], x[48], x[47], x[46], x[88], x[87], x[86], x[63], x[62], x[61]}), .y(y[68]));
  R2ind69 R2ind69_inst(.x({x[30], x[146], x[145], x[144], x[143], x[54], x[53], x[52], x[48], x[47], x[46], x[88], x[87], x[86], x[63], x[62], x[61]}), .y(y[69]));
  R2ind70 R2ind70_inst(.x({x[30], x[156], x[155], x[154], x[153], x[54], x[53], x[52], x[152], x[151], x[150], x[149], x[148], x[147], x[124], x[123], x[122]}), .y(y[70]));
  R2ind71 R2ind71_inst(.x({x[30], x[156], x[155], x[154], x[153], x[54], x[53], x[52], x[152], x[151], x[150], x[149], x[148], x[147], x[124], x[123], x[122]}), .y(y[71]));
  R2ind72 R2ind72_inst(.x({x[30], x[163], x[162], x[161], x[160], x[54], x[53], x[52], x[152], x[151], x[150], x[159], x[158], x[157], x[131], x[130], x[129]}), .y(y[72]));
  R2ind73 R2ind73_inst(.x({x[30], x[163], x[162], x[161], x[160], x[54], x[53], x[52], x[152], x[151], x[150], x[159], x[158], x[157], x[131], x[130], x[129]}), .y(y[73]));
  R2ind74 R2ind74_inst(.x({x[30], x[170], x[169], x[168], x[167], x[54], x[53], x[52], x[152], x[151], x[150], x[166], x[165], x[164], x[138], x[137], x[136]}), .y(y[74]));
  R2ind75 R2ind75_inst(.x({x[30], x[170], x[169], x[168], x[167], x[54], x[53], x[52], x[152], x[151], x[150], x[166], x[165], x[164], x[138], x[137], x[136]}), .y(y[75]));
  R2ind76 R2ind76_inst(.x({x[30], x[174], x[173], x[172], x[171], x[54], x[53], x[52], x[152], x[151], x[150], x[101], x[100], x[99], x[88], x[87], x[86]}), .y(y[76]));
  R2ind77 R2ind77_inst(.x({x[30], x[174], x[173], x[172], x[171], x[54], x[53], x[52], x[152], x[151], x[150], x[101], x[100], x[99], x[88], x[87], x[86]}), .y(y[77]));
  R2ind78 R2ind78_inst(.x({x[30], x[178], x[70], x[69], x[68], x[54], x[53], x[52], x[152], x[151], x[150], x[177], x[176], x[175], x[149], x[148], x[147]}), .y(y[78]));
  R2ind79 R2ind79_inst(.x({x[30], x[178], x[70], x[69], x[68], x[54], x[53], x[52], x[152], x[151], x[150], x[177], x[176], x[175], x[149], x[148], x[147]}), .y(y[79]));
  R2ind80 R2ind80_inst(.x({x[30], x[185], x[184], x[183], x[182], x[54], x[53], x[52], x[152], x[151], x[150], x[181], x[180], x[179], x[159], x[158], x[157]}), .y(y[80]));
  R2ind81 R2ind81_inst(.x({x[30], x[185], x[184], x[183], x[182], x[54], x[53], x[52], x[152], x[151], x[150], x[181], x[180], x[179], x[159], x[158], x[157]}), .y(y[81]));
  R2ind82 R2ind82_inst(.x({x[30], x[192], x[191], x[190], x[189], x[54], x[53], x[52], x[152], x[151], x[150], x[188], x[187], x[186], x[166], x[165], x[164]}), .y(y[82]));
  R2ind83 R2ind83_inst(.x({x[30], x[192], x[191], x[190], x[189], x[54], x[53], x[52], x[152], x[151], x[150], x[188], x[187], x[186], x[166], x[165], x[164]}), .y(y[83]));
  R2ind84 R2ind84_inst(.x({x[30], x[196], x[195], x[194], x[193], x[54], x[53], x[52], x[152], x[151], x[150], x[114], x[113], x[112], x[101], x[100], x[99]}), .y(y[84]));
  R2ind85 R2ind85_inst(.x({x[30], x[196], x[195], x[194], x[193], x[54], x[53], x[52], x[152], x[151], x[150], x[114], x[113], x[112], x[101], x[100], x[99]}), .y(y[85]));
  R2ind86 R2ind86_inst(.x({x[30], x[200], x[188], x[187], x[186], x[152], x[151], x[150], x[199], x[198], x[197], x[177], x[176], x[175], x[54], x[53], x[52]}), .y(y[86]));
  R2ind87 R2ind87_inst(.x({x[30], x[200], x[188], x[187], x[186], x[152], x[151], x[150], x[199], x[198], x[197], x[177], x[176], x[175], x[54], x[53], x[52]}), .y(y[87]));
  R2ind88 R2ind88_inst(.x({x[30], x[204], x[166], x[165], x[164], x[152], x[151], x[150], x[203], x[202], x[201], x[181], x[180], x[179], x[54], x[53], x[52]}), .y(y[88]));
  R2ind89 R2ind89_inst(.x({x[30], x[204], x[166], x[165], x[164], x[152], x[151], x[150], x[203], x[202], x[201], x[181], x[180], x[179], x[54], x[53], x[52]}), .y(y[89]));
  R2ind90 R2ind90_inst(.x({x[30], x[208], x[138], x[137], x[136], x[152], x[151], x[150], x[207], x[206], x[205], x[188], x[187], x[186], x[54], x[53], x[52]}), .y(y[90]));
  R2ind91 R2ind91_inst(.x({x[30], x[208], x[138], x[137], x[136], x[152], x[151], x[150], x[207], x[206], x[205], x[188], x[187], x[186], x[54], x[53], x[52]}), .y(y[91]));
  R2ind92 R2ind92_inst(.x({x[30], x[209], x[85], x[84], x[83], x[152], x[151], x[150], x[145], x[144], x[143], x[114], x[113], x[112], x[54], x[53], x[52]}), .y(y[92]));
  R2ind93 R2ind93_inst(.x({x[30], x[209], x[85], x[84], x[83], x[152], x[151], x[150], x[145], x[144], x[143], x[114], x[113], x[112], x[54], x[53], x[52]}), .y(y[93]));
  R2ind94 R2ind94_inst(.x({x[30], x[216], x[215], x[214], x[213], x[54], x[53], x[52], x[152], x[151], x[150], x[212], x[211], x[210], x[199], x[198], x[197]}), .y(y[94]));
  R2ind95 R2ind95_inst(.x({x[30], x[216], x[215], x[214], x[213], x[54], x[53], x[52], x[152], x[151], x[150], x[212], x[211], x[210], x[199], x[198], x[197]}), .y(y[95]));
  R2ind96 R2ind96_inst(.x({x[30], x[223], x[222], x[221], x[220], x[54], x[53], x[52], x[152], x[151], x[150], x[219], x[218], x[217], x[203], x[202], x[201]}), .y(y[96]));
  R2ind97 R2ind97_inst(.x({x[30], x[223], x[222], x[221], x[220], x[54], x[53], x[52], x[152], x[151], x[150], x[219], x[218], x[217], x[203], x[202], x[201]}), .y(y[97]));
  R2ind98 R2ind98_inst(.x({x[30], x[227], x[54], x[53], x[52], x[152], x[151], x[150], x[226], x[225], x[224], x[207], x[206], x[205]}), .y(y[98]));
  R2ind99 R2ind99_inst(.x({x[30], x[227], x[54], x[53], x[52], x[152], x[151], x[150], x[226], x[225], x[224], x[207], x[206], x[205]}), .y(y[99]));
  R2ind100 R2ind100_inst(.x({x[30], x[228], x[207], x[206], x[205], x[54], x[53], x[52], x[152], x[151], x[150], x[141], x[140], x[139], x[145], x[144], x[143]}), .y(y[100]));
  R2ind101 R2ind101_inst(.x({x[30], x[228], x[207], x[206], x[205], x[54], x[53], x[52], x[152], x[151], x[150], x[141], x[140], x[139], x[145], x[144], x[143]}), .y(y[101]));
  R2ind102 R2ind102_inst(.x({x[30], x[235], x[234], x[233], x[232], x[54], x[53], x[52], x[152], x[151], x[150], x[231], x[230], x[229], x[212], x[211], x[210]}), .y(y[102]));
  R2ind103 R2ind103_inst(.x({x[30], x[235], x[234], x[233], x[232], x[54], x[53], x[52], x[152], x[151], x[150], x[231], x[230], x[229], x[212], x[211], x[210]}), .y(y[103]));
  R2ind104 R2ind104_inst(.x({x[30], x[242], x[241], x[240], x[239], x[54], x[53], x[52], x[152], x[151], x[150], x[238], x[237], x[236], x[219], x[218], x[217]}), .y(y[104]));
  R2ind105 R2ind105_inst(.x({x[30], x[242], x[241], x[240], x[239], x[54], x[53], x[52], x[152], x[151], x[150], x[238], x[237], x[236], x[219], x[218], x[217]}), .y(y[105]));
  R2ind106 R2ind106_inst(.x({x[30], x[246], x[245], x[244], x[243], x[54], x[53], x[52], x[152], x[151], x[150], x[222], x[221], x[220], x[226], x[225], x[224]}), .y(y[106]));
  R2ind107 R2ind107_inst(.x({x[30], x[246], x[245], x[244], x[243], x[54], x[53], x[52], x[152], x[151], x[150], x[222], x[221], x[220], x[226], x[225], x[224]}), .y(y[107]));
  R2ind108 R2ind108_inst(.x({x[30], x[250], x[249], x[248], x[247], x[54], x[53], x[52], x[152], x[151], x[150], x[134], x[133], x[132], x[141], x[140], x[139]}), .y(y[108]));
  R2ind109 R2ind109_inst(.x({x[30], x[250], x[249], x[248], x[247], x[54], x[53], x[52], x[152], x[151], x[150], x[134], x[133], x[132], x[141], x[140], x[139]}), .y(y[109]));
  R2ind110 R2ind110_inst(.x({x[30], x[254], x[95], x[94], x[93], x[54], x[53], x[52], x[152], x[151], x[150], x[253], x[252], x[251], x[231], x[230], x[229]}), .y(y[110]));
  R2ind111 R2ind111_inst(.x({x[30], x[254], x[95], x[94], x[93], x[54], x[53], x[52], x[152], x[151], x[150], x[253], x[252], x[251], x[231], x[230], x[229]}), .y(y[111]));
  R2ind112 R2ind112_inst(.x({x[30], x[261], x[260], x[259], x[258], x[54], x[53], x[52], x[152], x[151], x[150], x[257], x[256], x[255], x[238], x[237], x[236]}), .y(y[112]));
  R2ind113 R2ind113_inst(.x({x[30], x[261], x[260], x[259], x[258], x[54], x[53], x[52], x[152], x[151], x[150], x[257], x[256], x[255], x[238], x[237], x[236]}), .y(y[113]));
  R2ind114 R2ind114_inst(.x({x[30], x[265], x[264], x[263], x[262], x[54], x[53], x[52], x[152], x[151], x[150], x[215], x[214], x[213], x[222], x[221], x[220]}), .y(y[114]));
  R2ind115 R2ind115_inst(.x({x[30], x[265], x[264], x[263], x[262], x[54], x[53], x[52], x[152], x[151], x[150], x[215], x[214], x[213], x[222], x[221], x[220]}), .y(y[115]));
  R2ind116 R2ind116_inst(.x({x[30], x[269], x[268], x[267], x[266], x[54], x[53], x[52], x[152], x[151], x[150], x[127], x[126], x[125], x[134], x[133], x[132]}), .y(y[116]));
  R2ind117 R2ind117_inst(.x({x[30], x[269], x[268], x[267], x[266], x[54], x[53], x[52], x[152], x[151], x[150], x[127], x[126], x[125], x[134], x[133], x[132]}), .y(y[117]));
  R2ind118 R2ind118_inst(.x({x[30], x[273], x[181], x[180], x[179], x[54], x[53], x[52], x[152], x[151], x[150], x[272], x[271], x[270], x[253], x[252], x[251]}), .y(y[118]));
  R2ind119 R2ind119_inst(.x({x[30], x[273], x[181], x[180], x[179], x[54], x[53], x[52], x[152], x[151], x[150], x[272], x[271], x[270], x[253], x[252], x[251]}), .y(y[119]));
  R2ind120 R2ind120_inst(.x({x[30], x[277], x[159], x[158], x[157], x[54], x[53], x[52], x[152], x[151], x[150], x[276], x[275], x[274], x[257], x[256], x[255]}), .y(y[120]));
  R2ind121 R2ind121_inst(.x({x[30], x[277], x[159], x[158], x[157], x[54], x[53], x[52], x[152], x[151], x[150], x[276], x[275], x[274], x[257], x[256], x[255]}), .y(y[121]));
  R2ind122 R2ind122_inst(.x({x[30], x[278], x[131], x[130], x[129], x[54], x[53], x[52], x[152], x[151], x[150], x[249], x[248], x[247], x[215], x[214], x[213]}), .y(y[122]));
  R2ind123 R2ind123_inst(.x({x[30], x[278], x[131], x[130], x[129], x[54], x[53], x[52], x[152], x[151], x[150], x[249], x[248], x[247], x[215], x[214], x[213]}), .y(y[123]));
  R2ind124 R2ind124_inst(.x({x[30], x[279], x[98], x[97], x[96], x[54], x[53], x[52], x[152], x[151], x[150], x[173], x[172], x[171], x[127], x[126], x[125]}), .y(y[124]));
  R2ind125 R2ind125_inst(.x({x[30], x[279], x[98], x[97], x[96], x[54], x[53], x[52], x[152], x[151], x[150], x[173], x[172], x[171], x[127], x[126], x[125]}), .y(y[125]));
  R2ind126 R2ind126_inst(.x({x[286], x[257], x[256], x[255], x[30], x[285], x[284], x[283], x[282], x[281], x[280], x[272], x[271], x[270], x[54], x[53], x[52]}), .y(y[126]));
  R2ind127 R2ind127_inst(.x({x[286], x[257], x[256], x[255], x[30], x[285], x[284], x[283], x[282], x[281], x[280], x[272], x[271], x[270], x[54], x[53], x[52]}), .y(y[127]));
  R2ind128 R2ind128_inst(.x({x[30], x[290], x[238], x[237], x[236], x[285], x[284], x[283], x[289], x[288], x[287], x[276], x[275], x[274], x[54], x[53], x[52]}), .y(y[128]));
  R2ind129 R2ind129_inst(.x({x[30], x[290], x[238], x[237], x[236], x[285], x[284], x[283], x[289], x[288], x[287], x[276], x[275], x[274], x[54], x[53], x[52]}), .y(y[129]));
  R2ind130 R2ind130_inst(.x({x[30], x[291], x[219], x[218], x[217], x[285], x[284], x[283], x[245], x[244], x[243], x[249], x[248], x[247], x[54], x[53], x[52]}), .y(y[130]));
  R2ind131 R2ind131_inst(.x({x[30], x[291], x[219], x[218], x[217], x[285], x[284], x[283], x[245], x[244], x[243], x[249], x[248], x[247], x[54], x[53], x[52]}), .y(y[131]));
  R2ind132 R2ind132_inst(.x({x[30], x[292], x[203], x[202], x[201], x[285], x[284], x[283], x[169], x[168], x[167], x[173], x[172], x[171], x[54], x[53], x[52]}), .y(y[132]));
  R2ind133 R2ind133_inst(.x({x[30], x[292], x[203], x[202], x[201], x[285], x[284], x[283], x[169], x[168], x[167], x[173], x[172], x[171], x[54], x[53], x[52]}), .y(y[133]));
  R2ind134 R2ind134_inst(.x({x[305], x[304], x[303], x[302], x[30], x[301], x[300], x[299], x[298], x[297], x[296], x[118], x[117], x[116], x[295], x[294], x[293]}), .y(y[134]));
  R2ind135 R2ind135_inst(.x({x[305], x[304], x[303], x[302], x[30], x[301], x[300], x[299], x[298], x[297], x[296], x[118], x[117], x[116], x[295], x[294], x[293]}), .y(y[135]));
  R2ind136 R2ind136_inst(.x({x[312], x[311], x[310], x[309], x[30], x[301], x[300], x[299], x[308], x[307], x[306], x[105], x[104], x[103], x[295], x[294], x[293]}), .y(y[136]));
  R2ind137 R2ind137_inst(.x({x[312], x[311], x[310], x[309], x[30], x[301], x[300], x[299], x[308], x[307], x[306], x[105], x[104], x[103], x[295], x[294], x[293]}), .y(y[137]));
  R2ind138 R2ind138_inst(.x({x[319], x[318], x[317], x[316], x[30], x[301], x[300], x[299], x[315], x[314], x[313], x[92], x[91], x[90], x[295], x[294], x[293]}), .y(y[138]));
  R2ind139 R2ind139_inst(.x({x[319], x[318], x[317], x[316], x[30], x[301], x[300], x[299], x[315], x[314], x[313], x[92], x[91], x[90], x[295], x[294], x[293]}), .y(y[139]));
  R2ind140 R2ind140_inst(.x({x[323], x[298], x[297], x[296], x[30], x[301], x[300], x[299], x[322], x[321], x[320], x[67], x[66], x[65], x[295], x[294], x[293]}), .y(y[140]));
  R2ind141 R2ind141_inst(.x({x[323], x[298], x[297], x[296], x[30], x[301], x[300], x[299], x[322], x[321], x[320], x[67], x[66], x[65], x[295], x[294], x[293]}), .y(y[141]));
  R2ind142 R2ind142_inst(.x({x[333], x[332], x[331], x[330], x[30], x[329], x[328], x[327], x[326], x[325], x[324], x[298], x[297], x[296], x[295], x[294], x[293]}), .y(y[142]));
  R2ind143 R2ind143_inst(.x({x[333], x[332], x[331], x[330], x[30], x[329], x[328], x[327], x[326], x[325], x[324], x[298], x[297], x[296], x[295], x[294], x[293]}), .y(y[143]));
  R2ind144 R2ind144_inst(.x({x[337], x[336], x[335], x[334], x[30], x[329], x[328], x[327], x[304], x[303], x[302], x[308], x[307], x[306], x[295], x[294], x[293]}), .y(y[144]));
  R2ind145 R2ind145_inst(.x({x[337], x[336], x[335], x[334], x[30], x[329], x[328], x[327], x[304], x[303], x[302], x[308], x[307], x[306], x[295], x[294], x[293]}), .y(y[145]));
  R2ind146 R2ind146_inst(.x({x[341], x[340], x[339], x[338], x[30], x[329], x[328], x[327], x[311], x[310], x[309], x[315], x[314], x[313], x[295], x[294], x[293]}), .y(y[146]));
  R2ind147 R2ind147_inst(.x({x[341], x[340], x[339], x[338], x[30], x[329], x[328], x[327], x[311], x[310], x[309], x[315], x[314], x[313], x[295], x[294], x[293]}), .y(y[147]));
  R2ind148 R2ind148_inst(.x({x[342], x[326], x[325], x[324], x[30], x[329], x[328], x[327], x[318], x[317], x[316], x[322], x[321], x[320], x[295], x[294], x[293]}), .y(y[148]));
  R2ind149 R2ind149_inst(.x({x[342], x[326], x[325], x[324], x[30], x[329], x[328], x[327], x[318], x[317], x[316], x[322], x[321], x[320], x[295], x[294], x[293]}), .y(y[149]));
  R2ind150 R2ind150_inst(.x({x[349], x[348], x[347], x[346], x[30], x[295], x[294], x[293], x[301], x[300], x[299], x[345], x[344], x[343], x[326], x[325], x[324]}), .y(y[150]));
  R2ind151 R2ind151_inst(.x({x[349], x[348], x[347], x[346], x[30], x[295], x[294], x[293], x[301], x[300], x[299], x[345], x[344], x[343], x[326], x[325], x[324]}), .y(y[151]));
  R2ind152 R2ind152_inst(.x({x[353], x[352], x[351], x[350], x[30], x[295], x[294], x[293], x[301], x[300], x[299], x[332], x[331], x[330], x[304], x[303], x[302]}), .y(y[152]));
  R2ind153 R2ind153_inst(.x({x[353], x[352], x[351], x[350], x[30], x[295], x[294], x[293], x[301], x[300], x[299], x[332], x[331], x[330], x[304], x[303], x[302]}), .y(y[153]));
  R2ind154 R2ind154_inst(.x({x[357], x[356], x[355], x[354], x[30], x[295], x[294], x[293], x[301], x[300], x[299], x[336], x[335], x[334], x[311], x[310], x[309]}), .y(y[154]));
  R2ind155 R2ind155_inst(.x({x[357], x[356], x[355], x[354], x[30], x[295], x[294], x[293], x[301], x[300], x[299], x[336], x[335], x[334], x[311], x[310], x[309]}), .y(y[155]));
  R2ind156 R2ind156_inst(.x({x[358], x[345], x[344], x[343], x[30], x[295], x[294], x[293], x[301], x[300], x[299], x[340], x[339], x[338], x[318], x[317], x[316]}), .y(y[156]));
  R2ind157 R2ind157_inst(.x({x[358], x[345], x[344], x[343], x[30], x[295], x[294], x[293], x[301], x[300], x[299], x[340], x[339], x[338], x[318], x[317], x[316]}), .y(y[157]));
  R2ind158 R2ind158_inst(.x({x[365], x[364], x[363], x[45], x[44], x[43], x[362], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[361], x[360], x[359], x[345], x[344], x[343]}), .y(y[158]));
  R2ind159 R2ind159_inst(.x({x[365], x[364], x[363], x[45], x[44], x[43], x[362], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[361], x[360], x[359], x[345], x[344], x[343]}), .y(y[159]));
  R2ind160 R2ind160_inst(.x({x[369], x[368], x[367], x[366], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[348], x[347], x[346], x[332], x[331], x[330]}), .y(y[160]));
  R2ind161 R2ind161_inst(.x({x[369], x[368], x[367], x[366], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[348], x[347], x[346], x[332], x[331], x[330]}), .y(y[161]));
  R2ind162 R2ind162_inst(.x({x[373], x[372], x[371], x[370], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[352], x[351], x[350], x[336], x[335], x[334]}), .y(y[162]));
  R2ind163 R2ind163_inst(.x({x[373], x[372], x[371], x[370], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[352], x[351], x[350], x[336], x[335], x[334]}), .y(y[163]));
  R2ind164 R2ind164_inst(.x({x[374], x[361], x[360], x[359], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[356], x[355], x[354], x[340], x[339], x[338]}), .y(y[164]));
  R2ind165 R2ind165_inst(.x({x[374], x[361], x[360], x[359], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[356], x[355], x[354], x[340], x[339], x[338]}), .y(y[165]));
  R2ind166 R2ind166_inst(.x({x[381], x[380], x[379], x[42], x[41], x[40], x[378], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[377], x[376], x[375], x[361], x[360], x[359]}), .y(y[166]));
  R2ind167 R2ind167_inst(.x({x[381], x[380], x[379], x[42], x[41], x[40], x[378], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[377], x[376], x[375], x[361], x[360], x[359]}), .y(y[167]));
  R2ind168 R2ind168_inst(.x({x[385], x[384], x[383], x[36], x[35], x[34], x[382], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[365], x[364], x[363], x[348], x[347], x[346]}), .y(y[168]));
  R2ind169 R2ind169_inst(.x({x[385], x[384], x[383], x[36], x[35], x[34], x[382], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[365], x[364], x[363], x[348], x[347], x[346]}), .y(y[169]));
  R2ind170 R2ind170_inst(.x({x[389], x[388], x[387], x[39], x[38], x[37], x[386], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[368], x[367], x[366], x[352], x[351], x[350]}), .y(y[170]));
  R2ind171 R2ind171_inst(.x({x[389], x[388], x[387], x[39], x[38], x[37], x[386], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[368], x[367], x[366], x[352], x[351], x[350]}), .y(y[171]));
  R2ind172 R2ind172_inst(.x({x[377], x[376], x[375], x[33], x[32], x[31], x[390], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[372], x[371], x[370], x[356], x[355], x[354]}), .y(y[172]));
  R2ind173 R2ind173_inst(.x({x[377], x[376], x[375], x[33], x[32], x[31], x[390], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[372], x[371], x[370], x[356], x[355], x[354]}), .y(y[173]));
  R2ind174 R2ind174_inst(.x({x[397], x[396], x[395], x[394], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[393], x[392], x[391], x[377], x[376], x[375]}), .y(y[174]));
  R2ind175 R2ind175_inst(.x({x[397], x[396], x[395], x[394], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[393], x[392], x[391], x[377], x[376], x[375]}), .y(y[175]));
  R2ind176 R2ind176_inst(.x({x[401], x[400], x[399], x[398], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[381], x[380], x[379], x[365], x[364], x[363]}), .y(y[176]));
  R2ind177 R2ind177_inst(.x({x[401], x[400], x[399], x[398], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[381], x[380], x[379], x[365], x[364], x[363]}), .y(y[177]));
  R2ind178 R2ind178_inst(.x({x[405], x[404], x[403], x[402], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[385], x[384], x[383], x[368], x[367], x[366]}), .y(y[178]));
  R2ind179 R2ind179_inst(.x({x[405], x[404], x[403], x[402], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[385], x[384], x[383], x[368], x[367], x[366]}), .y(y[179]));
  R2ind180 R2ind180_inst(.x({x[406], x[393], x[392], x[391], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[389], x[388], x[387], x[372], x[371], x[370]}), .y(y[180]));
  R2ind181 R2ind181_inst(.x({x[406], x[393], x[392], x[391], x[30], x[295], x[294], x[293], x[48], x[47], x[46], x[389], x[388], x[387], x[372], x[371], x[370]}), .y(y[181]));
  R2ind182 R2ind182_inst(.x({x[413], x[412], x[411], x[410], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[409], x[408], x[407], x[393], x[392], x[391]}), .y(y[182]));
  R2ind183 R2ind183_inst(.x({x[413], x[412], x[411], x[410], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[409], x[408], x[407], x[393], x[392], x[391]}), .y(y[183]));
  R2ind184 R2ind184_inst(.x({x[417], x[416], x[415], x[414], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[396], x[395], x[394], x[381], x[380], x[379]}), .y(y[184]));
  R2ind185 R2ind185_inst(.x({x[417], x[416], x[415], x[414], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[396], x[395], x[394], x[381], x[380], x[379]}), .y(y[185]));
  R2ind186 R2ind186_inst(.x({x[421], x[420], x[419], x[418], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[400], x[399], x[398], x[385], x[384], x[383]}), .y(y[186]));
  R2ind187 R2ind187_inst(.x({x[421], x[420], x[419], x[418], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[400], x[399], x[398], x[385], x[384], x[383]}), .y(y[187]));
  R2ind188 R2ind188_inst(.x({x[422], x[409], x[408], x[407], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[404], x[403], x[402], x[389], x[388], x[387]}), .y(y[188]));
  R2ind189 R2ind189_inst(.x({x[422], x[409], x[408], x[407], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[404], x[403], x[402], x[389], x[388], x[387]}), .y(y[189]));
  R2ind190 R2ind190_inst(.x({x[429], x[428], x[427], x[426], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[425], x[424], x[423], x[409], x[408], x[407]}), .y(y[190]));
  R2ind191 R2ind191_inst(.x({x[429], x[428], x[427], x[426], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[425], x[424], x[423], x[409], x[408], x[407]}), .y(y[191]));
  R2ind192 R2ind192_inst(.x({x[433], x[432], x[431], x[430], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[412], x[411], x[410], x[396], x[395], x[394]}), .y(y[192]));
  R2ind193 R2ind193_inst(.x({x[433], x[432], x[431], x[430], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[412], x[411], x[410], x[396], x[395], x[394]}), .y(y[193]));
  R2ind194 R2ind194_inst(.x({x[437], x[436], x[435], x[434], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[416], x[415], x[414], x[400], x[399], x[398]}), .y(y[194]));
  R2ind195 R2ind195_inst(.x({x[437], x[436], x[435], x[434], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[416], x[415], x[414], x[400], x[399], x[398]}), .y(y[195]));
  R2ind196 R2ind196_inst(.x({x[438], x[425], x[424], x[423], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[420], x[419], x[418], x[404], x[403], x[402]}), .y(y[196]));
  R2ind197 R2ind197_inst(.x({x[438], x[425], x[424], x[423], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[420], x[419], x[418], x[404], x[403], x[402]}), .y(y[197]));
  R2ind198 R2ind198_inst(.x({x[445], x[444], x[443], x[442], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[441], x[440], x[439], x[425], x[424], x[423]}), .y(y[198]));
  R2ind199 R2ind199_inst(.x({x[445], x[444], x[443], x[442], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[441], x[440], x[439], x[425], x[424], x[423]}), .y(y[199]));
  R2ind200 R2ind200_inst(.x({x[449], x[448], x[447], x[446], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[428], x[427], x[426], x[412], x[411], x[410]}), .y(y[200]));
  R2ind201 R2ind201_inst(.x({x[449], x[448], x[447], x[446], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[428], x[427], x[426], x[412], x[411], x[410]}), .y(y[201]));
  R2ind202 R2ind202_inst(.x({x[453], x[452], x[451], x[450], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[432], x[431], x[430], x[416], x[415], x[414]}), .y(y[202]));
  R2ind203 R2ind203_inst(.x({x[453], x[452], x[451], x[450], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[432], x[431], x[430], x[416], x[415], x[414]}), .y(y[203]));
  R2ind204 R2ind204_inst(.x({x[454], x[441], x[440], x[439], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[436], x[435], x[434], x[420], x[419], x[418]}), .y(y[204]));
  R2ind205 R2ind205_inst(.x({x[454], x[441], x[440], x[439], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[436], x[435], x[434], x[420], x[419], x[418]}), .y(y[205]));
  R2ind206 R2ind206_inst(.x({x[461], x[460], x[459], x[458], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[457], x[456], x[455], x[441], x[440], x[439]}), .y(y[206]));
  R2ind207 R2ind207_inst(.x({x[461], x[460], x[459], x[458], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[457], x[456], x[455], x[441], x[440], x[439]}), .y(y[207]));
  R2ind208 R2ind208_inst(.x({x[465], x[464], x[463], x[462], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[444], x[443], x[442], x[428], x[427], x[426]}), .y(y[208]));
  R2ind209 R2ind209_inst(.x({x[465], x[464], x[463], x[462], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[444], x[443], x[442], x[428], x[427], x[426]}), .y(y[209]));
  R2ind210 R2ind210_inst(.x({x[469], x[468], x[467], x[466], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[448], x[447], x[446], x[432], x[431], x[430]}), .y(y[210]));
  R2ind211 R2ind211_inst(.x({x[469], x[468], x[467], x[466], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[448], x[447], x[446], x[432], x[431], x[430]}), .y(y[211]));
  R2ind212 R2ind212_inst(.x({x[470], x[457], x[456], x[455], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[452], x[451], x[450], x[436], x[435], x[434]}), .y(y[212]));
  R2ind213 R2ind213_inst(.x({x[470], x[457], x[456], x[455], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[452], x[451], x[450], x[436], x[435], x[434]}), .y(y[213]));
  R2ind214 R2ind214_inst(.x({x[477], x[476], x[475], x[474], x[30], x[285], x[284], x[283], x[473], x[472], x[471], x[282], x[281], x[280], x[54], x[53], x[52]}), .y(y[214]));
  R2ind215 R2ind215_inst(.x({x[477], x[476], x[475], x[474], x[30], x[285], x[284], x[283], x[473], x[472], x[471], x[282], x[281], x[280], x[54], x[53], x[52]}), .y(y[215]));
  R2ind216 R2ind216_inst(.x({x[30], x[481], x[285], x[284], x[283], x[480], x[479], x[478], x[289], x[288], x[287], x[54], x[53], x[52]}), .y(y[216]));
  R2ind217 R2ind217_inst(.x({x[30], x[481], x[285], x[284], x[283], x[480], x[479], x[478], x[289], x[288], x[287], x[54], x[53], x[52]}), .y(y[217]));
  R2ind218 R2ind218_inst(.x({x[30], x[482], x[289], x[288], x[287], x[285], x[284], x[283], x[241], x[240], x[239], x[245], x[244], x[243], x[54], x[53], x[52]}), .y(y[218]));
  R2ind219 R2ind219_inst(.x({x[30], x[482], x[289], x[288], x[287], x[285], x[284], x[283], x[241], x[240], x[239], x[245], x[244], x[243], x[54], x[53], x[52]}), .y(y[219]));
  R2ind220 R2ind220_inst(.x({x[483], x[276], x[275], x[274], x[30], x[285], x[284], x[283], x[162], x[161], x[160], x[169], x[168], x[167], x[54], x[53], x[52]}), .y(y[220]));
  R2ind221 R2ind221_inst(.x({x[483], x[276], x[275], x[274], x[30], x[285], x[284], x[283], x[162], x[161], x[160], x[169], x[168], x[167], x[54], x[53], x[52]}), .y(y[221]));
  R2ind222 R2ind222_inst(.x({x[30], x[487], x[108], x[107], x[106], x[285], x[284], x[283], x[486], x[485], x[484], x[473], x[472], x[471], x[54], x[53], x[52]}), .y(y[222]));
  R2ind223 R2ind223_inst(.x({x[30], x[487], x[108], x[107], x[106], x[285], x[284], x[283], x[486], x[485], x[484], x[473], x[472], x[471], x[54], x[53], x[52]}), .y(y[223]));
  R2ind224 R2ind224_inst(.x({x[30], x[491], x[490], x[489], x[488], x[285], x[284], x[283], x[476], x[475], x[474], x[480], x[479], x[478], x[54], x[53], x[52]}), .y(y[224]));
  R2ind225 R2ind225_inst(.x({x[30], x[491], x[490], x[489], x[488], x[285], x[284], x[283], x[476], x[475], x[474], x[480], x[479], x[478], x[54], x[53], x[52]}), .y(y[225]));
  R2ind226 R2ind226_inst(.x({x[495], x[494], x[493], x[492], x[30], x[285], x[284], x[283], x[234], x[233], x[232], x[241], x[240], x[239], x[54], x[53], x[52]}), .y(y[226]));
  R2ind227 R2ind227_inst(.x({x[495], x[494], x[493], x[492], x[30], x[285], x[284], x[283], x[234], x[233], x[232], x[241], x[240], x[239], x[54], x[53], x[52]}), .y(y[227]));
  R2ind228 R2ind228_inst(.x({x[499], x[498], x[497], x[496], x[30], x[285], x[284], x[283], x[155], x[154], x[153], x[162], x[161], x[160], x[54], x[53], x[52]}), .y(y[228]));
  R2ind229 R2ind229_inst(.x({x[499], x[498], x[497], x[496], x[30], x[285], x[284], x[283], x[155], x[154], x[153], x[162], x[161], x[160], x[54], x[53], x[52]}), .y(y[229]));
  R2ind230 R2ind230_inst(.x({x[503], x[177], x[176], x[175], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[502], x[501], x[500], x[486], x[485], x[484]}), .y(y[230]));
  R2ind231 R2ind231_inst(.x({x[503], x[177], x[176], x[175], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[502], x[501], x[500], x[486], x[485], x[484]}), .y(y[231]));
  R2ind232 R2ind232_inst(.x({x[30], x[504], x[149], x[148], x[147], x[54], x[53], x[52], x[285], x[284], x[283], x[498], x[497], x[496], x[476], x[475], x[474]}), .y(y[232]));
  R2ind233 R2ind233_inst(.x({x[30], x[504], x[149], x[148], x[147], x[54], x[53], x[52], x[285], x[284], x[283], x[498], x[497], x[496], x[476], x[475], x[474]}), .y(y[233]));
  R2ind234 R2ind234_inst(.x({x[30], x[505], x[124], x[123], x[122], x[54], x[53], x[52], x[285], x[284], x[283], x[268], x[267], x[266], x[234], x[233], x[232]}), .y(y[234]));
  R2ind235 R2ind235_inst(.x({x[30], x[505], x[124], x[123], x[122], x[54], x[53], x[52], x[285], x[284], x[283], x[268], x[267], x[266], x[234], x[233], x[232]}), .y(y[235]));
  R2ind236 R2ind236_inst(.x({x[30], x[506], x[111], x[110], x[109], x[54], x[53], x[52], x[285], x[284], x[283], x[195], x[194], x[193], x[155], x[154], x[153]}), .y(y[236]));
  R2ind237 R2ind237_inst(.x({x[30], x[506], x[111], x[110], x[109], x[54], x[53], x[52], x[285], x[284], x[283], x[195], x[194], x[193], x[155], x[154], x[153]}), .y(y[237]));
  R2ind238 R2ind238_inst(.x({x[510], x[253], x[252], x[251], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[509], x[508], x[507], x[502], x[501], x[500]}), .y(y[238]));
  R2ind239 R2ind239_inst(.x({x[510], x[253], x[252], x[251], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[509], x[508], x[507], x[502], x[501], x[500]}), .y(y[239]));
  R2ind240 R2ind240_inst(.x({x[511], x[231], x[230], x[229], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[494], x[493], x[492], x[498], x[497], x[496]}), .y(y[240]));
  R2ind241 R2ind241_inst(.x({x[511], x[231], x[230], x[229], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[494], x[493], x[492], x[498], x[497], x[496]}), .y(y[241]));
  R2ind242 R2ind242_inst(.x({x[512], x[212], x[211], x[210], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[264], x[263], x[262], x[268], x[267], x[266]}), .y(y[242]));
  R2ind243 R2ind243_inst(.x({x[512], x[212], x[211], x[210], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[264], x[263], x[262], x[268], x[267], x[266]}), .y(y[243]));
  R2ind244 R2ind244_inst(.x({x[513], x[199], x[198], x[197], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[191], x[190], x[189], x[195], x[194], x[193]}), .y(y[244]));
  R2ind245 R2ind245_inst(.x({x[513], x[199], x[198], x[197], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[191], x[190], x[189], x[195], x[194], x[193]}), .y(y[245]));
  R2ind246 R2ind246_inst(.x({x[517], x[486], x[485], x[484], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[516], x[515], x[514], x[509], x[508], x[507]}), .y(y[246]));
  R2ind247 R2ind247_inst(.x({x[517], x[486], x[485], x[484], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[516], x[515], x[514], x[509], x[508], x[507]}), .y(y[247]));
  R2ind248 R2ind248_inst(.x({x[518], x[473], x[472], x[471], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[490], x[489], x[488], x[494], x[493], x[492]}), .y(y[248]));
  R2ind249 R2ind249_inst(.x({x[518], x[473], x[472], x[471], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[490], x[489], x[488], x[494], x[493], x[492]}), .y(y[249]));
  R2ind250 R2ind250_inst(.x({x[519], x[282], x[281], x[280], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[260], x[259], x[258], x[264], x[263], x[262]}), .y(y[250]));
  R2ind251 R2ind251_inst(.x({x[519], x[282], x[281], x[280], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[260], x[259], x[258], x[264], x[263], x[262]}), .y(y[251]));
  R2ind252 R2ind252_inst(.x({x[520], x[272], x[271], x[270], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[184], x[183], x[182], x[191], x[190], x[189]}), .y(y[252]));
  R2ind253 R2ind253_inst(.x({x[520], x[272], x[271], x[270], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[184], x[183], x[182], x[191], x[190], x[189]}), .y(y[253]));
  R2ind254 R2ind254_inst(.x({x[30], x[521], x[54], x[53], x[52], x[285], x[284], x[283], x[121], x[120], x[119], x[516], x[515], x[514]}), .y(y[254]));
  R2ind255 R2ind255_inst(.x({x[30], x[521], x[54], x[53], x[52], x[285], x[284], x[283], x[121], x[120], x[119], x[516], x[515], x[514]}), .y(y[255]));
  R2ind256 R2ind256_inst(.x({x[522], x[516], x[515], x[514], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[108], x[107], x[106], x[490], x[489], x[488]}), .y(y[256]));
  R2ind257 R2ind257_inst(.x({x[522], x[516], x[515], x[514], x[30], x[54], x[53], x[52], x[285], x[284], x[283], x[108], x[107], x[106], x[490], x[489], x[488]}), .y(y[257]));
  R2ind258 R2ind258_inst(.x({x[30], x[523], x[509], x[508], x[507], x[54], x[53], x[52], x[285], x[284], x[283], x[95], x[94], x[93], x[260], x[259], x[258]}), .y(y[258]));
  R2ind259 R2ind259_inst(.x({x[30], x[523], x[509], x[508], x[507], x[54], x[53], x[52], x[285], x[284], x[283], x[95], x[94], x[93], x[260], x[259], x[258]}), .y(y[259]));
  R2ind260 R2ind260_inst(.x({x[30], x[524], x[502], x[501], x[500], x[54], x[53], x[52], x[285], x[284], x[283], x[70], x[69], x[68], x[184], x[183], x[182]}), .y(y[260]));
  R2ind261 R2ind261_inst(.x({x[30], x[524], x[502], x[501], x[500], x[54], x[53], x[52], x[285], x[284], x[283], x[70], x[69], x[68], x[184], x[183], x[182]}), .y(y[261]));
  R2ind262 R2ind262_inst(.x({x[531], x[530], x[529], x[528], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[527], x[526], x[525], x[457], x[456], x[455]}), .y(y[262]));
  R2ind263 R2ind263_inst(.x({x[531], x[530], x[529], x[528], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[527], x[526], x[525], x[457], x[456], x[455]}), .y(y[263]));
  R2ind264 R2ind264_inst(.x({x[535], x[534], x[533], x[532], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[460], x[459], x[458], x[444], x[443], x[442]}), .y(y[264]));
  R2ind265 R2ind265_inst(.x({x[535], x[534], x[533], x[532], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[460], x[459], x[458], x[444], x[443], x[442]}), .y(y[265]));
  R2ind266 R2ind266_inst(.x({x[539], x[538], x[537], x[536], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[464], x[463], x[462], x[448], x[447], x[446]}), .y(y[266]));
  R2ind267 R2ind267_inst(.x({x[539], x[538], x[537], x[536], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[464], x[463], x[462], x[448], x[447], x[446]}), .y(y[267]));
  R2ind268 R2ind268_inst(.x({x[540], x[527], x[526], x[525], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[468], x[467], x[466], x[452], x[451], x[450]}), .y(y[268]));
  R2ind269 R2ind269_inst(.x({x[540], x[527], x[526], x[525], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[468], x[467], x[466], x[452], x[451], x[450]}), .y(y[269]));
  R2ind270 R2ind270_inst(.x({x[547], x[546], x[545], x[544], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[543], x[542], x[541], x[527], x[526], x[525]}), .y(y[270]));
  R2ind271 R2ind271_inst(.x({x[547], x[546], x[545], x[544], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[543], x[542], x[541], x[527], x[526], x[525]}), .y(y[271]));
  R2ind272 R2ind272_inst(.x({x[551], x[550], x[549], x[548], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[530], x[529], x[528], x[460], x[459], x[458]}), .y(y[272]));
  R2ind273 R2ind273_inst(.x({x[551], x[550], x[549], x[548], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[530], x[529], x[528], x[460], x[459], x[458]}), .y(y[273]));
  R2ind274 R2ind274_inst(.x({x[555], x[554], x[553], x[552], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[534], x[533], x[532], x[464], x[463], x[462]}), .y(y[274]));
  R2ind275 R2ind275_inst(.x({x[555], x[554], x[553], x[552], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[534], x[533], x[532], x[464], x[463], x[462]}), .y(y[275]));
  R2ind276 R2ind276_inst(.x({x[556], x[543], x[542], x[541], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[538], x[537], x[536], x[468], x[467], x[466]}), .y(y[276]));
  R2ind277 R2ind277_inst(.x({x[556], x[543], x[542], x[541], x[30], x[295], x[294], x[293], x[329], x[328], x[327], x[538], x[537], x[536], x[468], x[467], x[466]}), .y(y[277]));
  R2ind278 R2ind278_inst(.x({x[566], x[565], x[564], x[563], x[30], x[329], x[328], x[327], x[562], x[561], x[560], x[543], x[542], x[541], x[559], x[558], x[557]}), .y(y[278]));
  R2ind279 R2ind279_inst(.x({x[566], x[565], x[564], x[563], x[30], x[329], x[328], x[327], x[562], x[561], x[560], x[543], x[542], x[541], x[559], x[558], x[557]}), .y(y[279]));
  R2ind280 R2ind280_inst(.x({x[570], x[569], x[568], x[567], x[30], x[329], x[328], x[327], x[546], x[545], x[544], x[530], x[529], x[528], x[559], x[558], x[557]}), .y(y[280]));
  R2ind281 R2ind281_inst(.x({x[570], x[569], x[568], x[567], x[30], x[329], x[328], x[327], x[546], x[545], x[544], x[530], x[529], x[528], x[559], x[558], x[557]}), .y(y[281]));
  R2ind282 R2ind282_inst(.x({x[574], x[573], x[572], x[571], x[30], x[329], x[328], x[327], x[550], x[549], x[548], x[534], x[533], x[532], x[559], x[558], x[557]}), .y(y[282]));
  R2ind283 R2ind283_inst(.x({x[574], x[573], x[572], x[571], x[30], x[329], x[328], x[327], x[550], x[549], x[548], x[534], x[533], x[532], x[559], x[558], x[557]}), .y(y[283]));
  R2ind284 R2ind284_inst(.x({x[575], x[562], x[561], x[560], x[30], x[329], x[328], x[327], x[554], x[553], x[552], x[538], x[537], x[536], x[559], x[558], x[557]}), .y(y[284]));
  R2ind285 R2ind285_inst(.x({x[575], x[562], x[561], x[560], x[30], x[329], x[328], x[327], x[554], x[553], x[552], x[538], x[537], x[536], x[559], x[558], x[557]}), .y(y[285]));
  R2ind286 R2ind286_inst(.x({x[582], x[581], x[580], x[579], x[30], x[301], x[300], x[299], x[578], x[577], x[576], x[562], x[561], x[560], x[559], x[558], x[557]}), .y(y[286]));
  R2ind287 R2ind287_inst(.x({x[582], x[581], x[580], x[579], x[30], x[301], x[300], x[299], x[578], x[577], x[576], x[562], x[561], x[560], x[559], x[558], x[557]}), .y(y[287]));
  R2ind288 R2ind288_inst(.x({x[586], x[585], x[584], x[583], x[30], x[301], x[300], x[299], x[565], x[564], x[563], x[546], x[545], x[544], x[559], x[558], x[557]}), .y(y[288]));
  R2ind289 R2ind289_inst(.x({x[586], x[585], x[584], x[583], x[30], x[301], x[300], x[299], x[565], x[564], x[563], x[546], x[545], x[544], x[559], x[558], x[557]}), .y(y[289]));
  R2ind290 R2ind290_inst(.x({x[590], x[589], x[588], x[587], x[30], x[301], x[300], x[299], x[569], x[568], x[567], x[550], x[549], x[548], x[559], x[558], x[557]}), .y(y[290]));
  R2ind291 R2ind291_inst(.x({x[590], x[589], x[588], x[587], x[30], x[301], x[300], x[299], x[569], x[568], x[567], x[550], x[549], x[548], x[559], x[558], x[557]}), .y(y[291]));
  R2ind292 R2ind292_inst(.x({x[591], x[578], x[577], x[576], x[30], x[301], x[300], x[299], x[573], x[572], x[571], x[554], x[553], x[552], x[559], x[558], x[557]}), .y(y[292]));
  R2ind293 R2ind293_inst(.x({x[591], x[578], x[577], x[576], x[30], x[301], x[300], x[299], x[573], x[572], x[571], x[554], x[553], x[552], x[559], x[558], x[557]}), .y(y[293]));
  R2ind294 R2ind294_inst(.x({x[598], x[597], x[596], x[595], x[30], x[301], x[300], x[299], x[594], x[593], x[592], x[578], x[577], x[576], x[559], x[558], x[557]}), .y(y[294]));
  R2ind295 R2ind295_inst(.x({x[598], x[597], x[596], x[595], x[30], x[301], x[300], x[299], x[594], x[593], x[592], x[578], x[577], x[576], x[559], x[558], x[557]}), .y(y[295]));
  R2ind296 R2ind296_inst(.x({x[602], x[601], x[600], x[599], x[30], x[301], x[300], x[299], x[581], x[580], x[579], x[565], x[564], x[563], x[559], x[558], x[557]}), .y(y[296]));
  R2ind297 R2ind297_inst(.x({x[602], x[601], x[600], x[599], x[30], x[301], x[300], x[299], x[581], x[580], x[579], x[565], x[564], x[563], x[559], x[558], x[557]}), .y(y[297]));
  R2ind298 R2ind298_inst(.x({x[606], x[605], x[604], x[603], x[30], x[301], x[300], x[299], x[585], x[584], x[583], x[569], x[568], x[567], x[559], x[558], x[557]}), .y(y[298]));
  R2ind299 R2ind299_inst(.x({x[606], x[605], x[604], x[603], x[30], x[301], x[300], x[299], x[585], x[584], x[583], x[569], x[568], x[567], x[559], x[558], x[557]}), .y(y[299]));
  R2ind300 R2ind300_inst(.x({x[607], x[594], x[593], x[592], x[30], x[301], x[300], x[299], x[589], x[588], x[587], x[573], x[572], x[571], x[559], x[558], x[557]}), .y(y[300]));
  R2ind301 R2ind301_inst(.x({x[607], x[594], x[593], x[592], x[30], x[301], x[300], x[299], x[589], x[588], x[587], x[573], x[572], x[571], x[559], x[558], x[557]}), .y(y[301]));
  R2ind302 R2ind302_inst(.x({x[614], x[613], x[612], x[611], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[610], x[609], x[608], x[594], x[593], x[592]}), .y(y[302]));
  R2ind303 R2ind303_inst(.x({x[614], x[613], x[612], x[611], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[610], x[609], x[608], x[594], x[593], x[592]}), .y(y[303]));
  R2ind304 R2ind304_inst(.x({x[618], x[617], x[616], x[615], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[597], x[596], x[595], x[581], x[580], x[579]}), .y(y[304]));
  R2ind305 R2ind305_inst(.x({x[618], x[617], x[616], x[615], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[597], x[596], x[595], x[581], x[580], x[579]}), .y(y[305]));
  R2ind306 R2ind306_inst(.x({x[622], x[621], x[620], x[619], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[601], x[600], x[599], x[585], x[584], x[583]}), .y(y[306]));
  R2ind307 R2ind307_inst(.x({x[622], x[621], x[620], x[619], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[601], x[600], x[599], x[585], x[584], x[583]}), .y(y[307]));
  R2ind308 R2ind308_inst(.x({x[623], x[610], x[609], x[608], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[605], x[604], x[603], x[589], x[588], x[587]}), .y(y[308]));
  R2ind309 R2ind309_inst(.x({x[623], x[610], x[609], x[608], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[605], x[604], x[603], x[589], x[588], x[587]}), .y(y[309]));
  R2ind310 R2ind310_inst(.x({x[630], x[629], x[628], x[627], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[626], x[625], x[624], x[610], x[609], x[608]}), .y(y[310]));
  R2ind311 R2ind311_inst(.x({x[630], x[629], x[628], x[627], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[626], x[625], x[624], x[610], x[609], x[608]}), .y(y[311]));
  R2ind312 R2ind312_inst(.x({x[634], x[633], x[632], x[631], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[613], x[612], x[611], x[597], x[596], x[595]}), .y(y[312]));
  R2ind313 R2ind313_inst(.x({x[634], x[633], x[632], x[631], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[613], x[612], x[611], x[597], x[596], x[595]}), .y(y[313]));
  R2ind314 R2ind314_inst(.x({x[638], x[637], x[636], x[635], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[617], x[616], x[615], x[601], x[600], x[599]}), .y(y[314]));
  R2ind315 R2ind315_inst(.x({x[638], x[637], x[636], x[635], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[617], x[616], x[615], x[601], x[600], x[599]}), .y(y[315]));
  R2ind316 R2ind316_inst(.x({x[639], x[626], x[625], x[624], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[621], x[620], x[619], x[605], x[604], x[603]}), .y(y[316]));
  R2ind317 R2ind317_inst(.x({x[639], x[626], x[625], x[624], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[621], x[620], x[619], x[605], x[604], x[603]}), .y(y[317]));
  R2ind318 R2ind318_inst(.x({x[646], x[645], x[644], x[643], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[642], x[641], x[640], x[626], x[625], x[624]}), .y(y[318]));
  R2ind319 R2ind319_inst(.x({x[646], x[645], x[644], x[643], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[642], x[641], x[640], x[626], x[625], x[624]}), .y(y[319]));
  R2ind320 R2ind320_inst(.x({x[650], x[649], x[648], x[647], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[629], x[628], x[627], x[613], x[612], x[611]}), .y(y[320]));
  R2ind321 R2ind321_inst(.x({x[650], x[649], x[648], x[647], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[629], x[628], x[627], x[613], x[612], x[611]}), .y(y[321]));
  R2ind322 R2ind322_inst(.x({x[654], x[653], x[652], x[651], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[633], x[632], x[631], x[617], x[616], x[615]}), .y(y[322]));
  R2ind323 R2ind323_inst(.x({x[654], x[653], x[652], x[651], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[633], x[632], x[631], x[617], x[616], x[615]}), .y(y[323]));
  R2ind324 R2ind324_inst(.x({x[655], x[642], x[641], x[640], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[637], x[636], x[635], x[621], x[620], x[619]}), .y(y[324]));
  R2ind325 R2ind325_inst(.x({x[655], x[642], x[641], x[640], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[637], x[636], x[635], x[621], x[620], x[619]}), .y(y[325]));
  R2ind326 R2ind326_inst(.x({x[659], x[105], x[104], x[103], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[658], x[657], x[656], x[642], x[641], x[640]}), .y(y[326]));
  R2ind327 R2ind327_inst(.x({x[659], x[105], x[104], x[103], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[658], x[657], x[656], x[642], x[641], x[640]}), .y(y[327]));
  R2ind328 R2ind328_inst(.x({x[660], x[92], x[91], x[90], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[645], x[644], x[643], x[629], x[628], x[627]}), .y(y[328]));
  R2ind329 R2ind329_inst(.x({x[660], x[92], x[91], x[90], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[645], x[644], x[643], x[629], x[628], x[627]}), .y(y[329]));
  R2ind330 R2ind330_inst(.x({x[661], x[67], x[66], x[65], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[649], x[648], x[647], x[633], x[632], x[631]}), .y(y[330]));
  R2ind331 R2ind331_inst(.x({x[661], x[67], x[66], x[65], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[649], x[648], x[647], x[633], x[632], x[631]}), .y(y[331]));
  R2ind332 R2ind332_inst(.x({x[662], x[658], x[657], x[656], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[653], x[652], x[651], x[637], x[636], x[635]}), .y(y[332]));
  R2ind333 R2ind333_inst(.x({x[662], x[658], x[657], x[656], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[653], x[652], x[651], x[637], x[636], x[635]}), .y(y[333]));
  R2ind334 R2ind334_inst(.x({x[82], x[81], x[80], x[79], x[78], x[77], x[73], x[72], x[71], x[76], x[75], x[74], x[663], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[118], x[117], x[116], x[658], x[657], x[656]}), .y(y[334]));
  R2ind335 R2ind335_inst(.x({x[82], x[81], x[80], x[79], x[78], x[77], x[73], x[72], x[71], x[76], x[75], x[74], x[663], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[118], x[117], x[116], x[658], x[657], x[656]}), .y(y[335]));
  R2ind336 R2ind336_inst(.x({x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[82], x[81], x[80], x[664], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[105], x[104], x[103], x[645], x[644], x[643]}), .y(y[336]));
  R2ind337 R2ind337_inst(.x({x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[82], x[81], x[80], x[664], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[105], x[104], x[103], x[645], x[644], x[643]}), .y(y[337]));
  R2ind338 R2ind338_inst(.x({x[79], x[78], x[77], x[82], x[81], x[80], x[73], x[72], x[71], x[76], x[75], x[74], x[665], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[92], x[91], x[90], x[649], x[648], x[647]}), .y(y[338]));
  R2ind339 R2ind339_inst(.x({x[79], x[78], x[77], x[82], x[81], x[80], x[73], x[72], x[71], x[76], x[75], x[74], x[665], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[92], x[91], x[90], x[649], x[648], x[647]}), .y(y[339]));
  R2ind340 R2ind340_inst(.x({x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[666], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[67], x[66], x[65], x[653], x[652], x[651]}), .y(y[340]));
  R2ind341 R2ind341_inst(.x({x[82], x[81], x[80], x[79], x[78], x[77], x[76], x[75], x[74], x[73], x[72], x[71], x[666], x[30], x[559], x[558], x[557], x[301], x[300], x[299], x[67], x[66], x[65], x[653], x[652], x[651]}), .y(y[341]));
  R2ind342 R2ind342_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[70], x[69], x[68], x[67], x[66], x[65], x[118], x[117], x[116]}), .y(y[342]));
  R2ind343 R2ind343_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[70], x[69], x[68], x[67], x[66], x[65], x[118], x[117], x[116]}), .y(y[343]));
  R2ind344 R2ind344_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[95], x[94], x[93], x[92], x[91], x[90], x[322], x[321], x[320]}), .y(y[344]));
  R2ind345 R2ind345_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[95], x[94], x[93], x[92], x[91], x[90], x[322], x[321], x[320]}), .y(y[345]));
  R2ind346 R2ind346_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[108], x[107], x[106], x[105], x[104], x[103], x[315], x[314], x[313]}), .y(y[346]));
  R2ind347 R2ind347_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[108], x[107], x[106], x[105], x[104], x[103], x[315], x[314], x[313]}), .y(y[347]));
  R2ind348 R2ind348_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[121], x[120], x[119], x[118], x[117], x[116], x[308], x[307], x[306]}), .y(y[348]));
  R2ind349 R2ind349_inst(.x({x[14], x[13], x[12], x[11], x[10], x[9], x[17], x[16], x[15], x[8], x[7], x[6], x[121], x[120], x[119], x[118], x[117], x[116], x[308], x[307], x[306]}), .y(y[349]));
endmodule

