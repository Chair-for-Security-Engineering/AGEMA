/* modified netlist. Source: module sbox in file Designs/AESSbox/optBP2/AGEMA/sbox.v */
/* 8 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 9 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d2 (X_s0, clk, X_s1, X_s2, Fresh, Y_s0, Y_s1, Y_s2);
    input [7:0] X_s0 ;
    input clk ;
    input [7:0] X_s1 ;
    input [7:0] X_s2 ;
    input [101:0] Fresh ;
    output [7:0] Y_s0 ;
    output [7:0] Y_s1 ;
    output [7:0] Y_s2 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;
    wire signal_205 ;
    wire signal_206 ;
    wire signal_207 ;
    wire signal_208 ;
    wire signal_209 ;
    wire signal_210 ;
    wire signal_211 ;
    wire signal_212 ;
    wire signal_213 ;
    wire signal_214 ;
    wire signal_215 ;
    wire signal_216 ;
    wire signal_217 ;
    wire signal_218 ;
    wire signal_219 ;
    wire signal_220 ;
    wire signal_221 ;
    wire signal_222 ;
    wire signal_223 ;
    wire signal_224 ;
    wire signal_225 ;
    wire signal_226 ;
    wire signal_227 ;
    wire signal_228 ;
    wire signal_229 ;
    wire signal_230 ;
    wire signal_231 ;
    wire signal_232 ;
    wire signal_233 ;
    wire signal_234 ;
    wire signal_235 ;
    wire signal_236 ;
    wire signal_237 ;
    wire signal_238 ;
    wire signal_239 ;
    wire signal_240 ;
    wire signal_241 ;
    wire signal_242 ;
    wire signal_243 ;
    wire signal_244 ;
    wire signal_245 ;
    wire signal_246 ;
    wire signal_247 ;
    wire signal_248 ;
    wire signal_249 ;
    wire signal_250 ;
    wire signal_251 ;
    wire signal_252 ;
    wire signal_253 ;
    wire signal_254 ;
    wire signal_255 ;
    wire signal_256 ;
    wire signal_257 ;
    wire signal_258 ;
    wire signal_259 ;
    wire signal_260 ;
    wire signal_261 ;
    wire signal_262 ;
    wire signal_263 ;
    wire signal_264 ;
    wire signal_265 ;
    wire signal_266 ;
    wire signal_267 ;
    wire signal_268 ;
    wire signal_269 ;
    wire signal_270 ;
    wire signal_271 ;
    wire signal_272 ;
    wire signal_273 ;
    wire signal_274 ;
    wire signal_279 ;
    wire signal_280 ;
    wire signal_283 ;
    wire signal_284 ;
    wire signal_287 ;
    wire signal_288 ;
    wire signal_289 ;
    wire signal_290 ;
    wire signal_293 ;
    wire signal_294 ;
    wire signal_299 ;
    wire signal_300 ;
    wire signal_301 ;
    wire signal_302 ;
    wire signal_303 ;
    wire signal_304 ;
    wire signal_307 ;
    wire signal_308 ;
    wire signal_309 ;
    wire signal_310 ;
    wire signal_311 ;
    wire signal_312 ;
    wire signal_313 ;
    wire signal_314 ;
    wire signal_315 ;
    wire signal_316 ;
    wire signal_317 ;
    wire signal_318 ;
    wire signal_319 ;
    wire signal_320 ;
    wire signal_321 ;
    wire signal_322 ;
    wire signal_323 ;
    wire signal_324 ;
    wire signal_325 ;
    wire signal_326 ;
    wire signal_327 ;
    wire signal_328 ;
    wire signal_329 ;
    wire signal_330 ;
    wire signal_331 ;
    wire signal_332 ;
    wire signal_333 ;
    wire signal_334 ;
    wire signal_335 ;
    wire signal_336 ;
    wire signal_337 ;
    wire signal_338 ;
    wire signal_339 ;
    wire signal_340 ;
    wire signal_341 ;
    wire signal_342 ;
    wire signal_343 ;
    wire signal_344 ;
    wire signal_345 ;
    wire signal_346 ;
    wire signal_347 ;
    wire signal_348 ;
    wire signal_349 ;
    wire signal_350 ;
    wire signal_351 ;
    wire signal_352 ;
    wire signal_353 ;
    wire signal_354 ;
    wire signal_355 ;
    wire signal_356 ;
    wire signal_357 ;
    wire signal_358 ;
    wire signal_359 ;
    wire signal_360 ;
    wire signal_361 ;
    wire signal_362 ;
    wire signal_363 ;
    wire signal_364 ;
    wire signal_365 ;
    wire signal_366 ;
    wire signal_367 ;
    wire signal_368 ;
    wire signal_369 ;
    wire signal_370 ;
    wire signal_371 ;
    wire signal_372 ;
    wire signal_373 ;
    wire signal_374 ;
    wire signal_375 ;
    wire signal_376 ;
    wire signal_377 ;
    wire signal_378 ;
    wire signal_379 ;
    wire signal_380 ;
    wire signal_381 ;
    wire signal_382 ;
    wire signal_383 ;
    wire signal_384 ;
    wire signal_385 ;
    wire signal_386 ;
    wire signal_387 ;
    wire signal_388 ;
    wire signal_389 ;
    wire signal_390 ;
    wire signal_391 ;
    wire signal_392 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_415 ;
    wire signal_416 ;
    wire signal_417 ;
    wire signal_418 ;
    wire signal_419 ;
    wire signal_420 ;
    wire signal_421 ;
    wire signal_422 ;
    wire signal_423 ;
    wire signal_424 ;
    wire signal_425 ;
    wire signal_426 ;
    wire signal_427 ;
    wire signal_428 ;
    wire signal_429 ;
    wire signal_430 ;
    wire signal_431 ;
    wire signal_432 ;
    wire signal_433 ;
    wire signal_434 ;
    wire signal_435 ;
    wire signal_436 ;
    wire signal_437 ;
    wire signal_438 ;
    wire signal_439 ;
    wire signal_440 ;
    wire signal_441 ;
    wire signal_442 ;
    wire signal_443 ;
    wire signal_444 ;
    wire signal_445 ;
    wire signal_446 ;
    wire signal_447 ;
    wire signal_448 ;
    wire signal_449 ;
    wire signal_450 ;
    wire signal_451 ;
    wire signal_452 ;
    wire signal_453 ;
    wire signal_454 ;
    wire signal_455 ;
    wire signal_456 ;
    wire signal_457 ;
    wire signal_458 ;
    wire signal_459 ;
    wire signal_460 ;
    wire signal_461 ;
    wire signal_462 ;
    wire signal_463 ;
    wire signal_464 ;
    wire signal_465 ;
    wire signal_466 ;
    wire signal_467 ;
    wire signal_468 ;
    wire signal_469 ;
    wire signal_470 ;
    wire signal_471 ;
    wire signal_472 ;
    wire signal_473 ;
    wire signal_474 ;
    wire signal_475 ;
    wire signal_476 ;
    wire signal_477 ;
    wire signal_478 ;
    wire signal_479 ;
    wire signal_480 ;
    wire signal_481 ;
    wire signal_482 ;
    wire signal_483 ;
    wire signal_484 ;
    wire signal_485 ;
    wire signal_486 ;
    wire signal_487 ;
    wire signal_488 ;
    wire signal_489 ;
    wire signal_490 ;
    wire signal_491 ;
    wire signal_492 ;
    wire signal_493 ;
    wire signal_494 ;
    wire signal_495 ;
    wire signal_496 ;
    wire signal_497 ;
    wire signal_498 ;
    wire signal_499 ;
    wire signal_500 ;
    wire signal_501 ;
    wire signal_502 ;
    wire signal_503 ;
    wire signal_504 ;
    wire signal_505 ;
    wire signal_506 ;
    wire signal_507 ;
    wire signal_508 ;
    wire signal_509 ;
    wire signal_510 ;
    wire signal_511 ;
    wire signal_512 ;
    wire signal_513 ;
    wire signal_514 ;
    wire signal_515 ;
    wire signal_516 ;
    wire signal_517 ;
    wire signal_518 ;
    wire signal_519 ;
    wire signal_520 ;
    wire signal_521 ;
    wire signal_522 ;
    wire signal_523 ;
    wire signal_524 ;
    wire signal_525 ;
    wire signal_526 ;
    wire signal_527 ;
    wire signal_528 ;
    wire signal_529 ;
    wire signal_530 ;
    wire signal_531 ;
    wire signal_532 ;
    wire signal_533 ;
    wire signal_534 ;
    wire signal_535 ;
    wire signal_536 ;
    wire signal_537 ;
    wire signal_538 ;
    wire signal_539 ;
    wire signal_540 ;
    wire signal_541 ;
    wire signal_542 ;
    wire signal_543 ;
    wire signal_544 ;
    wire signal_545 ;
    wire signal_546 ;
    wire signal_547 ;
    wire signal_548 ;
    wire signal_549 ;
    wire signal_550 ;
    wire signal_551 ;
    wire signal_552 ;
    wire signal_553 ;
    wire signal_554 ;
    wire signal_673 ;
    wire signal_674 ;
    wire signal_675 ;
    wire signal_676 ;
    wire signal_677 ;
    wire signal_678 ;
    wire signal_679 ;
    wire signal_680 ;
    wire signal_681 ;
    wire signal_682 ;
    wire signal_683 ;
    wire signal_684 ;
    wire signal_685 ;
    wire signal_686 ;
    wire signal_687 ;
    wire signal_688 ;
    wire signal_689 ;
    wire signal_690 ;
    wire signal_691 ;
    wire signal_692 ;
    wire signal_693 ;
    wire signal_694 ;
    wire signal_695 ;
    wire signal_696 ;
    wire signal_697 ;
    wire signal_698 ;
    wire signal_699 ;
    wire signal_700 ;
    wire signal_701 ;
    wire signal_702 ;
    wire signal_703 ;
    wire signal_704 ;
    wire signal_705 ;
    wire signal_706 ;
    wire signal_707 ;
    wire signal_708 ;
    wire signal_709 ;
    wire signal_710 ;
    wire signal_711 ;
    wire signal_712 ;
    wire signal_713 ;
    wire signal_714 ;
    wire signal_715 ;
    wire signal_716 ;
    wire signal_717 ;
    wire signal_718 ;
    wire signal_719 ;
    wire signal_720 ;
    wire signal_721 ;
    wire signal_722 ;
    wire signal_723 ;
    wire signal_724 ;
    wire signal_725 ;
    wire signal_726 ;
    wire signal_727 ;
    wire signal_728 ;
    wire signal_729 ;
    wire signal_730 ;
    wire signal_731 ;
    wire signal_732 ;
    wire signal_733 ;
    wire signal_734 ;
    wire signal_735 ;
    wire signal_736 ;
    wire signal_737 ;
    wire signal_738 ;
    wire signal_739 ;
    wire signal_740 ;
    wire signal_741 ;
    wire signal_742 ;
    wire signal_743 ;
    wire signal_744 ;
    wire signal_745 ;
    wire signal_746 ;
    wire signal_747 ;
    wire signal_748 ;
    wire signal_749 ;
    wire signal_750 ;
    wire signal_751 ;
    wire signal_752 ;
    wire signal_753 ;
    wire signal_754 ;
    wire signal_755 ;
    wire signal_756 ;
    wire signal_757 ;
    wire signal_758 ;
    wire signal_759 ;
    wire signal_760 ;
    wire signal_761 ;
    wire signal_762 ;
    wire signal_763 ;
    wire signal_764 ;
    wire signal_765 ;
    wire signal_766 ;
    wire signal_767 ;
    wire signal_768 ;
    wire signal_769 ;
    wire signal_770 ;
    wire signal_771 ;
    wire signal_772 ;
    wire signal_773 ;
    wire signal_774 ;
    wire signal_775 ;
    wire signal_776 ;
    wire signal_777 ;
    wire signal_778 ;
    wire signal_779 ;
    wire signal_780 ;
    wire signal_781 ;
    wire signal_782 ;
    wire signal_783 ;
    wire signal_784 ;
    wire signal_785 ;
    wire signal_786 ;
    wire signal_787 ;
    wire signal_788 ;
    wire signal_789 ;
    wire signal_790 ;
    wire signal_791 ;
    wire signal_792 ;
    wire signal_793 ;
    wire signal_794 ;
    wire signal_795 ;
    wire signal_796 ;
    wire signal_797 ;
    wire signal_798 ;
    wire signal_799 ;
    wire signal_800 ;
    wire signal_801 ;
    wire signal_802 ;
    wire signal_803 ;
    wire signal_804 ;
    wire signal_805 ;
    wire signal_806 ;
    wire signal_807 ;
    wire signal_808 ;
    wire signal_809 ;
    wire signal_810 ;
    wire signal_811 ;
    wire signal_812 ;
    wire signal_813 ;
    wire signal_814 ;
    wire signal_815 ;
    wire signal_816 ;
    wire signal_817 ;
    wire signal_818 ;
    wire signal_819 ;
    wire signal_820 ;
    wire signal_821 ;
    wire signal_822 ;
    wire signal_823 ;
    wire signal_824 ;
    wire signal_825 ;
    wire signal_826 ;
    wire signal_827 ;
    wire signal_828 ;
    wire signal_829 ;
    wire signal_830 ;
    wire signal_831 ;
    wire signal_832 ;
    wire signal_833 ;
    wire signal_834 ;
    wire signal_835 ;
    wire signal_836 ;
    wire signal_837 ;
    wire signal_838 ;
    wire signal_839 ;
    wire signal_840 ;
    wire signal_841 ;
    wire signal_842 ;
    wire signal_843 ;
    wire signal_844 ;
    wire signal_845 ;
    wire signal_846 ;
    wire signal_847 ;
    wire signal_848 ;
    wire signal_849 ;
    wire signal_850 ;
    wire signal_851 ;
    wire signal_852 ;
    wire signal_853 ;
    wire signal_854 ;
    wire signal_855 ;
    wire signal_856 ;
    wire signal_857 ;
    wire signal_858 ;
    wire signal_859 ;
    wire signal_860 ;
    wire signal_861 ;
    wire signal_862 ;
    wire signal_863 ;
    wire signal_864 ;
    wire signal_865 ;
    wire signal_866 ;
    wire signal_867 ;
    wire signal_868 ;
    wire signal_869 ;
    wire signal_870 ;
    wire signal_871 ;
    wire signal_872 ;
    wire signal_873 ;
    wire signal_874 ;
    wire signal_875 ;
    wire signal_876 ;
    wire signal_877 ;
    wire signal_878 ;
    wire signal_879 ;
    wire signal_880 ;
    wire signal_881 ;
    wire signal_882 ;
    wire signal_883 ;
    wire signal_884 ;
    wire signal_885 ;
    wire signal_886 ;
    wire signal_887 ;
    wire signal_888 ;
    wire signal_889 ;
    wire signal_890 ;
    wire signal_891 ;
    wire signal_892 ;
    wire signal_893 ;
    wire signal_894 ;
    wire signal_895 ;
    wire signal_896 ;
    wire signal_897 ;
    wire signal_898 ;
    wire signal_899 ;
    wire signal_900 ;
    wire signal_901 ;
    wire signal_902 ;
    wire signal_903 ;
    wire signal_904 ;
    wire signal_905 ;
    wire signal_906 ;
    wire signal_907 ;
    wire signal_908 ;
    wire signal_909 ;
    wire signal_910 ;
    wire signal_911 ;
    wire signal_912 ;
    wire signal_913 ;
    wire signal_914 ;
    wire signal_915 ;
    wire signal_916 ;
    wire signal_917 ;
    wire signal_918 ;
    wire signal_919 ;
    wire signal_920 ;
    wire signal_921 ;
    wire signal_922 ;
    wire signal_923 ;
    wire signal_924 ;
    wire signal_925 ;
    wire signal_926 ;
    wire signal_927 ;
    wire signal_928 ;
    wire signal_929 ;
    wire signal_930 ;
    wire signal_931 ;
    wire signal_932 ;
    wire signal_933 ;
    wire signal_934 ;
    wire signal_935 ;
    wire signal_936 ;
    wire signal_937 ;
    wire signal_938 ;
    wire signal_939 ;
    wire signal_940 ;
    wire signal_941 ;
    wire signal_942 ;
    wire signal_943 ;
    wire signal_944 ;
    wire signal_945 ;
    wire signal_946 ;
    wire signal_947 ;
    wire signal_948 ;
    wire signal_949 ;
    wire signal_950 ;
    wire signal_951 ;
    wire signal_952 ;
    wire signal_953 ;
    wire signal_954 ;
    wire signal_955 ;
    wire signal_956 ;
    wire signal_957 ;
    wire signal_958 ;
    wire signal_959 ;
    wire signal_960 ;
    wire signal_961 ;
    wire signal_962 ;
    wire signal_963 ;
    wire signal_964 ;
    wire signal_965 ;
    wire signal_966 ;
    wire signal_967 ;
    wire signal_968 ;
    wire signal_969 ;
    wire signal_970 ;
    wire signal_971 ;
    wire signal_972 ;
    wire signal_973 ;
    wire signal_974 ;
    wire signal_975 ;
    wire signal_976 ;
    wire signal_977 ;
    wire signal_978 ;
    wire signal_979 ;
    wire signal_980 ;
    wire signal_981 ;
    wire signal_982 ;
    wire signal_983 ;
    wire signal_984 ;
    wire signal_985 ;
    wire signal_986 ;
    wire signal_987 ;
    wire signal_988 ;
    wire signal_989 ;
    wire signal_990 ;
    wire signal_991 ;
    wire signal_992 ;
    wire signal_993 ;
    wire signal_994 ;
    wire signal_995 ;
    wire signal_996 ;
    wire signal_997 ;
    wire signal_998 ;
    wire signal_999 ;
    wire signal_1000 ;
    wire signal_1001 ;
    wire signal_1002 ;
    wire signal_1003 ;
    wire signal_1004 ;
    wire signal_1005 ;
    wire signal_1006 ;
    wire signal_1007 ;
    wire signal_1008 ;
    wire signal_1009 ;
    wire signal_1010 ;
    wire signal_1011 ;
    wire signal_1012 ;
    wire signal_1013 ;
    wire signal_1014 ;
    wire signal_1015 ;
    wire signal_1016 ;
    wire signal_1017 ;
    wire signal_1018 ;
    wire signal_1019 ;
    wire signal_1020 ;
    wire signal_1021 ;
    wire signal_1022 ;
    wire signal_1023 ;
    wire signal_1024 ;
    wire signal_1025 ;
    wire signal_1026 ;
    wire signal_1027 ;
    wire signal_1028 ;
    wire signal_1029 ;
    wire signal_1030 ;
    wire signal_1031 ;
    wire signal_1032 ;
    wire signal_1033 ;
    wire signal_1034 ;
    wire signal_1035 ;
    wire signal_1036 ;
    wire signal_1037 ;
    wire signal_1038 ;
    wire signal_1039 ;
    wire signal_1040 ;
    wire signal_1041 ;
    wire signal_1042 ;
    wire signal_1043 ;
    wire signal_1044 ;
    wire signal_1045 ;
    wire signal_1046 ;
    wire signal_1047 ;
    wire signal_1048 ;
    wire signal_1049 ;
    wire signal_1050 ;
    wire signal_1051 ;
    wire signal_1052 ;
    wire signal_1053 ;
    wire signal_1054 ;
    wire signal_1055 ;
    wire signal_1056 ;
    wire signal_1057 ;
    wire signal_1058 ;
    wire signal_1059 ;
    wire signal_1060 ;
    wire signal_1061 ;
    wire signal_1062 ;
    wire signal_1063 ;
    wire signal_1064 ;
    wire signal_1065 ;
    wire signal_1066 ;
    wire signal_1067 ;
    wire signal_1068 ;

    /* cells in depth 0 */
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_136 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[4], X_s1[4], X_s0[4]}), .c ({signal_280, signal_279, signal_151}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_137 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_284, signal_283, signal_152}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_138 ( .a ({X_s2[7], X_s1[7], X_s0[7]}), .b ({X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_288, signal_287, signal_153}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_139 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_290, signal_289, signal_154}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_140 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_294, signal_293, signal_155}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_141 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[5], X_s1[5], X_s0[5]}), .c ({signal_300, signal_299, signal_156}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_142 ( .a ({X_s2[6], X_s1[6], X_s0[6]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_302, signal_301, signal_157}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_143 ( .a ({X_s2[5], X_s1[5], X_s0[5]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_304, signal_303, signal_158}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_144 ( .a ({X_s2[4], X_s1[4], X_s0[4]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_308, signal_307, signal_159}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_145 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_310, signal_309, signal_160}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_146 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_294, signal_293, signal_155}), .c ({signal_312, signal_311, signal_161}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_147 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_300, signal_299, signal_156}), .c ({signal_314, signal_313, signal_162}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_148 ( .a ({signal_288, signal_287, signal_153}), .b ({signal_290, signal_289, signal_154}), .c ({signal_316, signal_315, signal_163}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_149 ( .a ({signal_294, signal_293, signal_155}), .b ({signal_302, signal_301, signal_157}), .c ({signal_318, signal_317, signal_164}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_150 ( .a ({signal_294, signal_293, signal_155}), .b ({signal_304, signal_303, signal_158}), .c ({signal_320, signal_319, signal_165}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_151 ( .a ({signal_300, signal_299, signal_156}), .b ({signal_308, signal_307, signal_159}), .c ({signal_322, signal_321, signal_166}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_152 ( .a ({signal_300, signal_299, signal_156}), .b ({signal_310, signal_309, signal_160}), .c ({signal_324, signal_323, signal_167}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_153 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_304, signal_303, signal_158}), .c ({signal_326, signal_325, signal_168}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_160 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_312, signal_311, signal_161}), .c ({signal_340, signal_339, signal_175}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_161 ( .a ({signal_300, signal_299, signal_156}), .b ({signal_312, signal_311, signal_161}), .c ({signal_342, signal_341, signal_176}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_162 ( .a ({signal_302, signal_301, signal_157}), .b ({signal_312, signal_311, signal_161}), .c ({signal_344, signal_343, signal_177}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_163 ( .a ({signal_314, signal_313, signal_162}), .b ({signal_320, signal_319, signal_165}), .c ({signal_346, signal_345, signal_178}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_164 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_322, signal_321, signal_166}), .c ({signal_348, signal_347, signal_179}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_165 ( .a ({signal_284, signal_283, signal_152}), .b ({signal_324, signal_323, signal_167}), .c ({signal_350, signal_349, signal_180}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_166 ( .a ({signal_288, signal_287, signal_153}), .b ({signal_320, signal_319, signal_165}), .c ({signal_352, signal_351, signal_181}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_170 ( .a ({signal_284, signal_283, signal_152}), .b ({signal_342, signal_341, signal_176}), .c ({signal_360, signal_359, signal_185}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_171 ( .a ({signal_346, signal_345, signal_178}), .b ({signal_348, signal_347, signal_179}), .c ({signal_362, signal_361, signal_186}) ) ;

    /* cells in depth 1 */
    buf_clk cell_268 ( .C (clk), .D (signal_177), .Q (signal_673) ) ;
    buf_clk cell_270 ( .C (clk), .D (signal_343), .Q (signal_675) ) ;
    buf_clk cell_272 ( .C (clk), .D (signal_344), .Q (signal_677) ) ;
    buf_clk cell_274 ( .C (clk), .D (signal_181), .Q (signal_679) ) ;
    buf_clk cell_276 ( .C (clk), .D (signal_351), .Q (signal_681) ) ;
    buf_clk cell_278 ( .C (clk), .D (signal_352), .Q (signal_683) ) ;
    buf_clk cell_280 ( .C (clk), .D (signal_185), .Q (signal_685) ) ;
    buf_clk cell_282 ( .C (clk), .D (signal_359), .Q (signal_687) ) ;
    buf_clk cell_284 ( .C (clk), .D (signal_360), .Q (signal_689) ) ;
    buf_clk cell_286 ( .C (clk), .D (signal_186), .Q (signal_691) ) ;
    buf_clk cell_288 ( .C (clk), .D (signal_361), .Q (signal_693) ) ;
    buf_clk cell_290 ( .C (clk), .D (signal_362), .Q (signal_695) ) ;
    buf_clk cell_340 ( .C (clk), .D (signal_175), .Q (signal_745) ) ;
    buf_clk cell_346 ( .C (clk), .D (signal_339), .Q (signal_751) ) ;
    buf_clk cell_352 ( .C (clk), .D (signal_340), .Q (signal_757) ) ;
    buf_clk cell_358 ( .C (clk), .D (X_s0[0]), .Q (signal_763) ) ;
    buf_clk cell_364 ( .C (clk), .D (X_s1[0]), .Q (signal_769) ) ;
    buf_clk cell_370 ( .C (clk), .D (X_s2[0]), .Q (signal_775) ) ;
    buf_clk cell_376 ( .C (clk), .D (signal_162), .Q (signal_781) ) ;
    buf_clk cell_382 ( .C (clk), .D (signal_313), .Q (signal_787) ) ;
    buf_clk cell_388 ( .C (clk), .D (signal_314), .Q (signal_793) ) ;
    buf_clk cell_394 ( .C (clk), .D (signal_178), .Q (signal_799) ) ;
    buf_clk cell_400 ( .C (clk), .D (signal_345), .Q (signal_805) ) ;
    buf_clk cell_406 ( .C (clk), .D (signal_346), .Q (signal_811) ) ;
    buf_clk cell_412 ( .C (clk), .D (signal_180), .Q (signal_817) ) ;
    buf_clk cell_418 ( .C (clk), .D (signal_349), .Q (signal_823) ) ;
    buf_clk cell_424 ( .C (clk), .D (signal_350), .Q (signal_829) ) ;
    buf_clk cell_430 ( .C (clk), .D (signal_166), .Q (signal_835) ) ;
    buf_clk cell_436 ( .C (clk), .D (signal_321), .Q (signal_841) ) ;
    buf_clk cell_442 ( .C (clk), .D (signal_322), .Q (signal_847) ) ;
    buf_clk cell_448 ( .C (clk), .D (signal_167), .Q (signal_853) ) ;
    buf_clk cell_454 ( .C (clk), .D (signal_323), .Q (signal_859) ) ;
    buf_clk cell_460 ( .C (clk), .D (signal_324), .Q (signal_865) ) ;
    buf_clk cell_466 ( .C (clk), .D (signal_179), .Q (signal_871) ) ;
    buf_clk cell_472 ( .C (clk), .D (signal_347), .Q (signal_877) ) ;
    buf_clk cell_478 ( .C (clk), .D (signal_348), .Q (signal_883) ) ;
    buf_clk cell_484 ( .C (clk), .D (signal_161), .Q (signal_889) ) ;
    buf_clk cell_490 ( .C (clk), .D (signal_311), .Q (signal_895) ) ;
    buf_clk cell_496 ( .C (clk), .D (signal_312), .Q (signal_901) ) ;
    buf_clk cell_502 ( .C (clk), .D (signal_165), .Q (signal_907) ) ;
    buf_clk cell_508 ( .C (clk), .D (signal_319), .Q (signal_913) ) ;
    buf_clk cell_514 ( .C (clk), .D (signal_320), .Q (signal_919) ) ;
    buf_clk cell_520 ( .C (clk), .D (signal_164), .Q (signal_925) ) ;
    buf_clk cell_526 ( .C (clk), .D (signal_317), .Q (signal_931) ) ;
    buf_clk cell_532 ( .C (clk), .D (signal_318), .Q (signal_937) ) ;
    buf_clk cell_538 ( .C (clk), .D (signal_176), .Q (signal_943) ) ;
    buf_clk cell_544 ( .C (clk), .D (signal_341), .Q (signal_949) ) ;
    buf_clk cell_550 ( .C (clk), .D (signal_342), .Q (signal_955) ) ;
    buf_clk cell_556 ( .C (clk), .D (signal_163), .Q (signal_961) ) ;
    buf_clk cell_562 ( .C (clk), .D (signal_315), .Q (signal_967) ) ;
    buf_clk cell_568 ( .C (clk), .D (signal_316), .Q (signal_973) ) ;
    buf_clk cell_574 ( .C (clk), .D (signal_153), .Q (signal_979) ) ;
    buf_clk cell_580 ( .C (clk), .D (signal_287), .Q (signal_985) ) ;
    buf_clk cell_586 ( .C (clk), .D (signal_288), .Q (signal_991) ) ;
    buf_clk cell_592 ( .C (clk), .D (signal_151), .Q (signal_997) ) ;
    buf_clk cell_598 ( .C (clk), .D (signal_279), .Q (signal_1003) ) ;
    buf_clk cell_604 ( .C (clk), .D (signal_280), .Q (signal_1009) ) ;
    buf_clk cell_610 ( .C (clk), .D (signal_152), .Q (signal_1015) ) ;
    buf_clk cell_616 ( .C (clk), .D (signal_283), .Q (signal_1021) ) ;
    buf_clk cell_622 ( .C (clk), .D (signal_284), .Q (signal_1027) ) ;
    buf_clk cell_628 ( .C (clk), .D (signal_168), .Q (signal_1033) ) ;
    buf_clk cell_634 ( .C (clk), .D (signal_325), .Q (signal_1039) ) ;
    buf_clk cell_640 ( .C (clk), .D (signal_326), .Q (signal_1045) ) ;
    buf_clk cell_646 ( .C (clk), .D (signal_154), .Q (signal_1051) ) ;
    buf_clk cell_652 ( .C (clk), .D (signal_289), .Q (signal_1057) ) ;
    buf_clk cell_658 ( .C (clk), .D (signal_290), .Q (signal_1063) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_154 ( .a ({signal_312, signal_311, signal_161}), .b ({signal_316, signal_315, signal_163}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_328, signal_327, signal_169}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_155 ( .a ({X_s2[0], X_s1[0], X_s0[0]}), .b ({signal_322, signal_321, signal_166}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_330, signal_329, signal_170}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_156 ( .a ({signal_288, signal_287, signal_153}), .b ({signal_320, signal_319, signal_165}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_332, signal_331, signal_171}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_157 ( .a ({signal_314, signal_313, signal_162}), .b ({signal_324, signal_323, signal_167}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_334, signal_333, signal_172}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_158 ( .a ({signal_280, signal_279, signal_151}), .b ({signal_318, signal_317, signal_164}), .clk (clk), .r ({Fresh[14], Fresh[13], Fresh[12]}), .c ({signal_336, signal_335, signal_173}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_159 ( .a ({signal_290, signal_289, signal_154}), .b ({signal_326, signal_325, signal_168}), .clk (clk), .r ({Fresh[17], Fresh[16], Fresh[15]}), .c ({signal_338, signal_337, signal_174}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_167 ( .a ({signal_340, signal_339, signal_175}), .b ({signal_350, signal_349, signal_180}), .clk (clk), .r ({Fresh[20], Fresh[19], Fresh[18]}), .c ({signal_354, signal_353, signal_182}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_168 ( .a ({signal_346, signal_345, signal_178}), .b ({signal_348, signal_347, signal_179}), .clk (clk), .r ({Fresh[23], Fresh[22], Fresh[21]}), .c ({signal_356, signal_355, signal_183}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_169 ( .a ({signal_284, signal_283, signal_152}), .b ({signal_342, signal_341, signal_176}), .clk (clk), .r ({Fresh[26], Fresh[25], Fresh[24]}), .c ({signal_358, signal_357, signal_184}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_172 ( .a ({signal_678, signal_676, signal_674}), .b ({signal_328, signal_327, signal_169}), .c ({signal_364, signal_363, signal_187}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_173 ( .a ({signal_328, signal_327, signal_169}), .b ({signal_330, signal_329, signal_170}), .c ({signal_366, signal_365, signal_188}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_174 ( .a ({signal_684, signal_682, signal_680}), .b ({signal_332, signal_331, signal_171}), .c ({signal_368, signal_367, signal_189}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_175 ( .a ({signal_336, signal_335, signal_173}), .b ({signal_338, signal_337, signal_174}), .c ({signal_370, signal_369, signal_190}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_176 ( .a ({signal_332, signal_331, signal_171}), .b ({signal_356, signal_355, signal_183}), .c ({signal_372, signal_371, signal_191}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_177 ( .a ({signal_336, signal_335, signal_173}), .b ({signal_358, signal_357, signal_184}), .c ({signal_374, signal_373, signal_192}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_178 ( .a ({signal_354, signal_353, signal_182}), .b ({signal_364, signal_363, signal_187}), .c ({signal_376, signal_375, signal_193}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_179 ( .a ({signal_690, signal_688, signal_686}), .b ({signal_366, signal_365, signal_188}), .c ({signal_378, signal_377, signal_194}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_180 ( .a ({signal_334, signal_333, signal_172}), .b ({signal_368, signal_367, signal_189}), .c ({signal_380, signal_379, signal_195}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_181 ( .a ({signal_372, signal_371, signal_191}), .b ({signal_374, signal_373, signal_192}), .c ({signal_382, signal_381, signal_196}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_182 ( .a ({signal_370, signal_369, signal_190}), .b ({signal_376, signal_375, signal_193}), .c ({signal_384, signal_383, signal_197}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_183 ( .a ({signal_374, signal_373, signal_192}), .b ({signal_378, signal_377, signal_194}), .c ({signal_386, signal_385, signal_198}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_184 ( .a ({signal_370, signal_369, signal_190}), .b ({signal_380, signal_379, signal_195}), .c ({signal_388, signal_387, signal_199}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_187 ( .a ({signal_696, signal_694, signal_692}), .b ({signal_382, signal_381, signal_196}), .c ({signal_394, signal_393, signal_202}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_188 ( .a ({signal_384, signal_383, signal_197}), .b ({signal_386, signal_385, signal_198}), .c ({signal_396, signal_395, signal_203}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_190 ( .a ({signal_388, signal_387, signal_199}), .b ({signal_394, signal_393, signal_202}), .c ({signal_400, signal_399, signal_205}) ) ;
    buf_clk cell_269 ( .C (clk), .D (signal_673), .Q (signal_674) ) ;
    buf_clk cell_271 ( .C (clk), .D (signal_675), .Q (signal_676) ) ;
    buf_clk cell_273 ( .C (clk), .D (signal_677), .Q (signal_678) ) ;
    buf_clk cell_275 ( .C (clk), .D (signal_679), .Q (signal_680) ) ;
    buf_clk cell_277 ( .C (clk), .D (signal_681), .Q (signal_682) ) ;
    buf_clk cell_279 ( .C (clk), .D (signal_683), .Q (signal_684) ) ;
    buf_clk cell_281 ( .C (clk), .D (signal_685), .Q (signal_686) ) ;
    buf_clk cell_283 ( .C (clk), .D (signal_687), .Q (signal_688) ) ;
    buf_clk cell_285 ( .C (clk), .D (signal_689), .Q (signal_690) ) ;
    buf_clk cell_287 ( .C (clk), .D (signal_691), .Q (signal_692) ) ;
    buf_clk cell_289 ( .C (clk), .D (signal_693), .Q (signal_694) ) ;
    buf_clk cell_291 ( .C (clk), .D (signal_695), .Q (signal_696) ) ;
    buf_clk cell_341 ( .C (clk), .D (signal_745), .Q (signal_746) ) ;
    buf_clk cell_347 ( .C (clk), .D (signal_751), .Q (signal_752) ) ;
    buf_clk cell_353 ( .C (clk), .D (signal_757), .Q (signal_758) ) ;
    buf_clk cell_359 ( .C (clk), .D (signal_763), .Q (signal_764) ) ;
    buf_clk cell_365 ( .C (clk), .D (signal_769), .Q (signal_770) ) ;
    buf_clk cell_371 ( .C (clk), .D (signal_775), .Q (signal_776) ) ;
    buf_clk cell_377 ( .C (clk), .D (signal_781), .Q (signal_782) ) ;
    buf_clk cell_383 ( .C (clk), .D (signal_787), .Q (signal_788) ) ;
    buf_clk cell_389 ( .C (clk), .D (signal_793), .Q (signal_794) ) ;
    buf_clk cell_395 ( .C (clk), .D (signal_799), .Q (signal_800) ) ;
    buf_clk cell_401 ( .C (clk), .D (signal_805), .Q (signal_806) ) ;
    buf_clk cell_407 ( .C (clk), .D (signal_811), .Q (signal_812) ) ;
    buf_clk cell_413 ( .C (clk), .D (signal_817), .Q (signal_818) ) ;
    buf_clk cell_419 ( .C (clk), .D (signal_823), .Q (signal_824) ) ;
    buf_clk cell_425 ( .C (clk), .D (signal_829), .Q (signal_830) ) ;
    buf_clk cell_431 ( .C (clk), .D (signal_835), .Q (signal_836) ) ;
    buf_clk cell_437 ( .C (clk), .D (signal_841), .Q (signal_842) ) ;
    buf_clk cell_443 ( .C (clk), .D (signal_847), .Q (signal_848) ) ;
    buf_clk cell_449 ( .C (clk), .D (signal_853), .Q (signal_854) ) ;
    buf_clk cell_455 ( .C (clk), .D (signal_859), .Q (signal_860) ) ;
    buf_clk cell_461 ( .C (clk), .D (signal_865), .Q (signal_866) ) ;
    buf_clk cell_467 ( .C (clk), .D (signal_871), .Q (signal_872) ) ;
    buf_clk cell_473 ( .C (clk), .D (signal_877), .Q (signal_878) ) ;
    buf_clk cell_479 ( .C (clk), .D (signal_883), .Q (signal_884) ) ;
    buf_clk cell_485 ( .C (clk), .D (signal_889), .Q (signal_890) ) ;
    buf_clk cell_491 ( .C (clk), .D (signal_895), .Q (signal_896) ) ;
    buf_clk cell_497 ( .C (clk), .D (signal_901), .Q (signal_902) ) ;
    buf_clk cell_503 ( .C (clk), .D (signal_907), .Q (signal_908) ) ;
    buf_clk cell_509 ( .C (clk), .D (signal_913), .Q (signal_914) ) ;
    buf_clk cell_515 ( .C (clk), .D (signal_919), .Q (signal_920) ) ;
    buf_clk cell_521 ( .C (clk), .D (signal_925), .Q (signal_926) ) ;
    buf_clk cell_527 ( .C (clk), .D (signal_931), .Q (signal_932) ) ;
    buf_clk cell_533 ( .C (clk), .D (signal_937), .Q (signal_938) ) ;
    buf_clk cell_539 ( .C (clk), .D (signal_943), .Q (signal_944) ) ;
    buf_clk cell_545 ( .C (clk), .D (signal_949), .Q (signal_950) ) ;
    buf_clk cell_551 ( .C (clk), .D (signal_955), .Q (signal_956) ) ;
    buf_clk cell_557 ( .C (clk), .D (signal_961), .Q (signal_962) ) ;
    buf_clk cell_563 ( .C (clk), .D (signal_967), .Q (signal_968) ) ;
    buf_clk cell_569 ( .C (clk), .D (signal_973), .Q (signal_974) ) ;
    buf_clk cell_575 ( .C (clk), .D (signal_979), .Q (signal_980) ) ;
    buf_clk cell_581 ( .C (clk), .D (signal_985), .Q (signal_986) ) ;
    buf_clk cell_587 ( .C (clk), .D (signal_991), .Q (signal_992) ) ;
    buf_clk cell_593 ( .C (clk), .D (signal_997), .Q (signal_998) ) ;
    buf_clk cell_599 ( .C (clk), .D (signal_1003), .Q (signal_1004) ) ;
    buf_clk cell_605 ( .C (clk), .D (signal_1009), .Q (signal_1010) ) ;
    buf_clk cell_611 ( .C (clk), .D (signal_1015), .Q (signal_1016) ) ;
    buf_clk cell_617 ( .C (clk), .D (signal_1021), .Q (signal_1022) ) ;
    buf_clk cell_623 ( .C (clk), .D (signal_1027), .Q (signal_1028) ) ;
    buf_clk cell_629 ( .C (clk), .D (signal_1033), .Q (signal_1034) ) ;
    buf_clk cell_635 ( .C (clk), .D (signal_1039), .Q (signal_1040) ) ;
    buf_clk cell_641 ( .C (clk), .D (signal_1045), .Q (signal_1046) ) ;
    buf_clk cell_647 ( .C (clk), .D (signal_1051), .Q (signal_1052) ) ;
    buf_clk cell_653 ( .C (clk), .D (signal_1057), .Q (signal_1058) ) ;
    buf_clk cell_659 ( .C (clk), .D (signal_1063), .Q (signal_1064) ) ;

    /* cells in depth 3 */
    buf_clk cell_292 ( .C (clk), .D (signal_198), .Q (signal_697) ) ;
    buf_clk cell_294 ( .C (clk), .D (signal_385), .Q (signal_699) ) ;
    buf_clk cell_296 ( .C (clk), .D (signal_386), .Q (signal_701) ) ;
    buf_clk cell_298 ( .C (clk), .D (signal_202), .Q (signal_703) ) ;
    buf_clk cell_300 ( .C (clk), .D (signal_393), .Q (signal_705) ) ;
    buf_clk cell_302 ( .C (clk), .D (signal_394), .Q (signal_707) ) ;
    buf_clk cell_304 ( .C (clk), .D (signal_203), .Q (signal_709) ) ;
    buf_clk cell_306 ( .C (clk), .D (signal_395), .Q (signal_711) ) ;
    buf_clk cell_308 ( .C (clk), .D (signal_396), .Q (signal_713) ) ;
    buf_clk cell_310 ( .C (clk), .D (signal_205), .Q (signal_715) ) ;
    buf_clk cell_312 ( .C (clk), .D (signal_399), .Q (signal_717) ) ;
    buf_clk cell_314 ( .C (clk), .D (signal_400), .Q (signal_719) ) ;
    buf_clk cell_342 ( .C (clk), .D (signal_746), .Q (signal_747) ) ;
    buf_clk cell_348 ( .C (clk), .D (signal_752), .Q (signal_753) ) ;
    buf_clk cell_354 ( .C (clk), .D (signal_758), .Q (signal_759) ) ;
    buf_clk cell_360 ( .C (clk), .D (signal_764), .Q (signal_765) ) ;
    buf_clk cell_366 ( .C (clk), .D (signal_770), .Q (signal_771) ) ;
    buf_clk cell_372 ( .C (clk), .D (signal_776), .Q (signal_777) ) ;
    buf_clk cell_378 ( .C (clk), .D (signal_782), .Q (signal_783) ) ;
    buf_clk cell_384 ( .C (clk), .D (signal_788), .Q (signal_789) ) ;
    buf_clk cell_390 ( .C (clk), .D (signal_794), .Q (signal_795) ) ;
    buf_clk cell_396 ( .C (clk), .D (signal_800), .Q (signal_801) ) ;
    buf_clk cell_402 ( .C (clk), .D (signal_806), .Q (signal_807) ) ;
    buf_clk cell_408 ( .C (clk), .D (signal_812), .Q (signal_813) ) ;
    buf_clk cell_414 ( .C (clk), .D (signal_818), .Q (signal_819) ) ;
    buf_clk cell_420 ( .C (clk), .D (signal_824), .Q (signal_825) ) ;
    buf_clk cell_426 ( .C (clk), .D (signal_830), .Q (signal_831) ) ;
    buf_clk cell_432 ( .C (clk), .D (signal_836), .Q (signal_837) ) ;
    buf_clk cell_438 ( .C (clk), .D (signal_842), .Q (signal_843) ) ;
    buf_clk cell_444 ( .C (clk), .D (signal_848), .Q (signal_849) ) ;
    buf_clk cell_450 ( .C (clk), .D (signal_854), .Q (signal_855) ) ;
    buf_clk cell_456 ( .C (clk), .D (signal_860), .Q (signal_861) ) ;
    buf_clk cell_462 ( .C (clk), .D (signal_866), .Q (signal_867) ) ;
    buf_clk cell_468 ( .C (clk), .D (signal_872), .Q (signal_873) ) ;
    buf_clk cell_474 ( .C (clk), .D (signal_878), .Q (signal_879) ) ;
    buf_clk cell_480 ( .C (clk), .D (signal_884), .Q (signal_885) ) ;
    buf_clk cell_486 ( .C (clk), .D (signal_890), .Q (signal_891) ) ;
    buf_clk cell_492 ( .C (clk), .D (signal_896), .Q (signal_897) ) ;
    buf_clk cell_498 ( .C (clk), .D (signal_902), .Q (signal_903) ) ;
    buf_clk cell_504 ( .C (clk), .D (signal_908), .Q (signal_909) ) ;
    buf_clk cell_510 ( .C (clk), .D (signal_914), .Q (signal_915) ) ;
    buf_clk cell_516 ( .C (clk), .D (signal_920), .Q (signal_921) ) ;
    buf_clk cell_522 ( .C (clk), .D (signal_926), .Q (signal_927) ) ;
    buf_clk cell_528 ( .C (clk), .D (signal_932), .Q (signal_933) ) ;
    buf_clk cell_534 ( .C (clk), .D (signal_938), .Q (signal_939) ) ;
    buf_clk cell_540 ( .C (clk), .D (signal_944), .Q (signal_945) ) ;
    buf_clk cell_546 ( .C (clk), .D (signal_950), .Q (signal_951) ) ;
    buf_clk cell_552 ( .C (clk), .D (signal_956), .Q (signal_957) ) ;
    buf_clk cell_558 ( .C (clk), .D (signal_962), .Q (signal_963) ) ;
    buf_clk cell_564 ( .C (clk), .D (signal_968), .Q (signal_969) ) ;
    buf_clk cell_570 ( .C (clk), .D (signal_974), .Q (signal_975) ) ;
    buf_clk cell_576 ( .C (clk), .D (signal_980), .Q (signal_981) ) ;
    buf_clk cell_582 ( .C (clk), .D (signal_986), .Q (signal_987) ) ;
    buf_clk cell_588 ( .C (clk), .D (signal_992), .Q (signal_993) ) ;
    buf_clk cell_594 ( .C (clk), .D (signal_998), .Q (signal_999) ) ;
    buf_clk cell_600 ( .C (clk), .D (signal_1004), .Q (signal_1005) ) ;
    buf_clk cell_606 ( .C (clk), .D (signal_1010), .Q (signal_1011) ) ;
    buf_clk cell_612 ( .C (clk), .D (signal_1016), .Q (signal_1017) ) ;
    buf_clk cell_618 ( .C (clk), .D (signal_1022), .Q (signal_1023) ) ;
    buf_clk cell_624 ( .C (clk), .D (signal_1028), .Q (signal_1029) ) ;
    buf_clk cell_630 ( .C (clk), .D (signal_1034), .Q (signal_1035) ) ;
    buf_clk cell_636 ( .C (clk), .D (signal_1040), .Q (signal_1041) ) ;
    buf_clk cell_642 ( .C (clk), .D (signal_1046), .Q (signal_1047) ) ;
    buf_clk cell_648 ( .C (clk), .D (signal_1052), .Q (signal_1053) ) ;
    buf_clk cell_654 ( .C (clk), .D (signal_1058), .Q (signal_1059) ) ;
    buf_clk cell_660 ( .C (clk), .D (signal_1064), .Q (signal_1065) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_185 ( .a ({signal_384, signal_383, signal_197}), .b ({signal_388, signal_387, signal_199}), .clk (clk), .r ({Fresh[29], Fresh[28], Fresh[27]}), .c ({signal_390, signal_389, signal_200}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_186 ( .a ({signal_386, signal_385, signal_198}), .b ({signal_388, signal_387, signal_199}), .clk (clk), .r ({Fresh[32], Fresh[31], Fresh[30]}), .c ({signal_392, signal_391, signal_201}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_189 ( .a ({signal_384, signal_383, signal_197}), .b ({signal_394, signal_393, signal_202}), .clk (clk), .r ({Fresh[35], Fresh[34], Fresh[33]}), .c ({signal_398, signal_397, signal_204}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_191 ( .a ({signal_702, signal_700, signal_698}), .b ({signal_390, signal_389, signal_200}), .c ({signal_402, signal_401, signal_206}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_192 ( .a ({signal_708, signal_706, signal_704}), .b ({signal_390, signal_389, signal_200}), .c ({signal_404, signal_403, signal_207}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_193 ( .a ({signal_390, signal_389, signal_200}), .b ({signal_714, signal_712, signal_710}), .c ({signal_406, signal_405, signal_208}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_198 ( .a ({signal_390, signal_389, signal_200}), .b ({signal_720, signal_718, signal_716}), .c ({signal_416, signal_415, signal_213}) ) ;
    buf_clk cell_293 ( .C (clk), .D (signal_697), .Q (signal_698) ) ;
    buf_clk cell_295 ( .C (clk), .D (signal_699), .Q (signal_700) ) ;
    buf_clk cell_297 ( .C (clk), .D (signal_701), .Q (signal_702) ) ;
    buf_clk cell_299 ( .C (clk), .D (signal_703), .Q (signal_704) ) ;
    buf_clk cell_301 ( .C (clk), .D (signal_705), .Q (signal_706) ) ;
    buf_clk cell_303 ( .C (clk), .D (signal_707), .Q (signal_708) ) ;
    buf_clk cell_305 ( .C (clk), .D (signal_709), .Q (signal_710) ) ;
    buf_clk cell_307 ( .C (clk), .D (signal_711), .Q (signal_712) ) ;
    buf_clk cell_309 ( .C (clk), .D (signal_713), .Q (signal_714) ) ;
    buf_clk cell_311 ( .C (clk), .D (signal_715), .Q (signal_716) ) ;
    buf_clk cell_313 ( .C (clk), .D (signal_717), .Q (signal_718) ) ;
    buf_clk cell_315 ( .C (clk), .D (signal_719), .Q (signal_720) ) ;
    buf_clk cell_343 ( .C (clk), .D (signal_747), .Q (signal_748) ) ;
    buf_clk cell_349 ( .C (clk), .D (signal_753), .Q (signal_754) ) ;
    buf_clk cell_355 ( .C (clk), .D (signal_759), .Q (signal_760) ) ;
    buf_clk cell_361 ( .C (clk), .D (signal_765), .Q (signal_766) ) ;
    buf_clk cell_367 ( .C (clk), .D (signal_771), .Q (signal_772) ) ;
    buf_clk cell_373 ( .C (clk), .D (signal_777), .Q (signal_778) ) ;
    buf_clk cell_379 ( .C (clk), .D (signal_783), .Q (signal_784) ) ;
    buf_clk cell_385 ( .C (clk), .D (signal_789), .Q (signal_790) ) ;
    buf_clk cell_391 ( .C (clk), .D (signal_795), .Q (signal_796) ) ;
    buf_clk cell_397 ( .C (clk), .D (signal_801), .Q (signal_802) ) ;
    buf_clk cell_403 ( .C (clk), .D (signal_807), .Q (signal_808) ) ;
    buf_clk cell_409 ( .C (clk), .D (signal_813), .Q (signal_814) ) ;
    buf_clk cell_415 ( .C (clk), .D (signal_819), .Q (signal_820) ) ;
    buf_clk cell_421 ( .C (clk), .D (signal_825), .Q (signal_826) ) ;
    buf_clk cell_427 ( .C (clk), .D (signal_831), .Q (signal_832) ) ;
    buf_clk cell_433 ( .C (clk), .D (signal_837), .Q (signal_838) ) ;
    buf_clk cell_439 ( .C (clk), .D (signal_843), .Q (signal_844) ) ;
    buf_clk cell_445 ( .C (clk), .D (signal_849), .Q (signal_850) ) ;
    buf_clk cell_451 ( .C (clk), .D (signal_855), .Q (signal_856) ) ;
    buf_clk cell_457 ( .C (clk), .D (signal_861), .Q (signal_862) ) ;
    buf_clk cell_463 ( .C (clk), .D (signal_867), .Q (signal_868) ) ;
    buf_clk cell_469 ( .C (clk), .D (signal_873), .Q (signal_874) ) ;
    buf_clk cell_475 ( .C (clk), .D (signal_879), .Q (signal_880) ) ;
    buf_clk cell_481 ( .C (clk), .D (signal_885), .Q (signal_886) ) ;
    buf_clk cell_487 ( .C (clk), .D (signal_891), .Q (signal_892) ) ;
    buf_clk cell_493 ( .C (clk), .D (signal_897), .Q (signal_898) ) ;
    buf_clk cell_499 ( .C (clk), .D (signal_903), .Q (signal_904) ) ;
    buf_clk cell_505 ( .C (clk), .D (signal_909), .Q (signal_910) ) ;
    buf_clk cell_511 ( .C (clk), .D (signal_915), .Q (signal_916) ) ;
    buf_clk cell_517 ( .C (clk), .D (signal_921), .Q (signal_922) ) ;
    buf_clk cell_523 ( .C (clk), .D (signal_927), .Q (signal_928) ) ;
    buf_clk cell_529 ( .C (clk), .D (signal_933), .Q (signal_934) ) ;
    buf_clk cell_535 ( .C (clk), .D (signal_939), .Q (signal_940) ) ;
    buf_clk cell_541 ( .C (clk), .D (signal_945), .Q (signal_946) ) ;
    buf_clk cell_547 ( .C (clk), .D (signal_951), .Q (signal_952) ) ;
    buf_clk cell_553 ( .C (clk), .D (signal_957), .Q (signal_958) ) ;
    buf_clk cell_559 ( .C (clk), .D (signal_963), .Q (signal_964) ) ;
    buf_clk cell_565 ( .C (clk), .D (signal_969), .Q (signal_970) ) ;
    buf_clk cell_571 ( .C (clk), .D (signal_975), .Q (signal_976) ) ;
    buf_clk cell_577 ( .C (clk), .D (signal_981), .Q (signal_982) ) ;
    buf_clk cell_583 ( .C (clk), .D (signal_987), .Q (signal_988) ) ;
    buf_clk cell_589 ( .C (clk), .D (signal_993), .Q (signal_994) ) ;
    buf_clk cell_595 ( .C (clk), .D (signal_999), .Q (signal_1000) ) ;
    buf_clk cell_601 ( .C (clk), .D (signal_1005), .Q (signal_1006) ) ;
    buf_clk cell_607 ( .C (clk), .D (signal_1011), .Q (signal_1012) ) ;
    buf_clk cell_613 ( .C (clk), .D (signal_1017), .Q (signal_1018) ) ;
    buf_clk cell_619 ( .C (clk), .D (signal_1023), .Q (signal_1024) ) ;
    buf_clk cell_625 ( .C (clk), .D (signal_1029), .Q (signal_1030) ) ;
    buf_clk cell_631 ( .C (clk), .D (signal_1035), .Q (signal_1036) ) ;
    buf_clk cell_637 ( .C (clk), .D (signal_1041), .Q (signal_1042) ) ;
    buf_clk cell_643 ( .C (clk), .D (signal_1047), .Q (signal_1048) ) ;
    buf_clk cell_649 ( .C (clk), .D (signal_1053), .Q (signal_1054) ) ;
    buf_clk cell_655 ( .C (clk), .D (signal_1059), .Q (signal_1060) ) ;
    buf_clk cell_661 ( .C (clk), .D (signal_1065), .Q (signal_1066) ) ;

    /* cells in depth 5 */
    buf_clk cell_316 ( .C (clk), .D (signal_698), .Q (signal_721) ) ;
    buf_clk cell_318 ( .C (clk), .D (signal_700), .Q (signal_723) ) ;
    buf_clk cell_320 ( .C (clk), .D (signal_702), .Q (signal_725) ) ;
    buf_clk cell_322 ( .C (clk), .D (signal_208), .Q (signal_727) ) ;
    buf_clk cell_324 ( .C (clk), .D (signal_405), .Q (signal_729) ) ;
    buf_clk cell_326 ( .C (clk), .D (signal_406), .Q (signal_731) ) ;
    buf_clk cell_328 ( .C (clk), .D (signal_704), .Q (signal_733) ) ;
    buf_clk cell_330 ( .C (clk), .D (signal_706), .Q (signal_735) ) ;
    buf_clk cell_332 ( .C (clk), .D (signal_708), .Q (signal_737) ) ;
    buf_clk cell_334 ( .C (clk), .D (signal_213), .Q (signal_739) ) ;
    buf_clk cell_336 ( .C (clk), .D (signal_415), .Q (signal_741) ) ;
    buf_clk cell_338 ( .C (clk), .D (signal_416), .Q (signal_743) ) ;
    buf_clk cell_344 ( .C (clk), .D (signal_748), .Q (signal_749) ) ;
    buf_clk cell_350 ( .C (clk), .D (signal_754), .Q (signal_755) ) ;
    buf_clk cell_356 ( .C (clk), .D (signal_760), .Q (signal_761) ) ;
    buf_clk cell_362 ( .C (clk), .D (signal_766), .Q (signal_767) ) ;
    buf_clk cell_368 ( .C (clk), .D (signal_772), .Q (signal_773) ) ;
    buf_clk cell_374 ( .C (clk), .D (signal_778), .Q (signal_779) ) ;
    buf_clk cell_380 ( .C (clk), .D (signal_784), .Q (signal_785) ) ;
    buf_clk cell_386 ( .C (clk), .D (signal_790), .Q (signal_791) ) ;
    buf_clk cell_392 ( .C (clk), .D (signal_796), .Q (signal_797) ) ;
    buf_clk cell_398 ( .C (clk), .D (signal_802), .Q (signal_803) ) ;
    buf_clk cell_404 ( .C (clk), .D (signal_808), .Q (signal_809) ) ;
    buf_clk cell_410 ( .C (clk), .D (signal_814), .Q (signal_815) ) ;
    buf_clk cell_416 ( .C (clk), .D (signal_820), .Q (signal_821) ) ;
    buf_clk cell_422 ( .C (clk), .D (signal_826), .Q (signal_827) ) ;
    buf_clk cell_428 ( .C (clk), .D (signal_832), .Q (signal_833) ) ;
    buf_clk cell_434 ( .C (clk), .D (signal_838), .Q (signal_839) ) ;
    buf_clk cell_440 ( .C (clk), .D (signal_844), .Q (signal_845) ) ;
    buf_clk cell_446 ( .C (clk), .D (signal_850), .Q (signal_851) ) ;
    buf_clk cell_452 ( .C (clk), .D (signal_856), .Q (signal_857) ) ;
    buf_clk cell_458 ( .C (clk), .D (signal_862), .Q (signal_863) ) ;
    buf_clk cell_464 ( .C (clk), .D (signal_868), .Q (signal_869) ) ;
    buf_clk cell_470 ( .C (clk), .D (signal_874), .Q (signal_875) ) ;
    buf_clk cell_476 ( .C (clk), .D (signal_880), .Q (signal_881) ) ;
    buf_clk cell_482 ( .C (clk), .D (signal_886), .Q (signal_887) ) ;
    buf_clk cell_488 ( .C (clk), .D (signal_892), .Q (signal_893) ) ;
    buf_clk cell_494 ( .C (clk), .D (signal_898), .Q (signal_899) ) ;
    buf_clk cell_500 ( .C (clk), .D (signal_904), .Q (signal_905) ) ;
    buf_clk cell_506 ( .C (clk), .D (signal_910), .Q (signal_911) ) ;
    buf_clk cell_512 ( .C (clk), .D (signal_916), .Q (signal_917) ) ;
    buf_clk cell_518 ( .C (clk), .D (signal_922), .Q (signal_923) ) ;
    buf_clk cell_524 ( .C (clk), .D (signal_928), .Q (signal_929) ) ;
    buf_clk cell_530 ( .C (clk), .D (signal_934), .Q (signal_935) ) ;
    buf_clk cell_536 ( .C (clk), .D (signal_940), .Q (signal_941) ) ;
    buf_clk cell_542 ( .C (clk), .D (signal_946), .Q (signal_947) ) ;
    buf_clk cell_548 ( .C (clk), .D (signal_952), .Q (signal_953) ) ;
    buf_clk cell_554 ( .C (clk), .D (signal_958), .Q (signal_959) ) ;
    buf_clk cell_560 ( .C (clk), .D (signal_964), .Q (signal_965) ) ;
    buf_clk cell_566 ( .C (clk), .D (signal_970), .Q (signal_971) ) ;
    buf_clk cell_572 ( .C (clk), .D (signal_976), .Q (signal_977) ) ;
    buf_clk cell_578 ( .C (clk), .D (signal_982), .Q (signal_983) ) ;
    buf_clk cell_584 ( .C (clk), .D (signal_988), .Q (signal_989) ) ;
    buf_clk cell_590 ( .C (clk), .D (signal_994), .Q (signal_995) ) ;
    buf_clk cell_596 ( .C (clk), .D (signal_1000), .Q (signal_1001) ) ;
    buf_clk cell_602 ( .C (clk), .D (signal_1006), .Q (signal_1007) ) ;
    buf_clk cell_608 ( .C (clk), .D (signal_1012), .Q (signal_1013) ) ;
    buf_clk cell_614 ( .C (clk), .D (signal_1018), .Q (signal_1019) ) ;
    buf_clk cell_620 ( .C (clk), .D (signal_1024), .Q (signal_1025) ) ;
    buf_clk cell_626 ( .C (clk), .D (signal_1030), .Q (signal_1031) ) ;
    buf_clk cell_632 ( .C (clk), .D (signal_1036), .Q (signal_1037) ) ;
    buf_clk cell_638 ( .C (clk), .D (signal_1042), .Q (signal_1043) ) ;
    buf_clk cell_644 ( .C (clk), .D (signal_1048), .Q (signal_1049) ) ;
    buf_clk cell_650 ( .C (clk), .D (signal_1054), .Q (signal_1055) ) ;
    buf_clk cell_656 ( .C (clk), .D (signal_1060), .Q (signal_1061) ) ;
    buf_clk cell_662 ( .C (clk), .D (signal_1066), .Q (signal_1067) ) ;

    /* cells in depth 6 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_194 ( .a ({signal_714, signal_712, signal_710}), .b ({signal_404, signal_403, signal_207}), .clk (clk), .r ({Fresh[38], Fresh[37], Fresh[36]}), .c ({signal_408, signal_407, signal_209}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_195 ( .a ({signal_720, signal_718, signal_716}), .b ({signal_402, signal_401, signal_206}), .clk (clk), .r ({Fresh[41], Fresh[40], Fresh[39]}), .c ({signal_410, signal_409, signal_210}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_196 ( .a ({signal_714, signal_712, signal_710}), .b ({signal_398, signal_397, signal_204}), .clk (clk), .r ({Fresh[44], Fresh[43], Fresh[42]}), .c ({signal_412, signal_411, signal_211}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_197 ( .a ({signal_392, signal_391, signal_201}), .b ({signal_720, signal_718, signal_716}), .clk (clk), .r ({Fresh[47], Fresh[46], Fresh[45]}), .c ({signal_414, signal_413, signal_212}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_199 ( .a ({signal_726, signal_724, signal_722}), .b ({signal_408, signal_407, signal_209}), .c ({signal_418, signal_417, signal_214}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_200 ( .a ({signal_732, signal_730, signal_728}), .b ({signal_412, signal_411, signal_211}), .c ({signal_420, signal_419, signal_215}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_201 ( .a ({signal_738, signal_736, signal_734}), .b ({signal_410, signal_409, signal_210}), .c ({signal_422, signal_421, signal_216}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_202 ( .a ({signal_414, signal_413, signal_212}), .b ({signal_744, signal_742, signal_740}), .c ({signal_424, signal_423, signal_217}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_211 ( .a ({signal_420, signal_419, signal_215}), .b ({signal_424, signal_423, signal_217}), .c ({signal_442, signal_441, signal_226}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_212 ( .a ({signal_418, signal_417, signal_214}), .b ({signal_422, signal_421, signal_216}), .c ({signal_444, signal_443, signal_227}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_213 ( .a ({signal_418, signal_417, signal_214}), .b ({signal_420, signal_419, signal_215}), .c ({signal_446, signal_445, signal_228}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_214 ( .a ({signal_422, signal_421, signal_216}), .b ({signal_424, signal_423, signal_217}), .c ({signal_448, signal_447, signal_229}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_223 ( .a ({signal_442, signal_441, signal_226}), .b ({signal_444, signal_443, signal_227}), .c ({signal_466, signal_465, signal_238}) ) ;
    buf_clk cell_317 ( .C (clk), .D (signal_721), .Q (signal_722) ) ;
    buf_clk cell_319 ( .C (clk), .D (signal_723), .Q (signal_724) ) ;
    buf_clk cell_321 ( .C (clk), .D (signal_725), .Q (signal_726) ) ;
    buf_clk cell_323 ( .C (clk), .D (signal_727), .Q (signal_728) ) ;
    buf_clk cell_325 ( .C (clk), .D (signal_729), .Q (signal_730) ) ;
    buf_clk cell_327 ( .C (clk), .D (signal_731), .Q (signal_732) ) ;
    buf_clk cell_329 ( .C (clk), .D (signal_733), .Q (signal_734) ) ;
    buf_clk cell_331 ( .C (clk), .D (signal_735), .Q (signal_736) ) ;
    buf_clk cell_333 ( .C (clk), .D (signal_737), .Q (signal_738) ) ;
    buf_clk cell_335 ( .C (clk), .D (signal_739), .Q (signal_740) ) ;
    buf_clk cell_337 ( .C (clk), .D (signal_741), .Q (signal_742) ) ;
    buf_clk cell_339 ( .C (clk), .D (signal_743), .Q (signal_744) ) ;
    buf_clk cell_345 ( .C (clk), .D (signal_749), .Q (signal_750) ) ;
    buf_clk cell_351 ( .C (clk), .D (signal_755), .Q (signal_756) ) ;
    buf_clk cell_357 ( .C (clk), .D (signal_761), .Q (signal_762) ) ;
    buf_clk cell_363 ( .C (clk), .D (signal_767), .Q (signal_768) ) ;
    buf_clk cell_369 ( .C (clk), .D (signal_773), .Q (signal_774) ) ;
    buf_clk cell_375 ( .C (clk), .D (signal_779), .Q (signal_780) ) ;
    buf_clk cell_381 ( .C (clk), .D (signal_785), .Q (signal_786) ) ;
    buf_clk cell_387 ( .C (clk), .D (signal_791), .Q (signal_792) ) ;
    buf_clk cell_393 ( .C (clk), .D (signal_797), .Q (signal_798) ) ;
    buf_clk cell_399 ( .C (clk), .D (signal_803), .Q (signal_804) ) ;
    buf_clk cell_405 ( .C (clk), .D (signal_809), .Q (signal_810) ) ;
    buf_clk cell_411 ( .C (clk), .D (signal_815), .Q (signal_816) ) ;
    buf_clk cell_417 ( .C (clk), .D (signal_821), .Q (signal_822) ) ;
    buf_clk cell_423 ( .C (clk), .D (signal_827), .Q (signal_828) ) ;
    buf_clk cell_429 ( .C (clk), .D (signal_833), .Q (signal_834) ) ;
    buf_clk cell_435 ( .C (clk), .D (signal_839), .Q (signal_840) ) ;
    buf_clk cell_441 ( .C (clk), .D (signal_845), .Q (signal_846) ) ;
    buf_clk cell_447 ( .C (clk), .D (signal_851), .Q (signal_852) ) ;
    buf_clk cell_453 ( .C (clk), .D (signal_857), .Q (signal_858) ) ;
    buf_clk cell_459 ( .C (clk), .D (signal_863), .Q (signal_864) ) ;
    buf_clk cell_465 ( .C (clk), .D (signal_869), .Q (signal_870) ) ;
    buf_clk cell_471 ( .C (clk), .D (signal_875), .Q (signal_876) ) ;
    buf_clk cell_477 ( .C (clk), .D (signal_881), .Q (signal_882) ) ;
    buf_clk cell_483 ( .C (clk), .D (signal_887), .Q (signal_888) ) ;
    buf_clk cell_489 ( .C (clk), .D (signal_893), .Q (signal_894) ) ;
    buf_clk cell_495 ( .C (clk), .D (signal_899), .Q (signal_900) ) ;
    buf_clk cell_501 ( .C (clk), .D (signal_905), .Q (signal_906) ) ;
    buf_clk cell_507 ( .C (clk), .D (signal_911), .Q (signal_912) ) ;
    buf_clk cell_513 ( .C (clk), .D (signal_917), .Q (signal_918) ) ;
    buf_clk cell_519 ( .C (clk), .D (signal_923), .Q (signal_924) ) ;
    buf_clk cell_525 ( .C (clk), .D (signal_929), .Q (signal_930) ) ;
    buf_clk cell_531 ( .C (clk), .D (signal_935), .Q (signal_936) ) ;
    buf_clk cell_537 ( .C (clk), .D (signal_941), .Q (signal_942) ) ;
    buf_clk cell_543 ( .C (clk), .D (signal_947), .Q (signal_948) ) ;
    buf_clk cell_549 ( .C (clk), .D (signal_953), .Q (signal_954) ) ;
    buf_clk cell_555 ( .C (clk), .D (signal_959), .Q (signal_960) ) ;
    buf_clk cell_561 ( .C (clk), .D (signal_965), .Q (signal_966) ) ;
    buf_clk cell_567 ( .C (clk), .D (signal_971), .Q (signal_972) ) ;
    buf_clk cell_573 ( .C (clk), .D (signal_977), .Q (signal_978) ) ;
    buf_clk cell_579 ( .C (clk), .D (signal_983), .Q (signal_984) ) ;
    buf_clk cell_585 ( .C (clk), .D (signal_989), .Q (signal_990) ) ;
    buf_clk cell_591 ( .C (clk), .D (signal_995), .Q (signal_996) ) ;
    buf_clk cell_597 ( .C (clk), .D (signal_1001), .Q (signal_1002) ) ;
    buf_clk cell_603 ( .C (clk), .D (signal_1007), .Q (signal_1008) ) ;
    buf_clk cell_609 ( .C (clk), .D (signal_1013), .Q (signal_1014) ) ;
    buf_clk cell_615 ( .C (clk), .D (signal_1019), .Q (signal_1020) ) ;
    buf_clk cell_621 ( .C (clk), .D (signal_1025), .Q (signal_1026) ) ;
    buf_clk cell_627 ( .C (clk), .D (signal_1031), .Q (signal_1032) ) ;
    buf_clk cell_633 ( .C (clk), .D (signal_1037), .Q (signal_1038) ) ;
    buf_clk cell_639 ( .C (clk), .D (signal_1043), .Q (signal_1044) ) ;
    buf_clk cell_645 ( .C (clk), .D (signal_1049), .Q (signal_1050) ) ;
    buf_clk cell_651 ( .C (clk), .D (signal_1055), .Q (signal_1056) ) ;
    buf_clk cell_657 ( .C (clk), .D (signal_1061), .Q (signal_1062) ) ;
    buf_clk cell_663 ( .C (clk), .D (signal_1067), .Q (signal_1068) ) ;

    /* cells in depth 7 */

    /* cells in depth 8 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_203 ( .a ({signal_762, signal_756, signal_750}), .b ({signal_424, signal_423, signal_217}), .clk (clk), .r ({Fresh[50], Fresh[49], Fresh[48]}), .c ({signal_426, signal_425, signal_218}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_204 ( .a ({signal_780, signal_774, signal_768}), .b ({signal_422, signal_421, signal_216}), .clk (clk), .r ({Fresh[53], Fresh[52], Fresh[51]}), .c ({signal_428, signal_427, signal_219}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_205 ( .a ({signal_798, signal_792, signal_786}), .b ({signal_420, signal_419, signal_215}), .clk (clk), .r ({Fresh[56], Fresh[55], Fresh[54]}), .c ({signal_430, signal_429, signal_220}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_206 ( .a ({signal_816, signal_810, signal_804}), .b ({signal_418, signal_417, signal_214}), .clk (clk), .r ({Fresh[59], Fresh[58], Fresh[57]}), .c ({signal_432, signal_431, signal_221}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_207 ( .a ({signal_834, signal_828, signal_822}), .b ({signal_424, signal_423, signal_217}), .clk (clk), .r ({Fresh[62], Fresh[61], Fresh[60]}), .c ({signal_434, signal_433, signal_222}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_208 ( .a ({signal_852, signal_846, signal_840}), .b ({signal_422, signal_421, signal_216}), .clk (clk), .r ({Fresh[65], Fresh[64], Fresh[63]}), .c ({signal_436, signal_435, signal_223}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_209 ( .a ({signal_870, signal_864, signal_858}), .b ({signal_420, signal_419, signal_215}), .clk (clk), .r ({Fresh[68], Fresh[67], Fresh[66]}), .c ({signal_438, signal_437, signal_224}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_210 ( .a ({signal_888, signal_882, signal_876}), .b ({signal_418, signal_417, signal_214}), .clk (clk), .r ({Fresh[71], Fresh[70], Fresh[69]}), .c ({signal_440, signal_439, signal_225}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_215 ( .a ({signal_906, signal_900, signal_894}), .b ({signal_448, signal_447, signal_229}), .clk (clk), .r ({Fresh[74], Fresh[73], Fresh[72]}), .c ({signal_450, signal_449, signal_230}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_216 ( .a ({signal_924, signal_918, signal_912}), .b ({signal_446, signal_445, signal_228}), .clk (clk), .r ({Fresh[77], Fresh[76], Fresh[75]}), .c ({signal_452, signal_451, signal_231}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_217 ( .a ({signal_942, signal_936, signal_930}), .b ({signal_444, signal_443, signal_227}), .clk (clk), .r ({Fresh[80], Fresh[79], Fresh[78]}), .c ({signal_454, signal_453, signal_232}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_218 ( .a ({signal_960, signal_954, signal_948}), .b ({signal_442, signal_441, signal_226}), .clk (clk), .r ({Fresh[83], Fresh[82], Fresh[81]}), .c ({signal_456, signal_455, signal_233}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_219 ( .a ({signal_978, signal_972, signal_966}), .b ({signal_448, signal_447, signal_229}), .clk (clk), .r ({Fresh[86], Fresh[85], Fresh[84]}), .c ({signal_458, signal_457, signal_234}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_220 ( .a ({signal_996, signal_990, signal_984}), .b ({signal_446, signal_445, signal_228}), .clk (clk), .r ({Fresh[89], Fresh[88], Fresh[87]}), .c ({signal_460, signal_459, signal_235}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_221 ( .a ({signal_1014, signal_1008, signal_1002}), .b ({signal_444, signal_443, signal_227}), .clk (clk), .r ({Fresh[92], Fresh[91], Fresh[90]}), .c ({signal_462, signal_461, signal_236}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_222 ( .a ({signal_1032, signal_1026, signal_1020}), .b ({signal_442, signal_441, signal_226}), .clk (clk), .r ({Fresh[95], Fresh[94], Fresh[93]}), .c ({signal_464, signal_463, signal_237}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_224 ( .a ({signal_430, signal_429, signal_220}), .b ({signal_434, signal_433, signal_222}), .c ({signal_468, signal_467, signal_239}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_225 ( .a ({signal_432, signal_431, signal_221}), .b ({signal_438, signal_437, signal_224}), .c ({signal_470, signal_469, signal_240}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_226 ( .a ({signal_428, signal_427, signal_219}), .b ({signal_432, signal_431, signal_221}), .c ({signal_472, signal_471, signal_241}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_227 ( .a ({signal_1050, signal_1044, signal_1038}), .b ({signal_466, signal_465, signal_238}), .clk (clk), .r ({Fresh[98], Fresh[97], Fresh[96]}), .c ({signal_474, signal_473, signal_242}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_228 ( .a ({signal_1068, signal_1062, signal_1056}), .b ({signal_466, signal_465, signal_238}), .clk (clk), .r ({Fresh[101], Fresh[100], Fresh[99]}), .c ({signal_476, signal_475, signal_243}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_229 ( .a ({signal_428, signal_427, signal_219}), .b ({signal_450, signal_449, signal_230}), .c ({signal_478, signal_477, signal_244}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_230 ( .a ({signal_426, signal_425, signal_218}), .b ({signal_458, signal_457, signal_234}), .c ({signal_480, signal_479, signal_245}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_231 ( .a ({signal_456, signal_455, signal_233}), .b ({signal_460, signal_459, signal_235}), .c ({signal_482, signal_481, signal_246}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_232 ( .a ({signal_452, signal_451, signal_231}), .b ({signal_462, signal_461, signal_236}), .c ({signal_484, signal_483, signal_247}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_233 ( .a ({signal_454, signal_453, signal_232}), .b ({signal_462, signal_461, signal_236}), .c ({signal_486, signal_485, signal_248}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_234 ( .a ({signal_458, signal_457, signal_234}), .b ({signal_468, signal_467, signal_239}), .c ({signal_488, signal_487, signal_249}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_235 ( .a ({signal_436, signal_435, signal_223}), .b ({signal_468, signal_467, signal_239}), .c ({signal_490, signal_489, signal_250}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_236 ( .a ({signal_460, signal_459, signal_235}), .b ({signal_470, signal_469, signal_240}), .c ({signal_492, signal_491, signal_251}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_237 ( .a ({signal_462, signal_461, signal_236}), .b ({signal_476, signal_475, signal_243}), .c ({signal_494, signal_493, signal_252}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_238 ( .a ({signal_476, signal_475, signal_243}), .b ({signal_484, signal_483, signal_247}), .c ({signal_496, signal_495, signal_253}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_239 ( .a ({signal_450, signal_449, signal_230}), .b ({signal_480, signal_479, signal_245}), .c ({signal_498, signal_497, signal_254}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_240 ( .a ({signal_454, signal_453, signal_232}), .b ({signal_474, signal_473, signal_242}), .c ({signal_500, signal_499, signal_255}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_241 ( .a ({signal_474, signal_473, signal_242}), .b ({signal_482, signal_481, signal_246}), .c ({signal_502, signal_501, signal_256}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_242 ( .a ({signal_440, signal_439, signal_225}), .b ({signal_478, signal_477, signal_244}), .c ({signal_504, signal_503, signal_257}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_243 ( .a ({signal_464, signal_463, signal_237}), .b ({signal_482, signal_481, signal_246}), .c ({signal_506, signal_505, signal_258}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_244 ( .a ({signal_472, signal_471, signal_241}), .b ({signal_480, signal_479, signal_245}), .c ({signal_508, signal_507, signal_259}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_245 ( .a ({signal_478, signal_477, signal_244}), .b ({signal_492, signal_491, signal_251}), .c ({signal_510, signal_509, signal_260}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_246 ( .a ({signal_430, signal_429, signal_220}), .b ({signal_494, signal_493, signal_252}), .c ({signal_512, signal_511, signal_261}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_247 ( .a ({signal_434, signal_433, signal_222}), .b ({signal_494, signal_493, signal_252}), .c ({signal_514, signal_513, signal_262}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_248 ( .a ({signal_468, signal_467, signal_239}), .b ({signal_494, signal_493, signal_252}), .c ({signal_516, signal_515, signal_263}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_249 ( .a ({signal_468, signal_467, signal_239}), .b ({signal_498, signal_497, signal_254}), .c ({signal_518, signal_517, signal_264}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_250 ( .a ({signal_488, signal_487, signal_249}), .b ({signal_500, signal_499, signal_255}), .c ({signal_520, signal_519, signal_265}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_251 ( .a ({signal_496, signal_495, signal_253}), .b ({signal_502, signal_501, signal_256}), .c ({signal_522, signal_521, signal_266}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_252 ( .a ({signal_498, signal_497, signal_254}), .b ({signal_500, signal_499, signal_255}), .c ({signal_524, signal_523, signal_267}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_253 ( .a ({signal_470, signal_469, signal_240}), .b ({signal_502, signal_501, signal_256}), .c ({signal_526, signal_525, signal_268}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_254 ( .a ({signal_486, signal_485, signal_248}), .b ({signal_504, signal_503, signal_257}), .c ({signal_528, signal_527, signal_269}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_255 ( .a ({signal_490, signal_489, signal_250}), .b ({signal_504, signal_503, signal_257}), .c ({signal_530, signal_529, signal_270}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_256 ( .a ({signal_496, signal_495, signal_253}), .b ({signal_510, signal_509, signal_260}), .c ({signal_532, signal_531, signal_271}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_257 ( .a ({signal_532, signal_531, signal_271}), .b ({signal_534, signal_533, signal_150}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_258 ( .a ({signal_496, signal_495, signal_253}), .b ({signal_520, signal_519, signal_265}), .c ({signal_536, signal_535, signal_143}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_259 ( .a ({signal_514, signal_513, signal_262}), .b ({signal_524, signal_523, signal_267}), .c ({signal_538, signal_537, signal_272}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_260 ( .a ({signal_506, signal_505, signal_258}), .b ({signal_528, signal_527, signal_269}), .c ({signal_540, signal_539, signal_273}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_261 ( .a ({signal_496, signal_495, signal_253}), .b ({signal_518, signal_517, signal_264}), .c ({signal_542, signal_541, signal_146}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_262 ( .a ({signal_508, signal_507, signal_259}), .b ({signal_516, signal_515, signal_263}), .c ({signal_544, signal_543, signal_147}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_263 ( .a ({signal_522, signal_521, signal_266}), .b ({signal_530, signal_529, signal_270}), .c ({signal_546, signal_545, signal_148}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_264 ( .a ({signal_512, signal_511, signal_261}), .b ({signal_526, signal_525, signal_268}), .c ({signal_548, signal_547, signal_274}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_265 ( .a ({signal_538, signal_537, signal_272}), .b ({signal_550, signal_549, signal_144}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_266 ( .a ({signal_540, signal_539, signal_273}), .b ({signal_552, signal_551, signal_145}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_267 ( .a ({signal_548, signal_547, signal_274}), .b ({signal_554, signal_553, signal_149}) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_536, signal_535, signal_143}), .Q ({Y_s2[7], Y_s1[7], Y_s0[7]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_550, signal_549, signal_144}), .Q ({Y_s2[6], Y_s1[6], Y_s0[6]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_552, signal_551, signal_145}), .Q ({Y_s2[5], Y_s1[5], Y_s0[5]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_542, signal_541, signal_146}), .Q ({Y_s2[4], Y_s1[4], Y_s0[4]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_4 ( .clk (clk), .D ({signal_544, signal_543, signal_147}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_5 ( .clk (clk), .D ({signal_546, signal_545, signal_148}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_6 ( .clk (clk), .D ({signal_554, signal_553, signal_149}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_7 ( .clk (clk), .D ({signal_534, signal_533, signal_150}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
