/* modified netlist. Source: module sbox in file Designs/SkinnySbox/AGEMA/sbox_opt_correct/sbox.v */
/* 4 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 5 register stage(s) in total */

module sbox_HPC2_AIG_Pipeline_d2 (X_s0, clk, X_s1, X_s2, Fresh, Y_s0, Y_s1, Y_s2);
    input [3:0] X_s0 ;
    input clk ;
    input [3:0] X_s1 ;
    input [3:0] X_s2 ;
    input [11:0] Fresh ;
    output [3:0] Y_s0 ;
    output [3:0] Y_s1 ;
    output [3:0] Y_s2 ;
    wire signal_33 ;
    wire signal_34 ;
    wire signal_35 ;
    wire signal_36 ;
    wire signal_37 ;
    wire signal_38 ;
    wire signal_39 ;
    wire signal_40 ;
    wire signal_41 ;
    wire signal_42 ;
    wire signal_43 ;
    wire signal_44 ;
    wire signal_45 ;
    wire signal_46 ;
    wire signal_47 ;
    wire signal_48 ;
    wire signal_49 ;
    wire signal_50 ;
    wire signal_51 ;
    wire signal_52 ;
    wire signal_53 ;
    wire signal_54 ;
    wire signal_55 ;
    wire signal_56 ;
    wire signal_59 ;
    wire signal_60 ;
    wire signal_63 ;
    wire signal_64 ;
    wire signal_67 ;
    wire signal_68 ;
    wire signal_71 ;
    wire signal_72 ;
    wire signal_73 ;
    wire signal_74 ;
    wire signal_75 ;
    wire signal_76 ;
    wire signal_77 ;
    wire signal_78 ;
    wire signal_79 ;
    wire signal_80 ;
    wire signal_81 ;
    wire signal_82 ;
    wire signal_83 ;
    wire signal_84 ;
    wire signal_85 ;
    wire signal_86 ;
    wire signal_87 ;
    wire signal_88 ;
    wire signal_89 ;
    wire signal_90 ;
    wire signal_91 ;
    wire signal_92 ;
    wire signal_93 ;
    wire signal_94 ;
    wire signal_95 ;
    wire signal_96 ;
    wire signal_97 ;
    wire signal_98 ;
    wire signal_99 ;
    wire signal_100 ;
    wire signal_101 ;
    wire signal_102 ;
    wire signal_103 ;
    wire signal_104 ;
    wire signal_105 ;
    wire signal_106 ;
    wire signal_107 ;
    wire signal_108 ;
    wire signal_109 ;
    wire signal_110 ;
    wire signal_111 ;
    wire signal_112 ;
    wire signal_133 ;
    wire signal_134 ;
    wire signal_135 ;
    wire signal_136 ;
    wire signal_137 ;
    wire signal_138 ;
    wire signal_139 ;
    wire signal_140 ;
    wire signal_141 ;
    wire signal_142 ;
    wire signal_143 ;
    wire signal_144 ;
    wire signal_145 ;
    wire signal_146 ;
    wire signal_147 ;
    wire signal_148 ;
    wire signal_149 ;
    wire signal_150 ;
    wire signal_151 ;
    wire signal_152 ;
    wire signal_153 ;
    wire signal_154 ;
    wire signal_155 ;
    wire signal_156 ;
    wire signal_157 ;
    wire signal_158 ;
    wire signal_159 ;
    wire signal_160 ;
    wire signal_161 ;
    wire signal_162 ;
    wire signal_163 ;
    wire signal_164 ;
    wire signal_165 ;
    wire signal_166 ;
    wire signal_167 ;
    wire signal_168 ;
    wire signal_169 ;
    wire signal_170 ;
    wire signal_171 ;
    wire signal_172 ;
    wire signal_173 ;
    wire signal_174 ;
    wire signal_175 ;
    wire signal_176 ;
    wire signal_177 ;
    wire signal_178 ;
    wire signal_179 ;
    wire signal_180 ;
    wire signal_181 ;
    wire signal_182 ;
    wire signal_183 ;
    wire signal_184 ;
    wire signal_185 ;
    wire signal_186 ;
    wire signal_187 ;
    wire signal_188 ;
    wire signal_189 ;
    wire signal_190 ;
    wire signal_191 ;
    wire signal_192 ;
    wire signal_193 ;
    wire signal_194 ;
    wire signal_195 ;
    wire signal_196 ;
    wire signal_197 ;
    wire signal_198 ;
    wire signal_199 ;
    wire signal_200 ;
    wire signal_201 ;
    wire signal_202 ;
    wire signal_203 ;
    wire signal_204 ;

    /* cells in depth 0 */
    not_masked #(.security_order(2), .pipeline(1)) cell_26 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_60, signal_59, signal_37}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_27 ( .a ({X_s2[3], X_s1[3], X_s0[3]}), .b ({X_s2[2], X_s1[2], X_s0[2]}), .c ({signal_64, signal_63, signal_38}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_28 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s2[0], X_s1[0], X_s0[0]}), .c ({signal_68, signal_67, signal_39}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_29 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({X_s2[1], X_s1[1], X_s0[1]}), .c ({signal_72, signal_71, signal_40}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_31 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_68, signal_67, signal_39}), .c ({signal_76, signal_75, signal_42}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_32 ( .a ({X_s2[1], X_s1[1], X_s0[1]}), .b ({signal_64, signal_63, signal_38}), .c ({signal_78, signal_77, signal_43}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_33 ( .a ({X_s2[2], X_s1[2], X_s0[2]}), .b ({signal_68, signal_67, signal_39}), .c ({signal_80, signal_79, signal_44}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_34 ( .a ({signal_80, signal_79, signal_44}), .b ({signal_82, signal_81, signal_45}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_36 ( .a ({signal_78, signal_77, signal_43}), .b ({signal_80, signal_79, signal_44}), .c ({signal_86, signal_85, signal_47}) ) ;

    /* cells in depth 1 */
    buf_clk cell_50 ( .C (clk), .D (signal_38), .Q (signal_133) ) ;
    buf_clk cell_52 ( .C (clk), .D (signal_63), .Q (signal_135) ) ;
    buf_clk cell_54 ( .C (clk), .D (signal_64), .Q (signal_137) ) ;
    buf_clk cell_56 ( .C (clk), .D (signal_42), .Q (signal_139) ) ;
    buf_clk cell_58 ( .C (clk), .D (signal_75), .Q (signal_141) ) ;
    buf_clk cell_60 ( .C (clk), .D (signal_76), .Q (signal_143) ) ;
    buf_clk cell_62 ( .C (clk), .D (signal_47), .Q (signal_145) ) ;
    buf_clk cell_64 ( .C (clk), .D (signal_85), .Q (signal_147) ) ;
    buf_clk cell_66 ( .C (clk), .D (signal_86), .Q (signal_149) ) ;
    buf_clk cell_68 ( .C (clk), .D (signal_39), .Q (signal_151) ) ;
    buf_clk cell_70 ( .C (clk), .D (signal_67), .Q (signal_153) ) ;
    buf_clk cell_72 ( .C (clk), .D (signal_68), .Q (signal_155) ) ;
    buf_clk cell_74 ( .C (clk), .D (X_s0[1]), .Q (signal_157) ) ;
    buf_clk cell_76 ( .C (clk), .D (X_s1[1]), .Q (signal_159) ) ;
    buf_clk cell_78 ( .C (clk), .D (X_s2[1]), .Q (signal_161) ) ;
    buf_clk cell_80 ( .C (clk), .D (signal_45), .Q (signal_163) ) ;
    buf_clk cell_82 ( .C (clk), .D (signal_81), .Q (signal_165) ) ;
    buf_clk cell_84 ( .C (clk), .D (signal_82), .Q (signal_167) ) ;
    buf_clk cell_92 ( .C (clk), .D (signal_40), .Q (signal_175) ) ;
    buf_clk cell_96 ( .C (clk), .D (signal_71), .Q (signal_179) ) ;
    buf_clk cell_100 ( .C (clk), .D (signal_72), .Q (signal_183) ) ;

    /* cells in depth 2 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_30 ( .a ({signal_60, signal_59, signal_37}), .b ({signal_72, signal_71, signal_40}), .clk (clk), .r ({Fresh[2], Fresh[1], Fresh[0]}), .c ({signal_74, signal_73, signal_41}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_35 ( .a ({signal_60, signal_59, signal_37}), .b ({signal_78, signal_77, signal_43}), .clk (clk), .r ({Fresh[5], Fresh[4], Fresh[3]}), .c ({signal_84, signal_83, signal_46}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_37 ( .a ({signal_138, signal_136, signal_134}), .b ({signal_74, signal_73, signal_41}), .c ({signal_88, signal_87, signal_48}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_38 ( .a ({signal_88, signal_87, signal_48}), .b ({signal_90, signal_89, signal_36}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_39 ( .a ({signal_144, signal_142, signal_140}), .b ({signal_84, signal_83, signal_46}), .c ({signal_92, signal_91, signal_49}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_40 ( .a ({signal_74, signal_73, signal_41}), .b ({signal_150, signal_148, signal_146}), .c ({signal_94, signal_93, signal_50}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_41 ( .a ({signal_156, signal_154, signal_152}), .b ({signal_84, signal_83, signal_46}), .c ({signal_96, signal_95, signal_51}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_44 ( .a ({signal_74, signal_73, signal_41}), .b ({signal_96, signal_95, signal_51}), .c ({signal_102, signal_101, signal_54}) ) ;
    not_masked #(.security_order(2), .pipeline(1)) cell_45 ( .a ({signal_102, signal_101, signal_54}), .b ({signal_104, signal_103, signal_35}) ) ;
    buf_clk cell_51 ( .C (clk), .D (signal_133), .Q (signal_134) ) ;
    buf_clk cell_53 ( .C (clk), .D (signal_135), .Q (signal_136) ) ;
    buf_clk cell_55 ( .C (clk), .D (signal_137), .Q (signal_138) ) ;
    buf_clk cell_57 ( .C (clk), .D (signal_139), .Q (signal_140) ) ;
    buf_clk cell_59 ( .C (clk), .D (signal_141), .Q (signal_142) ) ;
    buf_clk cell_61 ( .C (clk), .D (signal_143), .Q (signal_144) ) ;
    buf_clk cell_63 ( .C (clk), .D (signal_145), .Q (signal_146) ) ;
    buf_clk cell_65 ( .C (clk), .D (signal_147), .Q (signal_148) ) ;
    buf_clk cell_67 ( .C (clk), .D (signal_149), .Q (signal_150) ) ;
    buf_clk cell_69 ( .C (clk), .D (signal_151), .Q (signal_152) ) ;
    buf_clk cell_71 ( .C (clk), .D (signal_153), .Q (signal_154) ) ;
    buf_clk cell_73 ( .C (clk), .D (signal_155), .Q (signal_156) ) ;
    buf_clk cell_75 ( .C (clk), .D (signal_157), .Q (signal_158) ) ;
    buf_clk cell_77 ( .C (clk), .D (signal_159), .Q (signal_160) ) ;
    buf_clk cell_79 ( .C (clk), .D (signal_161), .Q (signal_162) ) ;
    buf_clk cell_81 ( .C (clk), .D (signal_163), .Q (signal_164) ) ;
    buf_clk cell_83 ( .C (clk), .D (signal_165), .Q (signal_166) ) ;
    buf_clk cell_85 ( .C (clk), .D (signal_167), .Q (signal_168) ) ;
    buf_clk cell_93 ( .C (clk), .D (signal_175), .Q (signal_176) ) ;
    buf_clk cell_97 ( .C (clk), .D (signal_179), .Q (signal_180) ) ;
    buf_clk cell_101 ( .C (clk), .D (signal_183), .Q (signal_184) ) ;

    /* cells in depth 3 */
    buf_clk cell_86 ( .C (clk), .D (signal_41), .Q (signal_169) ) ;
    buf_clk cell_88 ( .C (clk), .D (signal_73), .Q (signal_171) ) ;
    buf_clk cell_90 ( .C (clk), .D (signal_74), .Q (signal_173) ) ;
    buf_clk cell_94 ( .C (clk), .D (signal_176), .Q (signal_177) ) ;
    buf_clk cell_98 ( .C (clk), .D (signal_180), .Q (signal_181) ) ;
    buf_clk cell_102 ( .C (clk), .D (signal_184), .Q (signal_185) ) ;
    buf_clk cell_104 ( .C (clk), .D (signal_51), .Q (signal_187) ) ;
    buf_clk cell_106 ( .C (clk), .D (signal_95), .Q (signal_189) ) ;
    buf_clk cell_108 ( .C (clk), .D (signal_96), .Q (signal_191) ) ;
    buf_clk cell_110 ( .C (clk), .D (signal_35), .Q (signal_193) ) ;
    buf_clk cell_112 ( .C (clk), .D (signal_103), .Q (signal_195) ) ;
    buf_clk cell_114 ( .C (clk), .D (signal_104), .Q (signal_197) ) ;
    buf_clk cell_116 ( .C (clk), .D (signal_36), .Q (signal_199) ) ;
    buf_clk cell_118 ( .C (clk), .D (signal_89), .Q (signal_201) ) ;
    buf_clk cell_120 ( .C (clk), .D (signal_90), .Q (signal_203) ) ;

    /* cells in depth 4 */
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_42 ( .a ({signal_162, signal_160, signal_158}), .b ({signal_92, signal_91, signal_49}), .clk (clk), .r ({Fresh[8], Fresh[7], Fresh[6]}), .c ({signal_98, signal_97, signal_52}) ) ;
    and_HPC2 #(.security_order(2), .pipeline(1)) cell_43 ( .a ({signal_168, signal_166, signal_164}), .b ({signal_94, signal_93, signal_50}), .clk (clk), .r ({Fresh[11], Fresh[10], Fresh[9]}), .c ({signal_100, signal_99, signal_53}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_46 ( .a ({signal_174, signal_172, signal_170}), .b ({signal_98, signal_97, signal_52}), .c ({signal_106, signal_105, signal_55}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_47 ( .a ({signal_186, signal_182, signal_178}), .b ({signal_98, signal_97, signal_52}), .c ({signal_108, signal_107, signal_56}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_48 ( .a ({signal_192, signal_190, signal_188}), .b ({signal_108, signal_107, signal_56}), .c ({signal_110, signal_109, signal_33}) ) ;
    xor_HPC2 #(.security_order(2), .pipeline(1)) cell_49 ( .a ({signal_100, signal_99, signal_53}), .b ({signal_106, signal_105, signal_55}), .c ({signal_112, signal_111, signal_34}) ) ;
    buf_clk cell_87 ( .C (clk), .D (signal_169), .Q (signal_170) ) ;
    buf_clk cell_89 ( .C (clk), .D (signal_171), .Q (signal_172) ) ;
    buf_clk cell_91 ( .C (clk), .D (signal_173), .Q (signal_174) ) ;
    buf_clk cell_95 ( .C (clk), .D (signal_177), .Q (signal_178) ) ;
    buf_clk cell_99 ( .C (clk), .D (signal_181), .Q (signal_182) ) ;
    buf_clk cell_103 ( .C (clk), .D (signal_185), .Q (signal_186) ) ;
    buf_clk cell_105 ( .C (clk), .D (signal_187), .Q (signal_188) ) ;
    buf_clk cell_107 ( .C (clk), .D (signal_189), .Q (signal_190) ) ;
    buf_clk cell_109 ( .C (clk), .D (signal_191), .Q (signal_192) ) ;
    buf_clk cell_111 ( .C (clk), .D (signal_193), .Q (signal_194) ) ;
    buf_clk cell_113 ( .C (clk), .D (signal_195), .Q (signal_196) ) ;
    buf_clk cell_115 ( .C (clk), .D (signal_197), .Q (signal_198) ) ;
    buf_clk cell_117 ( .C (clk), .D (signal_199), .Q (signal_200) ) ;
    buf_clk cell_119 ( .C (clk), .D (signal_201), .Q (signal_202) ) ;
    buf_clk cell_121 ( .C (clk), .D (signal_203), .Q (signal_204) ) ;

    /* register cells */
    reg_masked #(.security_order(2), .pipeline(1)) cell_0 ( .clk (clk), .D ({signal_198, signal_196, signal_194}), .Q ({Y_s2[3], Y_s1[3], Y_s0[3]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_1 ( .clk (clk), .D ({signal_204, signal_202, signal_200}), .Q ({Y_s2[2], Y_s1[2], Y_s0[2]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_2 ( .clk (clk), .D ({signal_110, signal_109, signal_33}), .Q ({Y_s2[1], Y_s1[1], Y_s0[1]}) ) ;
    reg_masked #(.security_order(2), .pipeline(1)) cell_3 ( .clk (clk), .D ({signal_112, signal_111, signal_34}), .Q ({Y_s2[0], Y_s1[0], Y_s0[0]}) ) ;
endmodule
