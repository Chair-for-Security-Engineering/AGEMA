/* modified netlist. Source: module AES in file AES.v */
/* 1 register stage(s) are added to the circuit and formed a pipeline design */
/* the circuit has 2 register stage(s) in total */

module AES_GHPCLL_ANF_Pipeline_d1 (plaintext_s0, key_s0, clk, reset, plaintext_s1, key_s1, Fresh, ciphertext_s0, done, ciphertext_s1);
    input [127:0] plaintext_s0 ;
    input [127:0] key_s0 ;
    input clk ;
    input reset ;
    input [127:0] plaintext_s1 ;
    input [127:0] key_s1 ;
    input [8191:0] Fresh ;
    output [127:0] ciphertext_s0 ;
    output done ;
    output [127:0] ciphertext_s1 ;
    wire signal_393 ;
    wire signal_394 ;
    wire signal_395 ;
    wire signal_396 ;
    wire signal_397 ;
    wire signal_398 ;
    wire signal_399 ;
    wire signal_400 ;
    wire signal_401 ;
    wire signal_402 ;
    wire signal_403 ;
    wire signal_404 ;
    wire signal_405 ;
    wire signal_406 ;
    wire signal_407 ;
    wire signal_408 ;
    wire signal_409 ;
    wire signal_410 ;
    wire signal_411 ;
    wire signal_412 ;
    wire signal_413 ;
    wire signal_414 ;
    wire signal_416 ;
    wire signal_418 ;
    wire signal_420 ;
    wire signal_422 ;
    wire signal_424 ;
    wire signal_426 ;
    wire signal_428 ;
    wire signal_430 ;
    wire signal_432 ;
    wire signal_434 ;
    wire signal_436 ;
    wire signal_438 ;
    wire signal_440 ;
    wire signal_442 ;
    wire signal_444 ;
    wire signal_446 ;
    wire signal_448 ;
    wire signal_450 ;
    wire signal_452 ;
    wire signal_454 ;
    wire signal_456 ;
    wire signal_458 ;
    wire signal_460 ;
    wire signal_462 ;
    wire signal_464 ;
    wire signal_466 ;
    wire signal_468 ;
    wire signal_470 ;
    wire signal_472 ;
    wire signal_474 ;
    wire signal_476 ;
    wire signal_478 ;
    wire signal_480 ;
    wire signal_482 ;
    wire signal_484 ;
    wire signal_486 ;
    wire signal_488 ;
    wire signal_490 ;
    wire signal_492 ;
    wire signal_494 ;
    wire signal_496 ;
    wire signal_498 ;
    wire signal_500 ;
    wire signal_502 ;
    wire signal_504 ;
    wire signal_506 ;
    wire signal_508 ;
    wire signal_510 ;
    wire signal_512 ;
    wire signal_514 ;
    wire signal_516 ;
    wire signal_518 ;
    wire signal_520 ;
    wire signal_522 ;
    wire signal_524 ;
    wire signal_526 ;
    wire signal_528 ;
    wire signal_530 ;
    wire signal_532 ;
    wire signal_534 ;
    wire signal_536 ;
    wire signal_538 ;
    wire signal_540 ;
    wire signal_542 ;
    wire signal_544 ;
    wire signal_546 ;
    wire signal_548 ;
    wire signal_550 ;
    wire signal_552 ;
    wire signal_554 ;
    wire signal_556 ;
    wire signal_558 ;
    wire signal_560 ;
    wire signal_562 ;
    wire signal_564 ;
    wire signal_566 ;
    wire signal_568 ;
    wire signal_570 ;
    wire signal_572 ;
    wire signal_574 ;
    wire signal_576 ;
    wire signal_578 ;
    wire signal_580 ;
    wire signal_582 ;
    wire signal_584 ;
    wire signal_586 ;
    wire signal_588 ;
    wire signal_590 ;
    wire signal_592 ;
    wire signal_594 ;
    wire signal_596 ;
    wire signal_598 ;
    wire signal_600 ;
    wire signal_602 ;
    wire signal_604 ;
    wire signal_606 ;
    wire signal_608 ;
    wire signal_610 ;
    wire signal_612 ;
    wire signal_614 ;
    wire signal_616 ;
    wire signal_618 ;
    wire signal_620 ;
    wire signal_622 ;
    wire signal_624 ;
    wire signal_626 ;
    wire signal_628 ;
    wire signal_630 ;
    wire signal_632 ;
    wire signal_634 ;
    wire signal_636 ;
    wire signal_638 ;
    wire signal_640 ;
    wire signal_642 ;
    wire signal_644 ;
    wire signal_646 ;
    wire signal_648 ;
    wire signal_650 ;
    wire signal_652 ;
    wire signal_654 ;
    wire signal_656 ;
    wire signal_658 ;
    wire signal_660 ;
    wire signal_662 ;
    wire signal_664 ;
    wire signal_666 ;
    wire signal_668 ;
    wire signal_670 ;
    wire signal_671 ;
    wire signal_672 ;
    wire signal_788 ;
    wire signal_908 ;
    wire signal_1028 ;
    wire signal_1148 ;
    wire signal_1153 ;
    wire signal_1216 ;
    wire signal_1217 ;
    wire signal_1218 ;
    wire signal_1219 ;
    wire signal_1220 ;
    wire signal_1221 ;
    wire signal_1222 ;
    wire signal_1223 ;
    wire signal_1224 ;
    wire signal_1225 ;
    wire signal_1226 ;
    wire signal_1227 ;
    wire signal_1229 ;
    wire signal_1231 ;
    wire signal_1233 ;
    wire signal_1235 ;
    wire signal_1237 ;
    wire signal_1239 ;
    wire signal_1241 ;
    wire signal_1243 ;
    wire signal_1245 ;
    wire signal_1247 ;
    wire signal_1249 ;
    wire signal_1251 ;
    wire signal_1253 ;
    wire signal_1255 ;
    wire signal_1257 ;
    wire signal_1259 ;
    wire signal_1261 ;
    wire signal_1263 ;
    wire signal_1265 ;
    wire signal_1267 ;
    wire signal_1269 ;
    wire signal_1271 ;
    wire signal_1273 ;
    wire signal_1275 ;
    wire signal_1277 ;
    wire signal_1279 ;
    wire signal_1281 ;
    wire signal_1283 ;
    wire signal_1285 ;
    wire signal_1287 ;
    wire signal_1289 ;
    wire signal_1291 ;
    wire signal_1293 ;
    wire signal_1295 ;
    wire signal_1297 ;
    wire signal_1299 ;
    wire signal_1301 ;
    wire signal_1303 ;
    wire signal_1305 ;
    wire signal_1307 ;
    wire signal_1309 ;
    wire signal_1311 ;
    wire signal_1313 ;
    wire signal_1315 ;
    wire signal_1317 ;
    wire signal_1319 ;
    wire signal_1321 ;
    wire signal_1323 ;
    wire signal_1325 ;
    wire signal_1327 ;
    wire signal_1329 ;
    wire signal_1331 ;
    wire signal_1333 ;
    wire signal_1335 ;
    wire signal_1337 ;
    wire signal_1339 ;
    wire signal_1341 ;
    wire signal_1343 ;
    wire signal_1345 ;
    wire signal_1347 ;
    wire signal_1349 ;
    wire signal_1351 ;
    wire signal_1353 ;
    wire signal_1355 ;
    wire signal_1357 ;
    wire signal_1359 ;
    wire signal_1361 ;
    wire signal_1363 ;
    wire signal_1365 ;
    wire signal_1367 ;
    wire signal_1369 ;
    wire signal_1371 ;
    wire signal_1373 ;
    wire signal_1375 ;
    wire signal_1377 ;
    wire signal_1379 ;
    wire signal_1381 ;
    wire signal_1383 ;
    wire signal_1385 ;
    wire signal_1387 ;
    wire signal_1389 ;
    wire signal_1391 ;
    wire signal_1393 ;
    wire signal_1395 ;
    wire signal_1397 ;
    wire signal_1399 ;
    wire signal_1401 ;
    wire signal_1403 ;
    wire signal_1405 ;
    wire signal_1407 ;
    wire signal_1409 ;
    wire signal_1411 ;
    wire signal_1413 ;
    wire signal_1415 ;
    wire signal_1417 ;
    wire signal_1419 ;
    wire signal_1421 ;
    wire signal_1423 ;
    wire signal_1425 ;
    wire signal_1427 ;
    wire signal_1429 ;
    wire signal_1431 ;
    wire signal_1433 ;
    wire signal_1435 ;
    wire signal_1437 ;
    wire signal_1439 ;
    wire signal_1441 ;
    wire signal_1443 ;
    wire signal_1445 ;
    wire signal_1447 ;
    wire signal_1449 ;
    wire signal_1451 ;
    wire signal_1453 ;
    wire signal_1455 ;
    wire signal_1457 ;
    wire signal_1459 ;
    wire signal_1461 ;
    wire signal_1463 ;
    wire signal_1465 ;
    wire signal_1467 ;
    wire signal_1469 ;
    wire signal_1471 ;
    wire signal_1473 ;
    wire signal_1475 ;
    wire signal_1477 ;
    wire signal_1479 ;
    wire signal_1481 ;
    wire signal_1483 ;
    wire signal_1484 ;
    wire signal_1485 ;
    wire signal_1486 ;
    wire signal_1487 ;
    wire signal_1488 ;
    wire signal_1489 ;
    wire signal_1490 ;
    wire signal_1491 ;
    wire signal_1492 ;
    wire signal_1493 ;
    wire signal_1494 ;
    wire signal_1495 ;
    wire signal_1496 ;
    wire signal_1497 ;
    wire signal_1498 ;
    wire signal_1499 ;
    wire signal_1500 ;
    wire signal_1501 ;
    wire signal_1502 ;
    wire signal_1506 ;
    wire signal_1507 ;
    wire signal_1508 ;
    wire signal_1509 ;
    wire signal_1510 ;
    wire signal_1511 ;
    wire signal_1512 ;
    wire signal_1513 ;
    wire signal_1514 ;
    wire signal_1515 ;
    wire signal_1516 ;
    wire signal_1517 ;
    wire signal_1518 ;
    wire signal_1519 ;
    wire signal_1520 ;
    wire signal_1522 ;
    wire signal_1523 ;
    wire signal_1524 ;
    wire signal_1525 ;
    wire signal_1526 ;
    wire signal_1527 ;
    wire signal_1528 ;
    wire signal_1529 ;
    wire signal_1530 ;
    wire signal_1531 ;
    wire signal_1532 ;
    wire signal_1533 ;
    wire signal_1534 ;
    wire signal_1535 ;
    wire signal_1536 ;
    wire signal_1537 ;
    wire signal_1538 ;
    wire signal_1539 ;
    wire signal_1540 ;
    wire signal_1541 ;
    wire signal_1542 ;
    wire signal_1543 ;
    wire signal_1544 ;
    wire signal_1545 ;
    wire signal_1546 ;
    wire signal_1547 ;
    wire signal_1548 ;
    wire signal_1549 ;
    wire signal_1550 ;
    wire signal_1551 ;
    wire signal_1552 ;
    wire signal_1553 ;
    wire signal_1554 ;
    wire signal_1555 ;
    wire signal_1556 ;
    wire signal_1557 ;
    wire signal_1558 ;
    wire signal_1559 ;
    wire signal_1560 ;
    wire signal_1561 ;
    wire signal_1562 ;
    wire signal_1563 ;
    wire signal_1564 ;
    wire signal_1565 ;
    wire signal_1566 ;
    wire signal_1567 ;
    wire signal_1568 ;
    wire signal_1569 ;
    wire signal_1570 ;
    wire signal_1571 ;
    wire signal_1572 ;
    wire signal_1573 ;
    wire signal_1574 ;
    wire signal_1575 ;
    wire signal_1576 ;
    wire signal_1577 ;
    wire signal_1578 ;
    wire signal_1579 ;
    wire signal_1580 ;
    wire signal_1581 ;
    wire signal_1582 ;
    wire signal_1583 ;
    wire signal_1584 ;
    wire signal_1585 ;
    wire signal_1586 ;
    wire signal_1587 ;
    wire signal_1588 ;
    wire signal_1589 ;
    wire signal_1590 ;
    wire signal_1591 ;
    wire signal_1592 ;
    wire signal_1593 ;
    wire signal_1594 ;
    wire signal_1595 ;
    wire signal_1596 ;
    wire signal_1597 ;
    wire signal_1598 ;
    wire signal_1599 ;
    wire signal_1600 ;
    wire signal_1601 ;
    wire signal_1602 ;
    wire signal_1603 ;
    wire signal_1604 ;
    wire signal_1605 ;
    wire signal_1606 ;
    wire signal_1607 ;
    wire signal_1608 ;
    wire signal_1609 ;
    wire signal_1610 ;
    wire signal_1611 ;
    wire signal_1612 ;
    wire signal_1613 ;
    wire signal_1614 ;
    wire signal_1615 ;
    wire signal_1616 ;
    wire signal_1617 ;
    wire signal_1618 ;
    wire signal_1619 ;
    wire signal_1620 ;
    wire signal_1621 ;
    wire signal_1622 ;
    wire signal_1623 ;
    wire signal_1624 ;
    wire signal_1625 ;
    wire signal_1626 ;
    wire signal_1627 ;
    wire signal_1628 ;
    wire signal_1629 ;
    wire signal_1630 ;
    wire signal_1631 ;
    wire signal_1632 ;
    wire signal_1633 ;
    wire signal_1634 ;
    wire signal_1635 ;
    wire signal_1636 ;
    wire signal_1637 ;
    wire signal_1638 ;
    wire signal_1639 ;
    wire signal_1640 ;
    wire signal_1641 ;
    wire signal_1642 ;
    wire signal_1643 ;
    wire signal_1644 ;
    wire signal_1645 ;
    wire signal_1646 ;
    wire signal_1647 ;
    wire signal_1648 ;
    wire signal_1649 ;
    wire signal_1650 ;
    wire signal_1651 ;
    wire signal_1652 ;
    wire signal_1653 ;
    wire signal_1654 ;
    wire signal_1655 ;
    wire signal_1656 ;
    wire signal_1657 ;
    wire signal_1658 ;
    wire signal_1659 ;
    wire signal_1660 ;
    wire signal_1661 ;
    wire signal_1662 ;
    wire signal_1663 ;
    wire signal_1664 ;
    wire signal_1665 ;
    wire signal_1666 ;
    wire signal_1667 ;
    wire signal_1668 ;
    wire signal_1669 ;
    wire signal_1670 ;
    wire signal_1671 ;
    wire signal_1672 ;
    wire signal_1673 ;
    wire signal_1674 ;
    wire signal_1675 ;
    wire signal_1676 ;
    wire signal_1677 ;
    wire signal_1678 ;
    wire signal_1679 ;
    wire signal_1680 ;
    wire signal_1681 ;
    wire signal_1682 ;
    wire signal_1683 ;
    wire signal_1684 ;
    wire signal_1685 ;
    wire signal_1686 ;
    wire signal_1687 ;
    wire signal_1688 ;
    wire signal_1689 ;
    wire signal_1690 ;
    wire signal_1691 ;
    wire signal_1692 ;
    wire signal_1693 ;
    wire signal_1694 ;
    wire signal_1695 ;
    wire signal_1696 ;
    wire signal_1697 ;
    wire signal_1698 ;
    wire signal_1699 ;
    wire signal_1700 ;
    wire signal_1701 ;
    wire signal_1702 ;
    wire signal_1703 ;
    wire signal_1704 ;
    wire signal_1705 ;
    wire signal_1706 ;
    wire signal_1707 ;
    wire signal_1708 ;
    wire signal_1709 ;
    wire signal_1710 ;
    wire signal_1711 ;
    wire signal_1712 ;
    wire signal_1713 ;
    wire signal_1714 ;
    wire signal_1715 ;
    wire signal_1716 ;
    wire signal_1717 ;
    wire signal_1718 ;
    wire signal_1719 ;
    wire signal_1720 ;
    wire signal_1721 ;
    wire signal_1722 ;
    wire signal_1723 ;
    wire signal_1724 ;
    wire signal_1725 ;
    wire signal_1726 ;
    wire signal_1727 ;
    wire signal_1728 ;
    wire signal_1729 ;
    wire signal_1730 ;
    wire signal_1731 ;
    wire signal_1732 ;
    wire signal_1733 ;
    wire signal_1734 ;
    wire signal_1735 ;
    wire signal_1736 ;
    wire signal_1737 ;
    wire signal_1738 ;
    wire signal_1739 ;
    wire signal_1740 ;
    wire signal_1741 ;
    wire signal_1742 ;
    wire signal_1743 ;
    wire signal_1744 ;
    wire signal_1745 ;
    wire signal_1746 ;
    wire signal_1747 ;
    wire signal_1748 ;
    wire signal_1749 ;
    wire signal_1750 ;
    wire signal_1751 ;
    wire signal_1752 ;
    wire signal_1753 ;
    wire signal_1754 ;
    wire signal_1755 ;
    wire signal_1756 ;
    wire signal_1757 ;
    wire signal_1758 ;
    wire signal_1759 ;
    wire signal_1760 ;
    wire signal_1761 ;
    wire signal_1762 ;
    wire signal_1763 ;
    wire signal_1764 ;
    wire signal_1765 ;
    wire signal_1766 ;
    wire signal_1767 ;
    wire signal_1768 ;
    wire signal_1769 ;
    wire signal_1770 ;
    wire signal_1771 ;
    wire signal_1772 ;
    wire signal_1773 ;
    wire signal_1774 ;
    wire signal_1775 ;
    wire signal_1776 ;
    wire signal_1777 ;
    wire signal_1778 ;
    wire signal_1779 ;
    wire signal_1780 ;
    wire signal_1781 ;
    wire signal_1782 ;
    wire signal_1783 ;
    wire signal_1784 ;
    wire signal_1785 ;
    wire signal_1786 ;
    wire signal_1787 ;
    wire signal_1788 ;
    wire signal_1789 ;
    wire signal_1790 ;
    wire signal_1791 ;
    wire signal_1792 ;
    wire signal_1793 ;
    wire signal_1794 ;
    wire signal_1795 ;
    wire signal_1796 ;
    wire signal_1797 ;
    wire signal_1798 ;
    wire signal_1799 ;
    wire signal_1800 ;
    wire signal_1801 ;
    wire signal_1802 ;
    wire signal_1803 ;
    wire signal_1804 ;
    wire signal_1805 ;
    wire signal_1806 ;
    wire signal_1807 ;
    wire signal_1808 ;
    wire signal_1809 ;
    wire signal_1810 ;
    wire signal_1811 ;
    wire signal_1812 ;
    wire signal_1813 ;
    wire signal_1814 ;
    wire signal_1815 ;
    wire signal_1816 ;
    wire signal_1817 ;
    wire signal_1818 ;
    wire signal_1819 ;
    wire signal_1820 ;
    wire signal_1821 ;
    wire signal_1822 ;
    wire signal_1823 ;
    wire signal_1824 ;
    wire signal_1825 ;
    wire signal_1826 ;
    wire signal_1827 ;
    wire signal_1828 ;
    wire signal_1829 ;
    wire signal_1830 ;
    wire signal_1831 ;
    wire signal_1832 ;
    wire signal_1833 ;
    wire signal_1834 ;
    wire signal_1835 ;
    wire signal_1836 ;
    wire signal_1837 ;
    wire signal_1838 ;
    wire signal_1839 ;
    wire signal_1840 ;
    wire signal_1841 ;
    wire signal_1842 ;
    wire signal_1843 ;
    wire signal_1845 ;
    wire signal_1846 ;
    wire signal_1847 ;
    wire signal_1848 ;
    wire signal_1849 ;
    wire signal_1850 ;
    wire signal_1851 ;
    wire signal_1852 ;
    wire signal_1853 ;
    wire signal_1854 ;
    wire signal_1855 ;
    wire signal_1856 ;
    wire signal_1857 ;
    wire signal_1858 ;
    wire signal_1859 ;
    wire signal_1860 ;
    wire signal_1861 ;
    wire signal_1862 ;
    wire signal_1863 ;
    wire signal_1864 ;
    wire signal_1865 ;
    wire signal_1866 ;
    wire signal_1867 ;
    wire signal_1868 ;
    wire signal_1869 ;
    wire signal_1870 ;
    wire signal_1871 ;
    wire signal_1872 ;
    wire signal_1873 ;
    wire signal_1874 ;
    wire signal_1875 ;
    wire signal_1876 ;
    wire signal_1877 ;
    wire signal_1878 ;
    wire signal_1879 ;
    wire signal_1880 ;
    wire signal_1881 ;
    wire signal_1882 ;
    wire signal_1883 ;
    wire signal_1884 ;
    wire signal_1885 ;
    wire signal_1886 ;
    wire signal_1887 ;
    wire signal_1888 ;
    wire signal_1889 ;
    wire signal_1890 ;
    wire signal_1891 ;
    wire signal_1892 ;
    wire signal_1893 ;
    wire signal_1894 ;
    wire signal_1895 ;
    wire signal_1896 ;
    wire signal_1897 ;
    wire signal_1898 ;
    wire signal_1899 ;
    wire signal_1900 ;
    wire signal_1901 ;
    wire signal_1902 ;
    wire signal_1903 ;
    wire signal_1904 ;
    wire signal_1905 ;
    wire signal_1906 ;
    wire signal_1907 ;
    wire signal_1908 ;
    wire signal_1909 ;
    wire signal_1910 ;
    wire signal_1911 ;
    wire signal_1912 ;
    wire signal_1913 ;
    wire signal_1914 ;
    wire signal_1915 ;
    wire signal_1916 ;
    wire signal_1917 ;
    wire signal_1918 ;
    wire signal_1919 ;
    wire signal_1920 ;
    wire signal_1921 ;
    wire signal_1922 ;
    wire signal_1923 ;
    wire signal_1924 ;
    wire signal_1925 ;
    wire signal_1926 ;
    wire signal_1927 ;
    wire signal_1928 ;
    wire signal_1929 ;
    wire signal_1930 ;
    wire signal_1931 ;
    wire signal_1932 ;
    wire signal_1933 ;
    wire signal_1934 ;
    wire signal_1935 ;
    wire signal_1936 ;
    wire signal_1937 ;
    wire signal_1938 ;
    wire signal_1939 ;
    wire signal_1940 ;
    wire signal_1941 ;
    wire signal_1942 ;
    wire signal_1943 ;
    wire signal_1944 ;
    wire signal_1945 ;
    wire signal_1946 ;
    wire signal_1947 ;
    wire signal_1948 ;
    wire signal_1949 ;
    wire signal_1950 ;
    wire signal_1951 ;
    wire signal_1952 ;
    wire signal_1953 ;
    wire signal_1954 ;
    wire signal_1955 ;
    wire signal_1956 ;
    wire signal_1957 ;
    wire signal_1958 ;
    wire signal_1959 ;
    wire signal_1960 ;
    wire signal_1961 ;
    wire signal_1962 ;
    wire signal_1963 ;
    wire signal_1964 ;
    wire signal_1965 ;
    wire signal_1966 ;
    wire signal_1967 ;
    wire signal_1968 ;
    wire signal_1969 ;
    wire signal_1970 ;
    wire signal_1971 ;
    wire signal_1972 ;
    wire signal_1973 ;
    wire signal_1974 ;
    wire signal_1975 ;
    wire signal_1976 ;
    wire signal_1977 ;
    wire signal_1978 ;
    wire signal_1979 ;
    wire signal_1980 ;
    wire signal_1981 ;
    wire signal_1982 ;
    wire signal_1983 ;
    wire signal_1984 ;
    wire signal_1985 ;
    wire signal_1986 ;
    wire signal_1987 ;
    wire signal_1988 ;
    wire signal_1989 ;
    wire signal_1990 ;
    wire signal_1991 ;
    wire signal_1992 ;
    wire signal_1993 ;
    wire signal_1994 ;
    wire signal_1995 ;
    wire signal_1996 ;
    wire signal_1997 ;
    wire signal_1998 ;
    wire signal_1999 ;
    wire signal_2000 ;
    wire signal_2001 ;
    wire signal_2002 ;
    wire signal_2003 ;
    wire signal_2004 ;
    wire signal_2005 ;
    wire signal_2006 ;
    wire signal_2007 ;
    wire signal_2008 ;
    wire signal_2009 ;
    wire signal_2010 ;
    wire signal_2011 ;
    wire signal_2012 ;
    wire signal_2013 ;
    wire signal_2014 ;
    wire signal_2015 ;
    wire signal_2016 ;
    wire signal_2017 ;
    wire signal_2018 ;
    wire signal_2019 ;
    wire signal_2020 ;
    wire signal_2021 ;
    wire signal_2022 ;
    wire signal_2023 ;
    wire signal_2024 ;
    wire signal_2025 ;
    wire signal_2026 ;
    wire signal_2027 ;
    wire signal_2028 ;
    wire signal_2029 ;
    wire signal_2030 ;
    wire signal_2031 ;
    wire signal_2032 ;
    wire signal_2033 ;
    wire signal_2034 ;
    wire signal_2035 ;
    wire signal_2036 ;
    wire signal_2037 ;
    wire signal_2038 ;
    wire signal_2039 ;
    wire signal_2040 ;
    wire signal_2041 ;
    wire signal_2042 ;
    wire signal_2043 ;
    wire signal_2044 ;
    wire signal_2045 ;
    wire signal_2046 ;
    wire signal_2047 ;
    wire signal_2048 ;
    wire signal_2049 ;
    wire signal_2050 ;
    wire signal_2051 ;
    wire signal_2052 ;
    wire signal_2053 ;
    wire signal_2054 ;
    wire signal_2055 ;
    wire signal_2056 ;
    wire signal_2057 ;
    wire signal_2058 ;
    wire signal_2059 ;
    wire signal_2060 ;
    wire signal_2061 ;
    wire signal_2062 ;
    wire signal_2063 ;
    wire signal_2064 ;
    wire signal_2065 ;
    wire signal_2066 ;
    wire signal_2067 ;
    wire signal_2068 ;
    wire signal_2069 ;
    wire signal_2070 ;
    wire signal_2071 ;
    wire signal_2072 ;
    wire signal_2073 ;
    wire signal_2074 ;
    wire signal_2075 ;
    wire signal_2076 ;
    wire signal_2077 ;
    wire signal_2078 ;
    wire signal_2079 ;
    wire signal_2080 ;
    wire signal_2081 ;
    wire signal_2082 ;
    wire signal_2083 ;
    wire signal_2084 ;
    wire signal_2085 ;
    wire signal_2086 ;
    wire signal_2087 ;
    wire signal_2088 ;
    wire signal_2089 ;
    wire signal_2090 ;
    wire signal_2091 ;
    wire signal_2092 ;
    wire signal_2093 ;
    wire signal_2094 ;
    wire signal_2095 ;
    wire signal_2096 ;
    wire signal_2097 ;
    wire signal_2098 ;
    wire signal_2099 ;
    wire signal_2100 ;
    wire signal_2101 ;
    wire signal_2102 ;
    wire signal_2103 ;
    wire signal_2104 ;
    wire signal_2105 ;
    wire signal_2106 ;
    wire signal_2107 ;
    wire signal_2108 ;
    wire signal_2109 ;
    wire signal_2110 ;
    wire signal_2111 ;
    wire signal_2112 ;
    wire signal_2113 ;
    wire signal_2114 ;
    wire signal_2115 ;
    wire signal_2116 ;
    wire signal_2117 ;
    wire signal_2118 ;
    wire signal_2119 ;
    wire signal_2120 ;
    wire signal_2121 ;
    wire signal_2122 ;
    wire signal_2123 ;
    wire signal_2124 ;
    wire signal_2125 ;
    wire signal_2126 ;
    wire signal_2127 ;
    wire signal_2128 ;
    wire signal_2129 ;
    wire signal_2130 ;
    wire signal_2131 ;
    wire signal_2132 ;
    wire signal_2133 ;
    wire signal_2134 ;
    wire signal_2135 ;
    wire signal_2136 ;
    wire signal_2137 ;
    wire signal_2138 ;
    wire signal_2139 ;
    wire signal_2140 ;
    wire signal_2141 ;
    wire signal_2142 ;
    wire signal_2143 ;
    wire signal_2144 ;
    wire signal_2145 ;
    wire signal_2146 ;
    wire signal_2147 ;
    wire signal_2148 ;
    wire signal_2149 ;
    wire signal_2150 ;
    wire signal_2151 ;
    wire signal_2152 ;
    wire signal_2153 ;
    wire signal_2154 ;
    wire signal_2155 ;
    wire signal_2156 ;
    wire signal_2157 ;
    wire signal_2158 ;
    wire signal_2159 ;
    wire signal_2160 ;
    wire signal_2161 ;
    wire signal_2162 ;
    wire signal_2163 ;
    wire signal_2164 ;
    wire signal_2165 ;
    wire signal_2166 ;
    wire signal_2167 ;
    wire signal_2168 ;
    wire signal_2169 ;
    wire signal_2170 ;
    wire signal_2171 ;
    wire signal_2172 ;
    wire signal_2173 ;
    wire signal_2174 ;
    wire signal_2175 ;
    wire signal_2176 ;
    wire signal_2177 ;
    wire signal_2178 ;
    wire signal_2179 ;
    wire signal_2180 ;
    wire signal_2181 ;
    wire signal_2182 ;
    wire signal_2183 ;
    wire signal_2184 ;
    wire signal_2185 ;
    wire signal_2186 ;
    wire signal_2187 ;
    wire signal_2188 ;
    wire signal_2189 ;
    wire signal_2190 ;
    wire signal_2191 ;
    wire signal_2192 ;
    wire signal_2193 ;
    wire signal_2194 ;
    wire signal_2195 ;
    wire signal_2196 ;
    wire signal_2197 ;
    wire signal_2198 ;
    wire signal_2199 ;
    wire signal_2200 ;
    wire signal_2201 ;
    wire signal_2202 ;
    wire signal_2203 ;
    wire signal_2204 ;
    wire signal_2205 ;
    wire signal_2206 ;
    wire signal_2207 ;
    wire signal_2208 ;
    wire signal_2209 ;
    wire signal_2210 ;
    wire signal_2211 ;
    wire signal_2212 ;
    wire signal_2213 ;
    wire signal_2214 ;
    wire signal_2215 ;
    wire signal_2216 ;
    wire signal_2217 ;
    wire signal_2218 ;
    wire signal_2219 ;
    wire signal_2220 ;
    wire signal_2221 ;
    wire signal_2222 ;
    wire signal_2223 ;
    wire signal_2224 ;
    wire signal_2225 ;
    wire signal_2226 ;
    wire signal_2227 ;
    wire signal_2228 ;
    wire signal_2229 ;
    wire signal_2230 ;
    wire signal_2231 ;
    wire signal_2232 ;
    wire signal_2233 ;
    wire signal_2234 ;
    wire signal_2235 ;
    wire signal_2236 ;
    wire signal_2237 ;
    wire signal_2238 ;
    wire signal_2239 ;
    wire signal_2240 ;
    wire signal_2241 ;
    wire signal_2242 ;
    wire signal_2243 ;
    wire signal_2244 ;
    wire signal_2245 ;
    wire signal_2246 ;
    wire signal_2247 ;
    wire signal_2248 ;
    wire signal_2249 ;
    wire signal_2250 ;
    wire signal_2251 ;
    wire signal_2252 ;
    wire signal_2253 ;
    wire signal_2254 ;
    wire signal_2255 ;
    wire signal_2256 ;
    wire signal_2257 ;
    wire signal_2258 ;
    wire signal_2259 ;
    wire signal_2260 ;
    wire signal_2261 ;
    wire signal_2262 ;
    wire signal_2263 ;
    wire signal_2264 ;
    wire signal_2265 ;
    wire signal_2266 ;
    wire signal_2267 ;
    wire signal_2268 ;
    wire signal_2269 ;
    wire signal_2270 ;
    wire signal_2271 ;
    wire signal_2272 ;
    wire signal_2273 ;
    wire signal_2274 ;
    wire signal_2275 ;
    wire signal_2276 ;
    wire signal_2298 ;
    wire signal_2299 ;
    wire signal_2300 ;
    wire signal_2303 ;
    wire signal_2305 ;
    wire signal_2306 ;
    wire signal_2307 ;
    wire signal_2308 ;
    wire signal_2309 ;
    wire signal_2310 ;
    wire signal_2311 ;
    wire signal_2312 ;
    wire signal_2313 ;
    wire signal_2314 ;
    wire signal_2315 ;
    wire signal_2316 ;
    wire signal_2317 ;
    wire signal_2318 ;
    wire signal_2319 ;
    wire signal_2320 ;
    wire signal_2321 ;
    wire signal_2322 ;
    wire signal_2323 ;
    wire signal_2324 ;
    wire signal_2325 ;
    wire signal_2326 ;
    wire signal_2327 ;
    wire signal_2328 ;
    wire signal_2329 ;
    wire signal_2330 ;
    wire signal_2331 ;
    wire signal_2332 ;
    wire signal_2333 ;
    wire signal_2334 ;
    wire signal_2335 ;
    wire signal_2336 ;
    wire signal_2337 ;
    wire signal_2339 ;
    wire signal_2340 ;
    wire signal_2342 ;
    wire signal_2343 ;
    wire signal_2345 ;
    wire signal_2346 ;
    wire signal_2348 ;
    wire signal_2349 ;
    wire signal_2351 ;
    wire signal_2352 ;
    wire signal_2354 ;
    wire signal_2355 ;
    wire signal_2357 ;
    wire signal_2358 ;
    wire signal_2360 ;
    wire signal_2361 ;
    wire signal_2363 ;
    wire signal_2364 ;
    wire signal_2366 ;
    wire signal_2367 ;
    wire signal_2369 ;
    wire signal_2370 ;
    wire signal_2372 ;
    wire signal_2373 ;
    wire signal_2375 ;
    wire signal_2376 ;
    wire signal_2378 ;
    wire signal_2379 ;
    wire signal_2381 ;
    wire signal_2382 ;
    wire signal_2384 ;
    wire signal_2385 ;
    wire signal_2387 ;
    wire signal_2388 ;
    wire signal_2390 ;
    wire signal_2391 ;
    wire signal_2393 ;
    wire signal_2394 ;
    wire signal_2396 ;
    wire signal_2397 ;
    wire signal_2399 ;
    wire signal_2400 ;
    wire signal_2402 ;
    wire signal_2403 ;
    wire signal_2405 ;
    wire signal_2406 ;
    wire signal_2408 ;
    wire signal_2409 ;
    wire signal_2411 ;
    wire signal_2412 ;
    wire signal_2414 ;
    wire signal_2415 ;
    wire signal_2417 ;
    wire signal_2418 ;
    wire signal_2420 ;
    wire signal_2421 ;
    wire signal_2423 ;
    wire signal_2424 ;
    wire signal_2426 ;
    wire signal_2427 ;
    wire signal_2429 ;
    wire signal_2430 ;
    wire signal_2432 ;
    wire signal_2433 ;
    wire signal_2435 ;
    wire signal_2436 ;
    wire signal_2438 ;
    wire signal_2439 ;
    wire signal_2441 ;
    wire signal_2442 ;
    wire signal_2444 ;
    wire signal_2445 ;
    wire signal_2447 ;
    wire signal_2448 ;
    wire signal_2450 ;
    wire signal_2451 ;
    wire signal_2453 ;
    wire signal_2454 ;
    wire signal_2456 ;
    wire signal_2457 ;
    wire signal_2459 ;
    wire signal_2460 ;
    wire signal_2462 ;
    wire signal_2463 ;
    wire signal_2465 ;
    wire signal_2466 ;
    wire signal_2468 ;
    wire signal_2469 ;
    wire signal_2471 ;
    wire signal_2472 ;
    wire signal_2474 ;
    wire signal_2475 ;
    wire signal_2477 ;
    wire signal_2478 ;
    wire signal_2480 ;
    wire signal_2481 ;
    wire signal_2483 ;
    wire signal_2484 ;
    wire signal_2486 ;
    wire signal_2487 ;
    wire signal_2489 ;
    wire signal_2490 ;
    wire signal_2492 ;
    wire signal_2493 ;
    wire signal_2495 ;
    wire signal_2496 ;
    wire signal_2498 ;
    wire signal_2499 ;
    wire signal_2501 ;
    wire signal_2502 ;
    wire signal_2504 ;
    wire signal_2505 ;
    wire signal_2507 ;
    wire signal_2508 ;
    wire signal_2510 ;
    wire signal_2511 ;
    wire signal_2513 ;
    wire signal_2514 ;
    wire signal_2516 ;
    wire signal_2517 ;
    wire signal_2519 ;
    wire signal_2520 ;
    wire signal_2522 ;
    wire signal_2523 ;
    wire signal_2525 ;
    wire signal_2526 ;
    wire signal_2528 ;
    wire signal_2529 ;
    wire signal_2531 ;
    wire signal_2532 ;
    wire signal_2534 ;
    wire signal_2535 ;
    wire signal_2537 ;
    wire signal_2538 ;
    wire signal_2540 ;
    wire signal_2541 ;
    wire signal_2543 ;
    wire signal_2544 ;
    wire signal_2546 ;
    wire signal_2547 ;
    wire signal_2549 ;
    wire signal_2550 ;
    wire signal_2552 ;
    wire signal_2553 ;
    wire signal_2555 ;
    wire signal_2556 ;
    wire signal_2558 ;
    wire signal_2559 ;
    wire signal_2561 ;
    wire signal_2562 ;
    wire signal_2564 ;
    wire signal_2565 ;
    wire signal_2567 ;
    wire signal_2568 ;
    wire signal_2570 ;
    wire signal_2571 ;
    wire signal_2573 ;
    wire signal_2574 ;
    wire signal_2576 ;
    wire signal_2577 ;
    wire signal_2579 ;
    wire signal_2580 ;
    wire signal_2582 ;
    wire signal_2583 ;
    wire signal_2585 ;
    wire signal_2586 ;
    wire signal_2588 ;
    wire signal_2589 ;
    wire signal_2591 ;
    wire signal_2592 ;
    wire signal_2594 ;
    wire signal_2595 ;
    wire signal_2597 ;
    wire signal_2598 ;
    wire signal_2600 ;
    wire signal_2601 ;
    wire signal_2603 ;
    wire signal_2604 ;
    wire signal_2606 ;
    wire signal_2607 ;
    wire signal_2609 ;
    wire signal_2610 ;
    wire signal_2612 ;
    wire signal_2613 ;
    wire signal_2615 ;
    wire signal_2616 ;
    wire signal_2618 ;
    wire signal_2619 ;
    wire signal_2621 ;
    wire signal_2622 ;
    wire signal_2624 ;
    wire signal_2625 ;
    wire signal_2627 ;
    wire signal_2628 ;
    wire signal_2630 ;
    wire signal_2631 ;
    wire signal_2633 ;
    wire signal_2634 ;
    wire signal_2636 ;
    wire signal_2637 ;
    wire signal_2639 ;
    wire signal_2640 ;
    wire signal_2642 ;
    wire signal_2643 ;
    wire signal_2645 ;
    wire signal_2646 ;
    wire signal_2648 ;
    wire signal_2649 ;
    wire signal_2651 ;
    wire signal_2652 ;
    wire signal_2654 ;
    wire signal_2655 ;
    wire signal_2657 ;
    wire signal_2658 ;
    wire signal_2660 ;
    wire signal_2661 ;
    wire signal_2663 ;
    wire signal_2664 ;
    wire signal_2666 ;
    wire signal_2667 ;
    wire signal_2669 ;
    wire signal_2670 ;
    wire signal_2672 ;
    wire signal_2673 ;
    wire signal_2675 ;
    wire signal_2676 ;
    wire signal_2678 ;
    wire signal_2679 ;
    wire signal_2681 ;
    wire signal_2682 ;
    wire signal_2684 ;
    wire signal_2685 ;
    wire signal_2687 ;
    wire signal_2688 ;
    wire signal_2690 ;
    wire signal_2691 ;
    wire signal_2693 ;
    wire signal_2694 ;
    wire signal_2696 ;
    wire signal_2697 ;
    wire signal_2699 ;
    wire signal_2700 ;
    wire signal_2702 ;
    wire signal_2703 ;
    wire signal_2705 ;
    wire signal_2706 ;
    wire signal_2708 ;
    wire signal_2709 ;
    wire signal_2711 ;
    wire signal_2712 ;
    wire signal_2714 ;
    wire signal_2715 ;
    wire signal_2717 ;
    wire signal_2718 ;
    wire signal_2720 ;
    wire signal_2721 ;
    wire signal_2722 ;
    wire signal_2723 ;
    wire signal_2724 ;
    wire signal_2725 ;
    wire signal_2726 ;
    wire signal_2727 ;
    wire signal_2728 ;
    wire signal_2729 ;
    wire signal_2730 ;
    wire signal_2731 ;
    wire signal_2732 ;
    wire signal_2733 ;
    wire signal_2734 ;
    wire signal_2735 ;
    wire signal_2736 ;
    wire signal_2737 ;
    wire signal_2738 ;
    wire signal_2739 ;
    wire signal_2740 ;
    wire signal_2741 ;
    wire signal_2742 ;
    wire signal_2743 ;
    wire signal_2744 ;
    wire signal_2745 ;
    wire signal_2746 ;
    wire signal_2747 ;
    wire signal_2748 ;
    wire signal_2749 ;
    wire signal_2750 ;
    wire signal_2751 ;
    wire signal_2752 ;
    wire signal_2753 ;
    wire signal_2754 ;
    wire signal_2755 ;
    wire signal_2756 ;
    wire signal_2757 ;
    wire signal_2758 ;
    wire signal_2759 ;
    wire signal_2760 ;
    wire signal_2761 ;
    wire signal_2762 ;
    wire signal_2763 ;
    wire signal_2764 ;
    wire signal_2765 ;
    wire signal_2766 ;
    wire signal_2767 ;
    wire signal_2768 ;
    wire signal_2769 ;
    wire signal_2770 ;
    wire signal_2771 ;
    wire signal_2772 ;
    wire signal_2773 ;
    wire signal_2774 ;
    wire signal_2775 ;
    wire signal_2776 ;
    wire signal_2777 ;
    wire signal_2778 ;
    wire signal_2779 ;
    wire signal_2780 ;
    wire signal_2781 ;
    wire signal_2782 ;
    wire signal_2783 ;
    wire signal_2784 ;
    wire signal_2785 ;
    wire signal_2786 ;
    wire signal_2787 ;
    wire signal_2788 ;
    wire signal_2789 ;
    wire signal_2790 ;
    wire signal_2791 ;
    wire signal_2792 ;
    wire signal_2793 ;
    wire signal_2794 ;
    wire signal_2795 ;
    wire signal_2796 ;
    wire signal_2797 ;
    wire signal_2798 ;
    wire signal_2799 ;
    wire signal_2800 ;
    wire signal_2801 ;
    wire signal_2802 ;
    wire signal_2803 ;
    wire signal_2804 ;
    wire signal_2805 ;
    wire signal_2806 ;
    wire signal_2807 ;
    wire signal_2808 ;
    wire signal_2809 ;
    wire signal_2810 ;
    wire signal_2811 ;
    wire signal_2812 ;
    wire signal_2813 ;
    wire signal_2814 ;
    wire signal_2815 ;
    wire signal_2816 ;
    wire signal_2817 ;
    wire signal_2818 ;
    wire signal_2819 ;
    wire signal_2820 ;
    wire signal_2821 ;
    wire signal_2822 ;
    wire signal_2823 ;
    wire signal_2824 ;
    wire signal_2825 ;
    wire signal_2826 ;
    wire signal_2827 ;
    wire signal_2828 ;
    wire signal_2829 ;
    wire signal_2830 ;
    wire signal_2831 ;
    wire signal_2832 ;
    wire signal_2833 ;
    wire signal_2834 ;
    wire signal_2835 ;
    wire signal_2836 ;
    wire signal_2837 ;
    wire signal_2838 ;
    wire signal_2839 ;
    wire signal_2840 ;
    wire signal_2841 ;
    wire signal_2842 ;
    wire signal_2843 ;
    wire signal_2844 ;
    wire signal_2845 ;
    wire signal_2846 ;
    wire signal_2847 ;
    wire signal_2848 ;
    wire signal_2849 ;
    wire signal_2851 ;
    wire signal_2853 ;
    wire signal_2855 ;
    wire signal_2857 ;
    wire signal_2859 ;
    wire signal_2861 ;
    wire signal_2863 ;
    wire signal_2865 ;
    wire signal_2867 ;
    wire signal_2869 ;
    wire signal_2871 ;
    wire signal_2873 ;
    wire signal_2875 ;
    wire signal_2877 ;
    wire signal_2879 ;
    wire signal_2881 ;
    wire signal_2883 ;
    wire signal_2885 ;
    wire signal_2887 ;
    wire signal_2889 ;
    wire signal_2891 ;
    wire signal_2893 ;
    wire signal_2895 ;
    wire signal_2897 ;
    wire signal_2899 ;
    wire signal_2901 ;
    wire signal_2903 ;
    wire signal_2905 ;
    wire signal_2907 ;
    wire signal_2909 ;
    wire signal_2911 ;
    wire signal_2913 ;
    wire signal_2915 ;
    wire signal_2917 ;
    wire signal_2919 ;
    wire signal_2921 ;
    wire signal_2923 ;
    wire signal_2925 ;
    wire signal_2927 ;
    wire signal_2929 ;
    wire signal_2931 ;
    wire signal_2933 ;
    wire signal_2935 ;
    wire signal_2937 ;
    wire signal_2939 ;
    wire signal_2941 ;
    wire signal_2943 ;
    wire signal_2945 ;
    wire signal_2947 ;
    wire signal_2949 ;
    wire signal_2951 ;
    wire signal_2953 ;
    wire signal_2955 ;
    wire signal_2957 ;
    wire signal_2959 ;
    wire signal_2961 ;
    wire signal_2963 ;
    wire signal_2965 ;
    wire signal_2967 ;
    wire signal_2969 ;
    wire signal_2971 ;
    wire signal_2973 ;
    wire signal_2975 ;
    wire signal_2977 ;
    wire signal_2979 ;
    wire signal_2981 ;
    wire signal_2983 ;
    wire signal_2985 ;
    wire signal_2987 ;
    wire signal_2989 ;
    wire signal_2991 ;
    wire signal_2993 ;
    wire signal_2995 ;
    wire signal_2997 ;
    wire signal_2999 ;
    wire signal_3001 ;
    wire signal_3003 ;
    wire signal_3005 ;
    wire signal_3007 ;
    wire signal_3009 ;
    wire signal_3011 ;
    wire signal_3013 ;
    wire signal_3015 ;
    wire signal_3017 ;
    wire signal_3019 ;
    wire signal_3021 ;
    wire signal_3023 ;
    wire signal_3025 ;
    wire signal_3027 ;
    wire signal_3029 ;
    wire signal_3031 ;
    wire signal_3033 ;
    wire signal_3035 ;
    wire signal_3037 ;
    wire signal_3039 ;
    wire signal_3041 ;
    wire signal_3042 ;
    wire signal_3043 ;
    wire signal_3044 ;
    wire signal_3045 ;
    wire signal_3046 ;
    wire signal_3047 ;
    wire signal_3048 ;
    wire signal_3049 ;
    wire signal_3050 ;
    wire signal_3051 ;
    wire signal_3052 ;
    wire signal_3053 ;
    wire signal_3054 ;
    wire signal_3055 ;
    wire signal_3056 ;
    wire signal_3057 ;
    wire signal_3058 ;
    wire signal_3059 ;
    wire signal_3060 ;
    wire signal_3061 ;
    wire signal_3062 ;
    wire signal_3063 ;
    wire signal_3064 ;
    wire signal_3065 ;
    wire signal_3066 ;
    wire signal_3067 ;
    wire signal_3068 ;
    wire signal_3069 ;
    wire signal_3070 ;
    wire signal_3071 ;
    wire signal_3072 ;
    wire signal_3073 ;
    wire signal_3074 ;
    wire signal_3075 ;
    wire signal_3076 ;
    wire signal_3077 ;
    wire signal_3078 ;
    wire signal_3079 ;
    wire signal_3080 ;
    wire signal_3081 ;
    wire signal_3082 ;
    wire signal_3083 ;
    wire signal_3084 ;
    wire signal_3085 ;
    wire signal_3086 ;
    wire signal_3087 ;
    wire signal_3088 ;
    wire signal_3089 ;
    wire signal_3090 ;
    wire signal_3091 ;
    wire signal_3092 ;
    wire signal_3093 ;
    wire signal_3094 ;
    wire signal_3095 ;
    wire signal_3096 ;
    wire signal_3097 ;
    wire signal_3098 ;
    wire signal_3099 ;
    wire signal_3100 ;
    wire signal_3101 ;
    wire signal_3102 ;
    wire signal_3103 ;
    wire signal_3104 ;
    wire signal_3105 ;
    wire signal_3106 ;
    wire signal_3107 ;
    wire signal_3108 ;
    wire signal_3109 ;
    wire signal_3110 ;
    wire signal_3111 ;
    wire signal_3112 ;
    wire signal_3113 ;
    wire signal_3114 ;
    wire signal_3115 ;
    wire signal_3116 ;
    wire signal_3117 ;
    wire signal_3118 ;
    wire signal_3119 ;
    wire signal_3120 ;
    wire signal_3121 ;
    wire signal_3122 ;
    wire signal_3123 ;
    wire signal_3124 ;
    wire signal_3125 ;
    wire signal_3126 ;
    wire signal_3127 ;
    wire signal_3128 ;
    wire signal_3129 ;
    wire signal_3130 ;
    wire signal_3131 ;
    wire signal_3132 ;
    wire signal_3133 ;
    wire signal_3134 ;
    wire signal_3135 ;
    wire signal_3136 ;
    wire signal_3137 ;
    wire signal_3138 ;
    wire signal_3139 ;
    wire signal_3140 ;
    wire signal_3141 ;
    wire signal_3142 ;
    wire signal_3143 ;
    wire signal_3144 ;
    wire signal_3145 ;
    wire signal_3146 ;
    wire signal_3147 ;
    wire signal_3148 ;
    wire signal_3149 ;
    wire signal_3150 ;
    wire signal_3151 ;
    wire signal_3152 ;
    wire signal_3153 ;
    wire signal_3154 ;
    wire signal_3155 ;
    wire signal_3156 ;
    wire signal_3157 ;
    wire signal_3158 ;
    wire signal_3159 ;
    wire signal_3160 ;
    wire signal_3161 ;
    wire signal_3162 ;
    wire signal_3163 ;
    wire signal_3164 ;
    wire signal_3165 ;
    wire signal_3166 ;
    wire signal_3167 ;
    wire signal_3168 ;
    wire signal_3169 ;
    wire signal_3170 ;
    wire signal_3171 ;
    wire signal_3172 ;
    wire signal_3173 ;
    wire signal_3174 ;
    wire signal_3175 ;
    wire signal_3176 ;
    wire signal_3177 ;
    wire signal_3178 ;
    wire signal_3179 ;
    wire signal_3180 ;
    wire signal_3181 ;
    wire signal_3182 ;
    wire signal_3183 ;
    wire signal_3184 ;
    wire signal_3185 ;
    wire signal_3186 ;
    wire signal_3187 ;
    wire signal_3188 ;
    wire signal_3189 ;
    wire signal_3190 ;
    wire signal_3191 ;
    wire signal_3192 ;
    wire signal_3193 ;
    wire signal_3194 ;
    wire signal_3195 ;
    wire signal_3196 ;
    wire signal_3197 ;
    wire signal_3198 ;
    wire signal_3199 ;
    wire signal_3200 ;
    wire signal_3201 ;
    wire signal_3202 ;
    wire signal_3203 ;
    wire signal_3204 ;
    wire signal_3205 ;
    wire signal_3206 ;
    wire signal_3207 ;
    wire signal_3208 ;
    wire signal_3209 ;
    wire signal_3210 ;
    wire signal_3211 ;
    wire signal_3212 ;
    wire signal_3213 ;
    wire signal_3214 ;
    wire signal_3215 ;
    wire signal_3216 ;
    wire signal_3217 ;
    wire signal_3218 ;
    wire signal_3219 ;
    wire signal_3220 ;
    wire signal_3221 ;
    wire signal_3222 ;
    wire signal_3223 ;
    wire signal_3224 ;
    wire signal_3225 ;
    wire signal_3226 ;
    wire signal_3227 ;
    wire signal_3228 ;
    wire signal_3229 ;
    wire signal_3230 ;
    wire signal_3231 ;
    wire signal_3232 ;
    wire signal_3233 ;
    wire signal_3234 ;
    wire signal_3235 ;
    wire signal_3236 ;
    wire signal_3237 ;
    wire signal_3238 ;
    wire signal_3239 ;
    wire signal_3240 ;
    wire signal_3241 ;
    wire signal_3242 ;
    wire signal_3243 ;
    wire signal_3244 ;
    wire signal_3245 ;
    wire signal_3246 ;
    wire signal_3247 ;
    wire signal_3248 ;
    wire signal_3249 ;
    wire signal_3250 ;
    wire signal_3251 ;
    wire signal_3252 ;
    wire signal_3253 ;
    wire signal_3254 ;
    wire signal_3255 ;
    wire signal_3256 ;
    wire signal_3257 ;
    wire signal_3258 ;
    wire signal_3259 ;
    wire signal_3260 ;
    wire signal_3261 ;
    wire signal_3263 ;
    wire signal_3265 ;
    wire signal_3267 ;
    wire signal_3269 ;
    wire signal_3271 ;
    wire signal_3273 ;
    wire signal_3275 ;
    wire signal_3277 ;
    wire signal_3279 ;
    wire signal_3281 ;
    wire signal_3283 ;
    wire signal_3285 ;
    wire signal_3287 ;
    wire signal_3289 ;
    wire signal_3291 ;
    wire signal_3293 ;
    wire signal_3295 ;
    wire signal_3297 ;
    wire signal_3299 ;
    wire signal_3301 ;
    wire signal_3303 ;
    wire signal_3305 ;
    wire signal_3307 ;
    wire signal_3309 ;
    wire signal_3311 ;
    wire signal_3313 ;
    wire signal_3315 ;
    wire signal_3317 ;
    wire signal_3319 ;
    wire signal_3321 ;
    wire signal_3322 ;
    wire signal_3323 ;
    wire signal_3325 ;
    wire signal_3327 ;
    wire signal_3329 ;
    wire signal_3331 ;
    wire signal_3333 ;
    wire signal_3335 ;
    wire signal_3337 ;
    wire signal_3339 ;
    wire signal_3341 ;
    wire signal_3343 ;
    wire signal_3345 ;
    wire signal_3347 ;
    wire signal_3349 ;
    wire signal_3351 ;
    wire signal_3353 ;
    wire signal_3355 ;
    wire signal_3357 ;
    wire signal_3359 ;
    wire signal_3361 ;
    wire signal_3363 ;
    wire signal_3365 ;
    wire signal_3367 ;
    wire signal_3369 ;
    wire signal_3371 ;
    wire signal_3372 ;
    wire signal_3373 ;
    wire signal_3374 ;
    wire signal_3375 ;
    wire signal_3376 ;
    wire signal_3377 ;
    wire signal_3378 ;
    wire signal_3379 ;
    wire signal_3380 ;
    wire signal_3381 ;
    wire signal_3382 ;
    wire signal_3383 ;
    wire signal_3384 ;
    wire signal_3385 ;
    wire signal_3386 ;
    wire signal_3387 ;
    wire signal_3388 ;
    wire signal_3389 ;
    wire signal_3390 ;
    wire signal_3391 ;
    wire signal_3392 ;
    wire signal_3393 ;
    wire signal_3394 ;
    wire signal_3395 ;
    wire signal_3396 ;
    wire signal_3397 ;
    wire signal_3398 ;
    wire signal_3399 ;
    wire signal_3400 ;
    wire signal_3401 ;
    wire signal_3402 ;
    wire signal_3403 ;
    wire signal_3404 ;
    wire signal_3405 ;
    wire signal_3406 ;
    wire signal_3407 ;
    wire signal_3408 ;
    wire signal_3409 ;
    wire signal_3410 ;
    wire signal_3411 ;
    wire signal_3412 ;
    wire signal_3413 ;
    wire signal_3414 ;
    wire signal_3415 ;
    wire signal_3416 ;
    wire signal_3417 ;
    wire signal_3418 ;
    wire signal_3419 ;
    wire signal_3420 ;
    wire signal_3421 ;
    wire signal_3422 ;
    wire signal_3423 ;
    wire signal_3424 ;
    wire signal_3425 ;
    wire signal_3426 ;
    wire signal_3427 ;
    wire signal_3428 ;
    wire signal_3429 ;
    wire signal_3430 ;
    wire signal_3431 ;
    wire signal_3432 ;
    wire signal_3433 ;
    wire signal_3434 ;
    wire signal_3435 ;
    wire signal_3437 ;
    wire signal_3439 ;
    wire signal_3441 ;
    wire signal_3443 ;
    wire signal_3445 ;
    wire signal_3447 ;
    wire signal_3449 ;
    wire signal_3451 ;
    wire signal_3453 ;
    wire signal_3455 ;
    wire signal_3457 ;
    wire signal_3459 ;
    wire signal_3461 ;
    wire signal_3463 ;
    wire signal_3465 ;
    wire signal_3467 ;
    wire signal_3469 ;
    wire signal_3471 ;
    wire signal_3473 ;
    wire signal_3475 ;
    wire signal_3477 ;
    wire signal_3479 ;
    wire signal_3481 ;
    wire signal_3483 ;
    wire signal_3485 ;
    wire signal_3487 ;
    wire signal_3489 ;
    wire signal_3491 ;
    wire signal_3493 ;
    wire signal_3495 ;
    wire signal_3497 ;
    wire signal_3499 ;
    wire signal_3501 ;
    wire signal_3503 ;
    wire signal_3504 ;
    wire signal_3505 ;
    wire signal_3506 ;
    wire signal_3507 ;
    wire signal_3508 ;
    wire signal_3509 ;
    wire signal_3510 ;
    wire signal_3511 ;
    wire signal_3512 ;
    wire signal_3513 ;
    wire signal_3514 ;
    wire signal_3515 ;
    wire signal_3516 ;
    wire signal_3517 ;
    wire signal_3518 ;
    wire signal_3519 ;
    wire signal_3520 ;
    wire signal_3521 ;
    wire signal_3522 ;
    wire signal_3523 ;
    wire signal_3524 ;
    wire signal_3525 ;
    wire signal_3526 ;
    wire signal_3527 ;
    wire signal_3528 ;
    wire signal_3529 ;
    wire signal_3530 ;
    wire signal_3531 ;
    wire signal_3532 ;
    wire signal_3533 ;
    wire signal_3534 ;
    wire signal_3535 ;
    wire signal_3536 ;
    wire signal_3537 ;
    wire signal_3538 ;
    wire signal_3539 ;
    wire signal_3540 ;
    wire signal_3541 ;
    wire signal_3542 ;
    wire signal_3543 ;
    wire signal_3544 ;
    wire signal_3545 ;
    wire signal_3546 ;
    wire signal_3547 ;
    wire signal_3548 ;
    wire signal_3549 ;
    wire signal_3550 ;
    wire signal_3551 ;
    wire signal_3552 ;
    wire signal_3553 ;
    wire signal_3554 ;
    wire signal_3555 ;
    wire signal_3556 ;
    wire signal_3557 ;
    wire signal_3558 ;
    wire signal_3559 ;
    wire signal_3560 ;
    wire signal_3561 ;
    wire signal_3562 ;
    wire signal_3563 ;
    wire signal_3564 ;
    wire signal_3565 ;
    wire signal_3566 ;
    wire signal_3567 ;
    wire signal_3569 ;
    wire signal_3571 ;
    wire signal_3573 ;
    wire signal_3575 ;
    wire signal_3577 ;
    wire signal_3579 ;
    wire signal_3581 ;
    wire signal_3583 ;
    wire signal_3585 ;
    wire signal_3587 ;
    wire signal_3589 ;
    wire signal_3591 ;
    wire signal_3593 ;
    wire signal_3595 ;
    wire signal_3597 ;
    wire signal_3599 ;
    wire signal_3601 ;
    wire signal_3603 ;
    wire signal_3605 ;
    wire signal_3607 ;
    wire signal_3609 ;
    wire signal_3611 ;
    wire signal_3613 ;
    wire signal_3615 ;
    wire signal_3617 ;
    wire signal_3619 ;
    wire signal_3621 ;
    wire signal_3623 ;
    wire signal_3625 ;
    wire signal_3627 ;
    wire signal_3629 ;
    wire signal_3631 ;
    wire signal_3632 ;
    wire signal_3633 ;
    wire signal_3634 ;
    wire signal_3635 ;
    wire signal_3636 ;
    wire signal_3637 ;
    wire signal_3638 ;
    wire signal_3639 ;
    wire signal_3640 ;
    wire signal_3641 ;
    wire signal_3642 ;
    wire signal_3643 ;
    wire signal_3644 ;
    wire signal_3645 ;
    wire signal_3646 ;
    wire signal_3647 ;
    wire signal_3648 ;
    wire signal_3649 ;
    wire signal_3650 ;
    wire signal_3651 ;
    wire signal_3652 ;
    wire signal_3653 ;
    wire signal_3654 ;
    wire signal_3655 ;
    wire signal_3656 ;
    wire signal_3657 ;
    wire signal_3658 ;
    wire signal_3659 ;
    wire signal_3660 ;
    wire signal_3661 ;
    wire signal_3662 ;
    wire signal_3663 ;
    wire signal_3664 ;
    wire signal_3665 ;
    wire signal_3666 ;
    wire signal_3667 ;
    wire signal_3668 ;
    wire signal_3669 ;
    wire signal_3670 ;
    wire signal_3671 ;
    wire signal_3673 ;
    wire signal_3675 ;
    wire signal_3677 ;
    wire signal_3679 ;
    wire signal_3681 ;
    wire signal_3683 ;
    wire signal_3685 ;
    wire signal_3687 ;
    wire signal_3689 ;
    wire signal_3691 ;
    wire signal_3693 ;
    wire signal_3695 ;
    wire signal_3697 ;
    wire signal_3699 ;
    wire signal_3701 ;
    wire signal_3703 ;
    wire signal_3705 ;
    wire signal_3707 ;
    wire signal_3709 ;
    wire signal_3711 ;
    wire signal_3713 ;
    wire signal_3715 ;
    wire signal_3717 ;
    wire signal_3719 ;
    wire signal_3721 ;
    wire signal_3723 ;
    wire signal_3725 ;
    wire signal_3727 ;
    wire signal_3729 ;
    wire signal_3731 ;
    wire signal_3733 ;
    wire signal_3735 ;
    wire signal_3736 ;
    wire signal_3737 ;
    wire signal_3738 ;
    wire signal_3739 ;
    wire signal_3740 ;
    wire signal_3741 ;
    wire signal_3742 ;
    wire signal_3743 ;
    wire signal_3745 ;
    wire signal_3747 ;
    wire signal_3749 ;
    wire signal_3751 ;
    wire signal_3753 ;
    wire signal_3755 ;
    wire signal_3757 ;
    wire signal_3759 ;
    wire signal_11952 ;
    wire signal_11953 ;
    wire signal_11954 ;
    wire signal_11955 ;
    wire signal_11956 ;
    wire signal_11957 ;
    wire signal_11958 ;
    wire signal_11959 ;
    wire signal_11960 ;
    wire signal_11961 ;
    wire signal_11962 ;
    wire signal_11963 ;
    wire signal_11964 ;
    wire signal_11965 ;
    wire signal_11966 ;
    wire signal_11967 ;
    wire signal_11968 ;
    wire signal_11969 ;
    wire signal_11970 ;
    wire signal_11971 ;
    wire signal_11972 ;
    wire signal_11973 ;
    wire signal_11974 ;
    wire signal_11975 ;
    wire signal_11976 ;
    wire signal_11977 ;
    wire signal_11978 ;
    wire signal_11979 ;
    wire signal_11980 ;
    wire signal_11981 ;
    wire signal_11982 ;
    wire signal_11983 ;
    wire signal_11984 ;
    wire signal_11985 ;
    wire signal_11986 ;
    wire signal_11987 ;
    wire signal_11988 ;
    wire signal_11989 ;
    wire signal_11990 ;
    wire signal_11991 ;
    wire signal_11992 ;
    wire signal_11993 ;
    wire signal_11994 ;
    wire signal_11995 ;
    wire signal_11996 ;
    wire signal_11997 ;
    wire signal_11998 ;
    wire signal_11999 ;
    wire signal_12000 ;
    wire signal_12001 ;
    wire signal_12002 ;
    wire signal_12003 ;
    wire signal_12004 ;
    wire signal_12005 ;
    wire signal_12006 ;
    wire signal_12007 ;
    wire signal_12008 ;
    wire signal_12009 ;
    wire signal_12010 ;
    wire signal_12011 ;
    wire signal_12012 ;
    wire signal_12013 ;
    wire signal_12014 ;
    wire signal_12015 ;
    wire signal_12016 ;
    wire signal_12017 ;
    wire signal_12018 ;
    wire signal_12019 ;
    wire signal_12020 ;
    wire signal_12021 ;
    wire signal_12022 ;
    wire signal_12023 ;
    wire signal_12024 ;
    wire signal_12025 ;
    wire signal_12026 ;
    wire signal_12027 ;
    wire signal_12028 ;
    wire signal_12029 ;
    wire signal_12030 ;
    wire signal_12031 ;
    wire signal_12032 ;
    wire signal_12033 ;
    wire signal_12034 ;
    wire signal_12035 ;
    wire signal_12036 ;
    wire signal_12037 ;
    wire signal_12038 ;
    wire signal_12039 ;
    wire signal_12040 ;
    wire signal_12041 ;
    wire signal_12042 ;
    wire signal_12043 ;
    wire signal_12044 ;
    wire signal_12045 ;
    wire signal_12046 ;
    wire signal_12047 ;
    wire signal_12048 ;
    wire signal_12049 ;
    wire signal_12050 ;
    wire signal_12051 ;
    wire signal_12052 ;
    wire signal_12053 ;
    wire signal_12054 ;
    wire signal_12055 ;
    wire signal_12056 ;
    wire signal_12057 ;
    wire signal_12058 ;
    wire signal_12059 ;
    wire signal_12060 ;
    wire signal_12061 ;
    wire signal_12062 ;
    wire signal_12063 ;
    wire signal_12064 ;
    wire signal_12065 ;
    wire signal_12066 ;
    wire signal_12067 ;
    wire signal_12068 ;
    wire signal_12069 ;
    wire signal_12070 ;
    wire signal_12071 ;
    wire signal_12072 ;
    wire signal_12073 ;
    wire signal_12074 ;
    wire signal_12075 ;
    wire signal_12076 ;
    wire signal_12077 ;
    wire signal_12078 ;
    wire signal_12079 ;
    wire signal_12080 ;
    wire signal_12081 ;
    wire signal_12082 ;
    wire signal_12083 ;
    wire signal_12084 ;
    wire signal_12085 ;
    wire signal_12086 ;
    wire signal_12087 ;
    wire signal_12088 ;
    wire signal_12089 ;
    wire signal_12090 ;
    wire signal_12091 ;
    wire signal_12092 ;
    wire signal_12093 ;
    wire signal_12094 ;
    wire signal_12095 ;
    wire signal_12096 ;
    wire signal_12097 ;
    wire signal_12098 ;
    wire signal_12099 ;
    wire signal_12100 ;
    wire signal_12101 ;
    wire signal_12102 ;
    wire signal_12103 ;
    wire signal_12104 ;
    wire signal_12105 ;
    wire signal_12106 ;
    wire signal_12107 ;
    wire signal_12108 ;
    wire signal_12109 ;
    wire signal_12110 ;
    wire signal_12111 ;
    wire signal_12112 ;
    wire signal_12113 ;
    wire signal_12114 ;
    wire signal_12115 ;
    wire signal_12116 ;
    wire signal_12117 ;
    wire signal_12118 ;
    wire signal_12119 ;
    wire signal_12120 ;
    wire signal_12121 ;
    wire signal_12122 ;
    wire signal_12123 ;
    wire signal_12124 ;
    wire signal_12125 ;
    wire signal_12126 ;
    wire signal_12127 ;
    wire signal_12128 ;
    wire signal_12129 ;
    wire signal_12130 ;
    wire signal_12131 ;
    wire signal_12132 ;
    wire signal_12133 ;
    wire signal_12134 ;
    wire signal_12135 ;
    wire signal_12136 ;
    wire signal_12137 ;
    wire signal_12138 ;
    wire signal_12139 ;
    wire signal_12140 ;
    wire signal_12141 ;
    wire signal_12142 ;
    wire signal_12143 ;
    wire signal_12144 ;
    wire signal_12145 ;
    wire signal_12146 ;
    wire signal_12147 ;
    wire signal_12148 ;
    wire signal_12149 ;
    wire signal_12150 ;
    wire signal_12151 ;
    wire signal_12152 ;
    wire signal_12153 ;
    wire signal_12154 ;
    wire signal_12155 ;
    wire signal_12156 ;
    wire signal_12157 ;
    wire signal_12158 ;
    wire signal_12159 ;
    wire signal_12160 ;
    wire signal_12161 ;
    wire signal_12162 ;
    wire signal_12163 ;
    wire signal_12164 ;
    wire signal_12165 ;
    wire signal_12166 ;
    wire signal_12167 ;
    wire signal_12168 ;
    wire signal_12169 ;
    wire signal_12170 ;
    wire signal_12171 ;
    wire signal_12172 ;
    wire signal_12173 ;
    wire signal_12174 ;
    wire signal_12175 ;
    wire signal_12176 ;
    wire signal_12177 ;
    wire signal_12178 ;
    wire signal_12179 ;
    wire signal_12180 ;
    wire signal_12181 ;
    wire signal_12182 ;
    wire signal_12183 ;
    wire signal_12184 ;
    wire signal_12185 ;
    wire signal_12186 ;
    wire signal_12187 ;
    wire signal_12188 ;
    wire signal_12189 ;
    wire signal_12190 ;
    wire signal_12191 ;
    wire signal_12192 ;
    wire signal_12193 ;
    wire signal_12194 ;
    wire signal_12195 ;
    wire signal_12196 ;
    wire signal_12197 ;
    wire signal_12198 ;
    wire signal_12199 ;
    wire signal_12200 ;
    wire signal_12201 ;
    wire signal_12202 ;
    wire signal_12203 ;
    wire signal_12204 ;
    wire signal_12205 ;
    wire signal_12206 ;
    wire signal_12207 ;
    wire signal_12208 ;
    wire signal_12209 ;
    wire signal_12210 ;
    wire signal_12211 ;
    wire signal_12212 ;
    wire signal_12213 ;
    wire signal_12214 ;
    wire signal_12215 ;
    wire signal_12216 ;
    wire signal_12217 ;
    wire signal_12218 ;
    wire signal_12219 ;
    wire signal_12220 ;
    wire signal_12221 ;
    wire signal_12222 ;
    wire signal_12223 ;
    wire signal_12224 ;
    wire signal_12225 ;
    wire signal_12226 ;
    wire signal_12227 ;
    wire signal_12228 ;
    wire signal_12229 ;
    wire signal_12230 ;
    wire signal_12231 ;
    wire signal_12232 ;
    wire signal_12233 ;
    wire signal_12234 ;
    wire signal_12235 ;
    wire signal_12236 ;
    wire signal_12237 ;
    wire signal_12238 ;
    wire signal_12239 ;
    wire signal_12240 ;
    wire signal_12241 ;
    wire signal_12242 ;
    wire signal_12243 ;
    wire signal_12244 ;
    wire signal_12245 ;
    wire signal_12246 ;
    wire signal_12247 ;
    wire signal_12248 ;
    wire signal_12249 ;
    wire signal_12250 ;
    wire signal_12251 ;
    wire signal_12252 ;
    wire signal_12253 ;
    wire signal_12254 ;
    wire signal_12255 ;
    wire signal_12256 ;
    wire signal_12257 ;
    wire signal_12258 ;
    wire signal_12259 ;
    wire signal_12260 ;
    wire signal_12261 ;
    wire signal_12262 ;
    wire signal_12263 ;
    wire signal_12264 ;
    wire signal_12265 ;
    wire signal_12266 ;
    wire signal_12267 ;
    wire signal_12268 ;
    wire signal_12269 ;
    wire signal_12270 ;
    wire signal_12271 ;
    wire signal_12272 ;
    wire signal_12273 ;
    wire signal_12274 ;
    wire signal_12275 ;
    wire signal_12276 ;
    wire signal_12277 ;
    wire signal_12278 ;
    wire signal_12279 ;
    wire signal_12280 ;
    wire signal_12281 ;
    wire signal_12282 ;
    wire signal_12283 ;
    wire signal_12284 ;
    wire signal_12285 ;
    wire signal_12286 ;
    wire signal_12287 ;
    wire signal_12288 ;
    wire signal_12289 ;
    wire signal_12290 ;
    wire signal_12291 ;
    wire signal_12292 ;
    wire signal_12293 ;
    wire signal_12294 ;
    wire signal_12295 ;
    wire signal_12296 ;
    wire signal_12297 ;
    wire signal_12298 ;
    wire signal_12299 ;
    wire signal_12300 ;
    wire signal_12301 ;
    wire signal_12302 ;
    wire signal_12303 ;
    wire signal_12304 ;
    wire signal_12305 ;
    wire signal_12306 ;
    wire signal_12307 ;
    wire signal_12308 ;
    wire signal_12309 ;
    wire signal_12310 ;
    wire signal_12311 ;
    wire signal_12312 ;
    wire signal_12313 ;
    wire signal_12314 ;
    wire signal_12315 ;
    wire signal_12316 ;
    wire signal_12317 ;
    wire signal_12318 ;
    wire signal_12319 ;
    wire signal_12320 ;
    wire signal_12321 ;
    wire signal_12322 ;
    wire signal_12323 ;
    wire signal_12324 ;
    wire signal_12325 ;
    wire signal_12326 ;
    wire signal_12327 ;
    wire signal_12328 ;
    wire signal_12329 ;
    wire signal_12330 ;
    wire signal_12331 ;
    wire signal_12332 ;
    wire signal_12333 ;
    wire signal_12334 ;
    wire signal_12335 ;
    wire signal_12336 ;
    wire signal_12337 ;
    wire signal_12338 ;
    wire signal_12339 ;
    wire signal_12340 ;
    wire signal_12341 ;
    wire signal_12342 ;
    wire signal_12343 ;
    wire signal_12344 ;
    wire signal_12345 ;
    wire signal_12346 ;
    wire signal_12347 ;
    wire signal_12348 ;
    wire signal_12349 ;
    wire signal_12350 ;
    wire signal_12351 ;
    wire signal_12352 ;
    wire signal_12353 ;
    wire signal_12354 ;
    wire signal_12355 ;
    wire signal_12356 ;
    wire signal_12357 ;
    wire signal_12358 ;
    wire signal_12359 ;
    wire signal_12360 ;
    wire signal_12361 ;
    wire signal_12362 ;
    wire signal_12363 ;
    wire signal_12364 ;
    wire signal_12365 ;
    wire signal_12366 ;
    wire signal_12367 ;
    wire signal_12368 ;
    wire signal_12369 ;
    wire signal_12370 ;
    wire signal_12371 ;
    wire signal_12372 ;
    wire signal_12373 ;
    wire signal_12374 ;
    wire signal_12375 ;
    wire signal_12376 ;
    wire signal_12377 ;
    wire signal_12378 ;
    wire signal_12379 ;
    wire signal_12380 ;
    wire signal_12381 ;
    wire signal_12382 ;
    wire signal_12383 ;
    wire signal_12384 ;
    wire signal_12385 ;
    wire signal_12386 ;
    wire signal_12387 ;
    wire signal_12388 ;
    wire signal_12389 ;
    wire signal_12390 ;
    wire signal_12391 ;
    wire signal_12392 ;
    wire signal_12393 ;
    wire signal_12394 ;
    wire signal_12395 ;
    wire signal_12396 ;
    wire signal_12397 ;
    wire signal_12398 ;
    wire signal_12399 ;
    wire signal_12400 ;
    wire signal_12401 ;
    wire signal_12402 ;
    wire signal_12403 ;
    wire signal_12404 ;
    wire signal_12405 ;
    wire signal_12406 ;
    wire signal_12407 ;
    wire signal_12408 ;
    wire signal_12409 ;
    wire signal_12410 ;
    wire signal_12411 ;
    wire signal_12412 ;
    wire signal_12413 ;
    wire signal_12414 ;
    wire signal_12415 ;
    wire signal_12416 ;
    wire signal_12417 ;
    wire signal_12418 ;
    wire signal_12419 ;
    wire signal_12420 ;
    wire signal_12421 ;
    wire signal_12422 ;
    wire signal_12423 ;
    wire signal_12424 ;
    wire signal_12425 ;
    wire signal_12426 ;
    wire signal_12427 ;
    wire signal_12428 ;
    wire signal_12429 ;
    wire signal_12430 ;
    wire signal_12431 ;
    wire signal_12432 ;
    wire signal_12433 ;
    wire signal_12434 ;
    wire signal_12435 ;
    wire signal_12436 ;
    wire signal_12437 ;
    wire signal_12438 ;
    wire signal_12439 ;
    wire signal_12440 ;
    wire signal_12441 ;
    wire signal_12442 ;
    wire signal_12443 ;
    wire signal_12444 ;
    wire signal_12445 ;
    wire signal_12446 ;
    wire signal_12447 ;
    wire signal_12448 ;
    wire signal_12449 ;
    wire signal_12450 ;
    wire signal_12451 ;
    wire signal_12452 ;
    wire signal_12453 ;
    wire signal_12454 ;
    wire signal_12455 ;
    wire signal_12456 ;
    wire signal_12457 ;
    wire signal_12458 ;
    wire signal_12459 ;
    wire signal_12460 ;
    wire signal_12461 ;
    wire signal_12462 ;
    wire signal_12463 ;
    wire signal_12464 ;
    wire signal_12465 ;
    wire signal_12466 ;
    wire signal_12467 ;
    wire signal_12468 ;
    wire signal_12469 ;
    wire signal_12470 ;
    wire signal_12471 ;
    wire signal_12472 ;
    wire signal_12473 ;
    wire signal_12474 ;
    wire signal_12475 ;
    wire signal_12476 ;
    wire signal_12477 ;
    wire signal_12478 ;
    wire signal_12479 ;
    wire signal_12480 ;
    wire signal_12481 ;
    wire signal_12482 ;
    wire signal_12483 ;
    wire signal_12484 ;
    wire signal_12485 ;
    wire signal_12486 ;
    wire signal_12487 ;
    wire signal_12488 ;
    wire signal_12489 ;
    wire signal_12490 ;
    wire signal_12491 ;
    wire signal_12492 ;
    wire signal_12493 ;
    wire signal_12494 ;
    wire signal_12495 ;
    wire signal_12496 ;
    wire signal_12497 ;
    wire signal_12498 ;
    wire signal_12499 ;
    wire signal_12500 ;
    wire signal_12501 ;
    wire signal_12502 ;
    wire signal_12503 ;
    wire signal_12504 ;
    wire signal_12505 ;
    wire signal_12506 ;
    wire signal_12507 ;
    wire signal_12508 ;
    wire signal_12509 ;
    wire signal_12510 ;
    wire signal_12511 ;
    wire signal_12512 ;
    wire signal_12513 ;
    wire signal_12514 ;
    wire signal_12515 ;
    wire signal_12516 ;
    wire signal_12517 ;
    wire signal_12518 ;
    wire signal_12519 ;
    wire signal_12520 ;
    wire signal_12521 ;
    wire signal_12522 ;
    wire signal_12523 ;
    wire signal_12524 ;
    wire signal_12525 ;
    wire signal_12526 ;
    wire signal_12527 ;
    wire signal_12528 ;
    wire signal_12529 ;
    wire signal_12530 ;
    wire signal_12531 ;
    wire signal_12532 ;
    wire signal_12533 ;
    wire signal_12534 ;
    wire signal_12535 ;
    wire signal_12536 ;
    wire signal_12537 ;
    wire signal_12538 ;
    wire signal_12539 ;
    wire signal_12540 ;
    wire signal_12541 ;
    wire signal_12542 ;
    wire signal_12543 ;
    wire signal_12544 ;
    wire signal_12545 ;
    wire signal_12546 ;
    wire signal_12547 ;
    wire signal_12548 ;
    wire signal_12549 ;
    wire signal_12550 ;
    wire signal_12551 ;
    wire signal_12552 ;
    wire signal_12553 ;
    wire signal_12554 ;
    wire signal_12555 ;
    wire signal_12556 ;
    wire signal_12557 ;
    wire signal_12558 ;
    wire signal_12559 ;
    wire signal_12560 ;
    wire signal_12561 ;
    wire signal_12562 ;
    wire signal_12563 ;
    wire signal_12564 ;
    wire signal_12565 ;
    wire signal_12566 ;
    wire signal_12567 ;
    wire signal_12568 ;
    wire signal_12569 ;
    wire signal_12570 ;
    wire signal_12571 ;
    wire signal_12572 ;
    wire signal_12573 ;
    wire signal_12574 ;
    wire signal_12575 ;
    wire signal_12576 ;
    wire signal_12577 ;
    wire signal_12578 ;
    wire signal_12579 ;
    wire signal_12580 ;
    wire signal_12581 ;
    wire signal_12582 ;
    wire signal_12583 ;
    wire signal_12584 ;
    wire signal_12585 ;
    wire signal_12586 ;
    wire signal_12587 ;
    wire signal_12588 ;
    wire signal_12589 ;
    wire signal_12590 ;
    wire signal_12591 ;
    wire signal_12592 ;
    wire signal_12593 ;
    wire signal_12594 ;
    wire signal_12595 ;
    wire signal_12596 ;
    wire signal_12597 ;
    wire signal_12598 ;
    wire signal_12599 ;
    wire signal_12600 ;
    wire signal_12601 ;
    wire signal_12602 ;
    wire signal_12603 ;
    wire signal_12604 ;
    wire signal_12605 ;
    wire signal_12606 ;
    wire signal_12607 ;
    wire signal_12608 ;
    wire signal_12609 ;
    wire signal_12610 ;
    wire signal_12611 ;
    wire signal_12612 ;
    wire signal_12613 ;
    wire signal_12614 ;
    wire signal_12615 ;
    wire signal_12616 ;
    wire signal_12617 ;
    wire signal_12618 ;
    wire signal_12619 ;
    wire signal_12620 ;
    wire signal_12621 ;
    wire signal_12622 ;
    wire signal_12623 ;
    wire signal_12624 ;
    wire signal_12625 ;
    wire signal_12626 ;
    wire signal_12627 ;
    wire signal_12628 ;
    wire signal_12629 ;
    wire signal_12630 ;
    wire signal_12631 ;
    wire signal_12632 ;
    wire signal_12633 ;
    wire signal_12634 ;
    wire signal_12635 ;
    wire signal_12636 ;
    wire signal_12637 ;
    wire signal_12638 ;
    wire signal_12639 ;
    wire signal_12640 ;
    wire signal_12641 ;
    wire signal_12642 ;
    wire signal_12643 ;
    wire signal_12644 ;
    wire signal_12645 ;
    wire signal_12646 ;
    wire signal_12647 ;
    wire signal_12648 ;
    wire signal_12649 ;
    wire signal_12650 ;
    wire signal_12651 ;
    wire signal_12652 ;
    wire signal_12653 ;
    wire signal_12654 ;
    wire signal_12655 ;
    wire signal_12656 ;
    wire signal_12657 ;
    wire signal_12658 ;
    wire signal_12659 ;
    wire signal_12660 ;
    wire signal_12661 ;
    wire signal_12662 ;
    wire signal_12663 ;
    wire signal_12664 ;
    wire signal_12665 ;
    wire signal_12666 ;
    wire signal_12667 ;
    wire signal_12668 ;
    wire signal_12669 ;
    wire signal_12670 ;
    wire signal_12671 ;
    wire signal_12672 ;
    wire signal_12673 ;
    wire signal_12674 ;
    wire signal_12675 ;
    wire signal_12676 ;
    wire signal_12677 ;
    wire signal_12678 ;
    wire signal_12679 ;
    wire signal_12680 ;
    wire signal_12681 ;
    wire signal_12682 ;
    wire signal_12683 ;
    wire signal_12684 ;
    wire signal_12685 ;
    wire signal_12686 ;
    wire signal_12687 ;
    wire signal_12688 ;
    wire signal_12689 ;
    wire signal_12690 ;
    wire signal_12691 ;
    wire signal_12692 ;
    wire signal_12693 ;
    wire signal_12694 ;
    wire signal_12695 ;
    wire signal_12696 ;
    wire signal_12697 ;
    wire signal_12698 ;
    wire signal_12699 ;
    wire signal_12700 ;
    wire signal_12701 ;
    wire signal_12702 ;
    wire signal_12703 ;
    wire signal_12704 ;
    wire signal_12705 ;
    wire signal_12706 ;
    wire signal_12707 ;
    wire signal_12708 ;
    wire signal_12709 ;
    wire signal_12710 ;
    wire signal_12711 ;
    wire signal_12712 ;
    wire signal_12713 ;
    wire signal_12714 ;
    wire signal_12715 ;
    wire signal_12716 ;
    wire signal_12717 ;
    wire signal_12718 ;
    wire signal_12719 ;
    wire signal_12720 ;
    wire signal_12721 ;
    wire signal_12722 ;
    wire signal_12723 ;
    wire signal_12724 ;
    wire signal_12725 ;
    wire signal_12726 ;
    wire signal_12727 ;
    wire signal_12728 ;
    wire signal_12729 ;
    wire signal_12730 ;
    wire signal_12731 ;
    wire signal_12732 ;
    wire signal_12733 ;
    wire signal_12734 ;
    wire signal_12735 ;
    wire signal_12736 ;
    wire signal_12737 ;
    wire signal_12738 ;
    wire signal_12739 ;
    wire signal_12740 ;
    wire signal_12741 ;
    wire signal_12742 ;
    wire signal_12743 ;
    wire signal_12744 ;
    wire signal_12745 ;
    wire signal_12746 ;
    wire signal_12747 ;
    wire signal_12748 ;
    wire signal_12749 ;
    wire signal_12750 ;
    wire signal_12751 ;
    wire signal_12752 ;
    wire signal_12753 ;
    wire signal_12754 ;
    wire signal_12755 ;
    wire signal_12756 ;
    wire signal_12757 ;
    wire signal_12758 ;
    wire signal_12759 ;
    wire signal_12760 ;
    wire signal_12761 ;
    wire signal_12762 ;
    wire signal_12763 ;
    wire signal_12764 ;
    wire signal_12765 ;
    wire signal_12766 ;
    wire signal_12767 ;
    wire signal_12768 ;
    wire signal_12769 ;
    wire signal_12770 ;
    wire signal_12771 ;
    wire signal_12772 ;
    wire signal_12773 ;
    wire signal_12774 ;
    wire signal_12775 ;
    wire signal_12776 ;
    wire signal_12777 ;
    wire signal_12778 ;
    wire signal_12779 ;
    wire signal_12780 ;
    wire signal_12781 ;
    wire signal_12782 ;
    wire signal_12783 ;
    wire signal_12784 ;
    wire signal_12785 ;
    wire signal_12786 ;
    wire signal_12787 ;
    wire signal_12788 ;
    wire signal_12789 ;
    wire signal_12790 ;
    wire signal_12791 ;
    wire signal_12792 ;
    wire signal_12793 ;
    wire signal_12794 ;
    wire signal_12795 ;
    wire signal_12796 ;
    wire signal_12797 ;
    wire signal_12798 ;
    wire signal_12799 ;
    wire signal_12800 ;
    wire signal_12801 ;
    wire signal_12802 ;
    wire signal_12803 ;
    wire signal_12804 ;
    wire signal_12805 ;
    wire signal_12806 ;
    wire signal_12807 ;
    wire signal_12808 ;
    wire signal_12809 ;
    wire signal_12810 ;
    wire signal_12811 ;
    wire signal_12812 ;
    wire signal_12813 ;
    wire signal_12814 ;
    wire signal_12815 ;
    wire signal_12816 ;

    /* cells in depth 0 */
    AND2_X1 cell_0 ( .A1 (signal_396), .A2 (signal_395), .ZN (signal_393) ) ;
    NOR2_X1 cell_1 ( .A1 (signal_411), .A2 (signal_400), .ZN (signal_394) ) ;
    AND2_X1 cell_2 ( .A1 (signal_2273), .A2 (signal_394), .ZN (done) ) ;
    INV_X1 cell_3 ( .A (signal_2270), .ZN (signal_411) ) ;
    NOR2_X1 cell_4 ( .A1 (signal_2276), .A2 (signal_2275), .ZN (signal_396) ) ;
    INV_X1 cell_5 ( .A (signal_2271), .ZN (signal_397) ) ;
    NAND2_X1 cell_6 ( .A1 (signal_2272), .A2 (signal_397), .ZN (signal_400) ) ;
    NOR2_X1 cell_7 ( .A1 (done), .A2 (signal_2274), .ZN (signal_395) ) ;
    INV_X1 cell_8 ( .A (signal_2272), .ZN (signal_406) ) ;
    NAND2_X1 cell_9 ( .A1 (signal_406), .A2 (signal_397), .ZN (signal_398) ) ;
    NOR2_X1 cell_10 ( .A1 (signal_2273), .A2 (signal_398), .ZN (signal_2141) ) ;
    NOR2_X1 cell_11 ( .A1 (signal_2273), .A2 (signal_2270), .ZN (signal_409) ) ;
    NOR2_X1 cell_12 ( .A1 (signal_409), .A2 (signal_398), .ZN (signal_2140) ) ;
    NOR2_X1 cell_13 ( .A1 (signal_2270), .A2 (signal_400), .ZN (signal_399) ) ;
    NOR2_X1 cell_14 ( .A1 (signal_411), .A2 (signal_398), .ZN (signal_405) ) ;
    MUX2_X1 cell_15 ( .S (signal_2273), .A (signal_399), .B (signal_405), .Z (signal_2139) ) ;
    INV_X1 cell_16 ( .A (signal_2273), .ZN (signal_401) ) ;
    NOR2_X1 cell_17 ( .A1 (signal_401), .A2 (signal_400), .ZN (signal_402) ) ;
    MUX2_X1 cell_18 ( .S (signal_2270), .A (signal_402), .B (signal_2141), .Z (signal_2138) ) ;
    NAND2_X1 cell_19 ( .A1 (signal_2271), .A2 (signal_409), .ZN (signal_403) ) ;
    NOR2_X1 cell_20 ( .A1 (signal_2272), .A2 (signal_403), .ZN (signal_404) ) ;
    OR2_X1 cell_21 ( .A1 (signal_405), .A2 (signal_404), .ZN (signal_2137) ) ;
    XNOR2_X1 cell_22 ( .A (signal_2271), .B (signal_2270), .ZN (signal_408) ) ;
    NAND2_X1 cell_23 ( .A1 (signal_2273), .A2 (signal_406), .ZN (signal_407) ) ;
    NOR2_X1 cell_24 ( .A1 (signal_408), .A2 (signal_407), .ZN (signal_2136) ) ;
    INV_X1 cell_25 ( .A (signal_409), .ZN (signal_410) ) ;
    NAND2_X1 cell_26 ( .A1 (signal_2272), .A2 (signal_2271), .ZN (signal_412) ) ;
    NOR2_X1 cell_27 ( .A1 (signal_410), .A2 (signal_412), .ZN (signal_2135) ) ;
    NAND2_X1 cell_28 ( .A1 (signal_2273), .A2 (signal_411), .ZN (signal_413) ) ;
    NOR2_X1 cell_29 ( .A1 (signal_413), .A2 (signal_412), .ZN (signal_2134) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_30 ( .a ({ciphertext_s1[32], ciphertext_s0[32]}), .b ({signal_2339, signal_1793}), .c ({signal_2340, signal_1681}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_31 ( .a ({ciphertext_s1[4], ciphertext_s0[4]}), .b ({signal_2342, signal_2065}), .c ({signal_2343, signal_1709}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_32 ( .a ({ciphertext_s1[5], ciphertext_s0[5]}), .b ({signal_2345, signal_2064}), .c ({signal_2346, signal_1708}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_33 ( .a ({ciphertext_s1[6], ciphertext_s0[6]}), .b ({signal_2348, signal_2063}), .c ({signal_2349, signal_1707}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_34 ( .a ({ciphertext_s1[7], ciphertext_s0[7]}), .b ({signal_2351, signal_2062}), .c ({signal_2352, signal_1706}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_35 ( .a ({ciphertext_s1[40], ciphertext_s0[40]}), .b ({signal_2354, signal_2061}), .c ({signal_2355, signal_1737}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_36 ( .a ({ciphertext_s1[41], ciphertext_s0[41]}), .b ({signal_2357, signal_2060}), .c ({signal_2358, signal_1736}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_37 ( .a ({ciphertext_s1[42], ciphertext_s0[42]}), .b ({signal_2360, signal_2059}), .c ({signal_2361, signal_1735}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_38 ( .a ({ciphertext_s1[43], ciphertext_s0[43]}), .b ({signal_2363, signal_2058}), .c ({signal_2364, signal_1734}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_39 ( .a ({ciphertext_s1[44], ciphertext_s0[44]}), .b ({signal_2366, signal_2057}), .c ({signal_2367, signal_1733}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_40 ( .a ({ciphertext_s1[45], ciphertext_s0[45]}), .b ({signal_2369, signal_2056}), .c ({signal_2370, signal_1732}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_41 ( .a ({ciphertext_s1[74], ciphertext_s0[74]}), .b ({signal_2372, signal_1799}), .c ({signal_2373, signal_1703}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_42 ( .a ({ciphertext_s1[46], ciphertext_s0[46]}), .b ({signal_2375, signal_2055}), .c ({signal_2376, signal_1731}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_43 ( .a ({ciphertext_s1[47], ciphertext_s0[47]}), .b ({signal_2378, signal_2054}), .c ({signal_2379, signal_1730}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_44 ( .a ({ciphertext_s1[80], ciphertext_s0[80]}), .b ({signal_2381, signal_2053}), .c ({signal_2382, signal_1761}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_45 ( .a ({ciphertext_s1[81], ciphertext_s0[81]}), .b ({signal_2384, signal_2052}), .c ({signal_2385, signal_1760}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_46 ( .a ({ciphertext_s1[82], ciphertext_s0[82]}), .b ({signal_2387, signal_2051}), .c ({signal_2388, signal_1759}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_47 ( .a ({ciphertext_s1[83], ciphertext_s0[83]}), .b ({signal_2390, signal_2050}), .c ({signal_2391, signal_1758}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_48 ( .a ({ciphertext_s1[84], ciphertext_s0[84]}), .b ({signal_2393, signal_2049}), .c ({signal_2394, signal_1757}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_49 ( .a ({ciphertext_s1[85], ciphertext_s0[85]}), .b ({signal_2396, signal_2048}), .c ({signal_2397, signal_1756}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_50 ( .a ({ciphertext_s1[86], ciphertext_s0[86]}), .b ({signal_2399, signal_2047}), .c ({signal_2400, signal_1755}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_51 ( .a ({ciphertext_s1[87], ciphertext_s0[87]}), .b ({signal_2402, signal_2046}), .c ({signal_2403, signal_1754}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_52 ( .a ({ciphertext_s1[75], ciphertext_s0[75]}), .b ({signal_2405, signal_1798}), .c ({signal_2406, signal_1702}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_53 ( .a ({ciphertext_s1[120], ciphertext_s0[120]}), .b ({signal_2408, signal_2045}), .c ({signal_2409, signal_1657}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_54 ( .a ({ciphertext_s1[121], ciphertext_s0[121]}), .b ({signal_2411, signal_2044}), .c ({signal_2412, signal_1656}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_55 ( .a ({ciphertext_s1[122], ciphertext_s0[122]}), .b ({signal_2414, signal_2043}), .c ({signal_2415, signal_1655}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_56 ( .a ({ciphertext_s1[123], ciphertext_s0[123]}), .b ({signal_2417, signal_2042}), .c ({signal_2418, signal_1654}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_57 ( .a ({ciphertext_s1[124], ciphertext_s0[124]}), .b ({signal_2420, signal_2041}), .c ({signal_2421, signal_1653}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_58 ( .a ({ciphertext_s1[125], ciphertext_s0[125]}), .b ({signal_2423, signal_2040}), .c ({signal_2424, signal_1652}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_59 ( .a ({ciphertext_s1[126], ciphertext_s0[126]}), .b ({signal_2426, signal_2039}), .c ({signal_2427, signal_1651}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_60 ( .a ({ciphertext_s1[127], ciphertext_s0[127]}), .b ({signal_2429, signal_2038}), .c ({signal_2430, signal_1650}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_61 ( .a ({ciphertext_s1[76], ciphertext_s0[76]}), .b ({signal_2432, signal_1797}), .c ({signal_2433, signal_1701}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_62 ( .a ({ciphertext_s1[77], ciphertext_s0[77]}), .b ({signal_2435, signal_1796}), .c ({signal_2436, signal_1700}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_63 ( .a ({ciphertext_s1[78], ciphertext_s0[78]}), .b ({signal_2438, signal_1795}), .c ({signal_2439, signal_1699}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_64 ( .a ({ciphertext_s1[79], ciphertext_s0[79]}), .b ({signal_2441, signal_1794}), .c ({signal_2442, signal_1698}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_65 ( .a ({ciphertext_s1[112], ciphertext_s0[112]}), .b ({signal_2444, signal_1809}), .c ({signal_2445, signal_1729}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_66 ( .a ({ciphertext_s1[113], ciphertext_s0[113]}), .b ({signal_2447, signal_1808}), .c ({signal_2448, signal_1728}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_67 ( .a ({ciphertext_s1[114], ciphertext_s0[114]}), .b ({signal_2450, signal_1807}), .c ({signal_2451, signal_1727}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_68 ( .a ({ciphertext_s1[115], ciphertext_s0[115]}), .b ({signal_2453, signal_1806}), .c ({signal_2454, signal_1726}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_69 ( .a ({ciphertext_s1[33], ciphertext_s0[33]}), .b ({signal_2456, signal_1792}), .c ({signal_2457, signal_1680}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_70 ( .a ({ciphertext_s1[116], ciphertext_s0[116]}), .b ({signal_2459, signal_1805}), .c ({signal_2460, signal_1725}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_71 ( .a ({ciphertext_s1[117], ciphertext_s0[117]}), .b ({signal_2462, signal_1804}), .c ({signal_2463, signal_1724}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_72 ( .a ({ciphertext_s1[118], ciphertext_s0[118]}), .b ({signal_2465, signal_1803}), .c ({signal_2466, signal_1723}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_73 ( .a ({ciphertext_s1[119], ciphertext_s0[119]}), .b ({signal_2468, signal_1802}), .c ({signal_2469, signal_1722}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_74 ( .a ({ciphertext_s1[24], ciphertext_s0[24]}), .b ({signal_2471, signal_1785}), .c ({signal_2472, signal_1753}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_75 ( .a ({ciphertext_s1[25], ciphertext_s0[25]}), .b ({signal_2474, signal_1784}), .c ({signal_2475, signal_1752}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_76 ( .a ({ciphertext_s1[26], ciphertext_s0[26]}), .b ({signal_2477, signal_1783}), .c ({signal_2478, signal_1751}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_77 ( .a ({ciphertext_s1[27], ciphertext_s0[27]}), .b ({signal_2480, signal_1782}), .c ({signal_2481, signal_1750}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_78 ( .a ({ciphertext_s1[28], ciphertext_s0[28]}), .b ({signal_2483, signal_1781}), .c ({signal_2484, signal_1749}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_79 ( .a ({ciphertext_s1[29], ciphertext_s0[29]}), .b ({signal_2486, signal_1780}), .c ({signal_2487, signal_1748}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_80 ( .a ({ciphertext_s1[34], ciphertext_s0[34]}), .b ({signal_2489, signal_1791}), .c ({signal_2490, signal_1679}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_81 ( .a ({ciphertext_s1[30], ciphertext_s0[30]}), .b ({signal_2492, signal_1779}), .c ({signal_2493, signal_1747}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_82 ( .a ({ciphertext_s1[31], ciphertext_s0[31]}), .b ({signal_2495, signal_1778}), .c ({signal_2496, signal_1746}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_83 ( .a ({ciphertext_s1[64], ciphertext_s0[64]}), .b ({signal_2498, signal_2133}), .c ({signal_2499, signal_1777}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_84 ( .a ({ciphertext_s1[65], ciphertext_s0[65]}), .b ({signal_2501, signal_2132}), .c ({signal_2502, signal_1776}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_85 ( .a ({ciphertext_s1[66], ciphertext_s0[66]}), .b ({signal_2504, signal_2131}), .c ({signal_2505, signal_1775}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_86 ( .a ({ciphertext_s1[67], ciphertext_s0[67]}), .b ({signal_2507, signal_2130}), .c ({signal_2508, signal_1774}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_87 ( .a ({ciphertext_s1[68], ciphertext_s0[68]}), .b ({signal_2510, signal_2129}), .c ({signal_2511, signal_1773}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_88 ( .a ({ciphertext_s1[69], ciphertext_s0[69]}), .b ({signal_2513, signal_2128}), .c ({signal_2514, signal_1772}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_89 ( .a ({ciphertext_s1[70], ciphertext_s0[70]}), .b ({signal_2516, signal_2127}), .c ({signal_2517, signal_1771}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_90 ( .a ({ciphertext_s1[71], ciphertext_s0[71]}), .b ({signal_2519, signal_2126}), .c ({signal_2520, signal_1770}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_91 ( .a ({ciphertext_s1[35], ciphertext_s0[35]}), .b ({signal_2522, signal_1790}), .c ({signal_2523, signal_1678}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_92 ( .a ({ciphertext_s1[104], ciphertext_s0[104]}), .b ({signal_2525, signal_2125}), .c ({signal_2526, signal_1673}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_93 ( .a ({ciphertext_s1[105], ciphertext_s0[105]}), .b ({signal_2528, signal_2124}), .c ({signal_2529, signal_1672}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_94 ( .a ({ciphertext_s1[106], ciphertext_s0[106]}), .b ({signal_2531, signal_2123}), .c ({signal_2532, signal_1671}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_95 ( .a ({ciphertext_s1[107], ciphertext_s0[107]}), .b ({signal_2534, signal_2122}), .c ({signal_2535, signal_1670}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_96 ( .a ({ciphertext_s1[108], ciphertext_s0[108]}), .b ({signal_2537, signal_2121}), .c ({signal_2538, signal_1669}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_97 ( .a ({ciphertext_s1[109], ciphertext_s0[109]}), .b ({signal_2540, signal_2120}), .c ({signal_2541, signal_1668}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_98 ( .a ({ciphertext_s1[110], ciphertext_s0[110]}), .b ({signal_2543, signal_2119}), .c ({signal_2544, signal_1667}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_99 ( .a ({ciphertext_s1[111], ciphertext_s0[111]}), .b ({signal_2546, signal_2118}), .c ({signal_2547, signal_1666}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_100 ( .a ({ciphertext_s1[16], ciphertext_s0[16]}), .b ({signal_2549, signal_2117}), .c ({signal_2550, signal_1697}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_101 ( .a ({ciphertext_s1[17], ciphertext_s0[17]}), .b ({signal_2552, signal_2116}), .c ({signal_2553, signal_1696}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_102 ( .a ({ciphertext_s1[36], ciphertext_s0[36]}), .b ({signal_2555, signal_1789}), .c ({signal_2556, signal_1677}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_103 ( .a ({ciphertext_s1[18], ciphertext_s0[18]}), .b ({signal_2558, signal_2115}), .c ({signal_2559, signal_1695}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_104 ( .a ({ciphertext_s1[19], ciphertext_s0[19]}), .b ({signal_2561, signal_2114}), .c ({signal_2562, signal_1694}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_105 ( .a ({ciphertext_s1[20], ciphertext_s0[20]}), .b ({signal_2564, signal_2113}), .c ({signal_2565, signal_1693}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_106 ( .a ({ciphertext_s1[21], ciphertext_s0[21]}), .b ({signal_2567, signal_2112}), .c ({signal_2568, signal_1692}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_107 ( .a ({ciphertext_s1[22], ciphertext_s0[22]}), .b ({signal_2570, signal_2111}), .c ({signal_2571, signal_1691}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_108 ( .a ({ciphertext_s1[23], ciphertext_s0[23]}), .b ({signal_2573, signal_2110}), .c ({signal_2574, signal_1690}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_109 ( .a ({ciphertext_s1[56], ciphertext_s0[56]}), .b ({signal_2576, signal_2109}), .c ({signal_2577, signal_1721}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_110 ( .a ({ciphertext_s1[57], ciphertext_s0[57]}), .b ({signal_2579, signal_2108}), .c ({signal_2580, signal_1720}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_111 ( .a ({ciphertext_s1[58], ciphertext_s0[58]}), .b ({signal_2582, signal_2107}), .c ({signal_2583, signal_1719}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_112 ( .a ({ciphertext_s1[59], ciphertext_s0[59]}), .b ({signal_2585, signal_2106}), .c ({signal_2586, signal_1718}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_113 ( .a ({ciphertext_s1[37], ciphertext_s0[37]}), .b ({signal_2588, signal_1788}), .c ({signal_2589, signal_1676}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_114 ( .a ({ciphertext_s1[60], ciphertext_s0[60]}), .b ({signal_2591, signal_2105}), .c ({signal_2592, signal_1717}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_115 ( .a ({ciphertext_s1[61], ciphertext_s0[61]}), .b ({signal_2594, signal_2104}), .c ({signal_2595, signal_1716}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_116 ( .a ({ciphertext_s1[62], ciphertext_s0[62]}), .b ({signal_2597, signal_2103}), .c ({signal_2598, signal_1715}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_117 ( .a ({ciphertext_s1[63], ciphertext_s0[63]}), .b ({signal_2600, signal_2102}), .c ({signal_2601, signal_1714}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_118 ( .a ({ciphertext_s1[96], ciphertext_s0[96]}), .b ({signal_2603, signal_2101}), .c ({signal_2604, signal_1745}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_119 ( .a ({ciphertext_s1[97], ciphertext_s0[97]}), .b ({signal_2606, signal_2100}), .c ({signal_2607, signal_1744}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_120 ( .a ({ciphertext_s1[98], ciphertext_s0[98]}), .b ({signal_2609, signal_2099}), .c ({signal_2610, signal_1743}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_121 ( .a ({ciphertext_s1[99], ciphertext_s0[99]}), .b ({signal_2612, signal_2098}), .c ({signal_2613, signal_1742}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_122 ( .a ({ciphertext_s1[100], ciphertext_s0[100]}), .b ({signal_2615, signal_2097}), .c ({signal_2616, signal_1741}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_123 ( .a ({ciphertext_s1[101], ciphertext_s0[101]}), .b ({signal_2618, signal_2096}), .c ({signal_2619, signal_1740}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_124 ( .a ({ciphertext_s1[38], ciphertext_s0[38]}), .b ({signal_2621, signal_1787}), .c ({signal_2622, signal_1675}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_125 ( .a ({ciphertext_s1[102], ciphertext_s0[102]}), .b ({signal_2624, signal_2095}), .c ({signal_2625, signal_1739}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_126 ( .a ({ciphertext_s1[103], ciphertext_s0[103]}), .b ({signal_2627, signal_2094}), .c ({signal_2628, signal_1738}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_127 ( .a ({ciphertext_s1[8], ciphertext_s0[8]}), .b ({signal_2630, signal_2093}), .c ({signal_2631, signal_1769}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_128 ( .a ({ciphertext_s1[9], ciphertext_s0[9]}), .b ({signal_2633, signal_2092}), .c ({signal_2634, signal_1768}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_129 ( .a ({ciphertext_s1[10], ciphertext_s0[10]}), .b ({signal_2636, signal_2091}), .c ({signal_2637, signal_1767}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_130 ( .a ({ciphertext_s1[11], ciphertext_s0[11]}), .b ({signal_2639, signal_2090}), .c ({signal_2640, signal_1766}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_131 ( .a ({ciphertext_s1[12], ciphertext_s0[12]}), .b ({signal_2642, signal_2089}), .c ({signal_2643, signal_1765}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_132 ( .a ({ciphertext_s1[13], ciphertext_s0[13]}), .b ({signal_2645, signal_2088}), .c ({signal_2646, signal_1764}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_133 ( .a ({ciphertext_s1[14], ciphertext_s0[14]}), .b ({signal_2648, signal_2087}), .c ({signal_2649, signal_1763}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_134 ( .a ({ciphertext_s1[15], ciphertext_s0[15]}), .b ({signal_2651, signal_2086}), .c ({signal_2652, signal_1762}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_135 ( .a ({ciphertext_s1[39], ciphertext_s0[39]}), .b ({signal_2654, signal_1786}), .c ({signal_2655, signal_1674}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_136 ( .a ({ciphertext_s1[48], ciphertext_s0[48]}), .b ({signal_2657, signal_2085}), .c ({signal_2658, signal_1665}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_137 ( .a ({ciphertext_s1[49], ciphertext_s0[49]}), .b ({signal_2660, signal_2084}), .c ({signal_2661, signal_1664}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_138 ( .a ({ciphertext_s1[50], ciphertext_s0[50]}), .b ({signal_2663, signal_2083}), .c ({signal_2664, signal_1663}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_139 ( .a ({ciphertext_s1[51], ciphertext_s0[51]}), .b ({signal_2666, signal_2082}), .c ({signal_2667, signal_1662}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_140 ( .a ({ciphertext_s1[52], ciphertext_s0[52]}), .b ({signal_2669, signal_2081}), .c ({signal_2670, signal_1661}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_141 ( .a ({ciphertext_s1[53], ciphertext_s0[53]}), .b ({signal_2672, signal_2080}), .c ({signal_2673, signal_1660}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_142 ( .a ({ciphertext_s1[54], ciphertext_s0[54]}), .b ({signal_2675, signal_2079}), .c ({signal_2676, signal_1659}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_143 ( .a ({ciphertext_s1[55], ciphertext_s0[55]}), .b ({signal_2678, signal_2078}), .c ({signal_2679, signal_1658}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_144 ( .a ({ciphertext_s1[88], ciphertext_s0[88]}), .b ({signal_2681, signal_2077}), .c ({signal_2682, signal_1689}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_145 ( .a ({ciphertext_s1[89], ciphertext_s0[89]}), .b ({signal_2684, signal_2076}), .c ({signal_2685, signal_1688}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_146 ( .a ({ciphertext_s1[72], ciphertext_s0[72]}), .b ({signal_2687, signal_1801}), .c ({signal_2688, signal_1705}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_147 ( .a ({ciphertext_s1[90], ciphertext_s0[90]}), .b ({signal_2690, signal_2075}), .c ({signal_2691, signal_1687}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_148 ( .a ({ciphertext_s1[91], ciphertext_s0[91]}), .b ({signal_2693, signal_2074}), .c ({signal_2694, signal_1686}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_149 ( .a ({ciphertext_s1[92], ciphertext_s0[92]}), .b ({signal_2696, signal_2073}), .c ({signal_2697, signal_1685}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_150 ( .a ({ciphertext_s1[93], ciphertext_s0[93]}), .b ({signal_2699, signal_2072}), .c ({signal_2700, signal_1684}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_151 ( .a ({ciphertext_s1[94], ciphertext_s0[94]}), .b ({signal_2702, signal_2071}), .c ({signal_2703, signal_1683}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_152 ( .a ({ciphertext_s1[95], ciphertext_s0[95]}), .b ({signal_2705, signal_2070}), .c ({signal_2706, signal_1682}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_153 ( .a ({ciphertext_s1[0], ciphertext_s0[0]}), .b ({signal_2708, signal_2069}), .c ({signal_2709, signal_1713}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_154 ( .a ({ciphertext_s1[1], ciphertext_s0[1]}), .b ({signal_2711, signal_2068}), .c ({signal_2712, signal_1712}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_155 ( .a ({ciphertext_s1[2], ciphertext_s0[2]}), .b ({signal_2714, signal_2067}), .c ({signal_2715, signal_1711}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_156 ( .a ({ciphertext_s1[3], ciphertext_s0[3]}), .b ({signal_2717, signal_2066}), .c ({signal_2718, signal_1710}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_157 ( .a ({ciphertext_s1[73], ciphertext_s0[73]}), .b ({signal_2720, signal_1800}), .c ({signal_2721, signal_1704}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_256 ( .s (reset), .b ({signal_2754, signal_1617}), .a ({plaintext_s1[32], plaintext_s0[32]}), .c ({signal_2851, signal_478}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_259 ( .s (reset), .b ({signal_2755, signal_1616}), .a ({plaintext_s1[33], plaintext_s0[33]}), .c ({signal_2853, signal_480}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_262 ( .s (reset), .b ({signal_2756, signal_1615}), .a ({plaintext_s1[34], plaintext_s0[34]}), .c ({signal_2855, signal_482}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_265 ( .s (reset), .b ({signal_2757, signal_1614}), .a ({plaintext_s1[35], plaintext_s0[35]}), .c ({signal_2857, signal_484}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_268 ( .s (reset), .b ({signal_2758, signal_1613}), .a ({plaintext_s1[36], plaintext_s0[36]}), .c ({signal_2859, signal_486}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_271 ( .s (reset), .b ({signal_2759, signal_1612}), .a ({plaintext_s1[37], plaintext_s0[37]}), .c ({signal_2861, signal_488}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_274 ( .s (reset), .b ({signal_2760, signal_1611}), .a ({plaintext_s1[38], plaintext_s0[38]}), .c ({signal_2863, signal_490}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_277 ( .s (reset), .b ({signal_2761, signal_1610}), .a ({plaintext_s1[39], plaintext_s0[39]}), .c ({signal_2865, signal_492}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_280 ( .s (reset), .b ({signal_2762, signal_1609}), .a ({plaintext_s1[40], plaintext_s0[40]}), .c ({signal_2867, signal_494}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_283 ( .s (reset), .b ({signal_2763, signal_1608}), .a ({plaintext_s1[41], plaintext_s0[41]}), .c ({signal_2869, signal_496}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_286 ( .s (reset), .b ({signal_2764, signal_1607}), .a ({plaintext_s1[42], plaintext_s0[42]}), .c ({signal_2871, signal_498}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_289 ( .s (reset), .b ({signal_2765, signal_1606}), .a ({plaintext_s1[43], plaintext_s0[43]}), .c ({signal_2873, signal_500}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_292 ( .s (reset), .b ({signal_2766, signal_1605}), .a ({plaintext_s1[44], plaintext_s0[44]}), .c ({signal_2875, signal_502}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_295 ( .s (reset), .b ({signal_2767, signal_1604}), .a ({plaintext_s1[45], plaintext_s0[45]}), .c ({signal_2877, signal_504}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_298 ( .s (reset), .b ({signal_2768, signal_1603}), .a ({plaintext_s1[46], plaintext_s0[46]}), .c ({signal_2879, signal_506}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_301 ( .s (reset), .b ({signal_2769, signal_1602}), .a ({plaintext_s1[47], plaintext_s0[47]}), .c ({signal_2881, signal_508}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_304 ( .s (reset), .b ({signal_2770, signal_1601}), .a ({plaintext_s1[48], plaintext_s0[48]}), .c ({signal_2883, signal_510}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_307 ( .s (reset), .b ({signal_2771, signal_1600}), .a ({plaintext_s1[49], plaintext_s0[49]}), .c ({signal_2885, signal_512}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_310 ( .s (reset), .b ({signal_2772, signal_1599}), .a ({plaintext_s1[50], plaintext_s0[50]}), .c ({signal_2887, signal_514}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_313 ( .s (reset), .b ({signal_2773, signal_1598}), .a ({plaintext_s1[51], plaintext_s0[51]}), .c ({signal_2889, signal_516}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_316 ( .s (reset), .b ({signal_2774, signal_1597}), .a ({plaintext_s1[52], plaintext_s0[52]}), .c ({signal_2891, signal_518}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_319 ( .s (reset), .b ({signal_2775, signal_1596}), .a ({plaintext_s1[53], plaintext_s0[53]}), .c ({signal_2893, signal_520}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_322 ( .s (reset), .b ({signal_2776, signal_1595}), .a ({plaintext_s1[54], plaintext_s0[54]}), .c ({signal_2895, signal_522}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_325 ( .s (reset), .b ({signal_2777, signal_1594}), .a ({plaintext_s1[55], plaintext_s0[55]}), .c ({signal_2897, signal_524}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_328 ( .s (reset), .b ({signal_2778, signal_1593}), .a ({plaintext_s1[56], plaintext_s0[56]}), .c ({signal_2899, signal_526}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_331 ( .s (reset), .b ({signal_2779, signal_1592}), .a ({plaintext_s1[57], plaintext_s0[57]}), .c ({signal_2901, signal_528}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_334 ( .s (reset), .b ({signal_2780, signal_1591}), .a ({plaintext_s1[58], plaintext_s0[58]}), .c ({signal_2903, signal_530}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_337 ( .s (reset), .b ({signal_2781, signal_1590}), .a ({plaintext_s1[59], plaintext_s0[59]}), .c ({signal_2905, signal_532}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_340 ( .s (reset), .b ({signal_2782, signal_1589}), .a ({plaintext_s1[60], plaintext_s0[60]}), .c ({signal_2907, signal_534}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_343 ( .s (reset), .b ({signal_2783, signal_1588}), .a ({plaintext_s1[61], plaintext_s0[61]}), .c ({signal_2909, signal_536}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_346 ( .s (reset), .b ({signal_2784, signal_1587}), .a ({plaintext_s1[62], plaintext_s0[62]}), .c ({signal_2911, signal_538}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_349 ( .s (reset), .b ({signal_2785, signal_1586}), .a ({plaintext_s1[63], plaintext_s0[63]}), .c ({signal_2913, signal_540}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_352 ( .s (reset), .b ({signal_2786, signal_1585}), .a ({plaintext_s1[64], plaintext_s0[64]}), .c ({signal_2915, signal_542}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_355 ( .s (reset), .b ({signal_2787, signal_1584}), .a ({plaintext_s1[65], plaintext_s0[65]}), .c ({signal_2917, signal_544}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_358 ( .s (reset), .b ({signal_2788, signal_1583}), .a ({plaintext_s1[66], plaintext_s0[66]}), .c ({signal_2919, signal_546}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_361 ( .s (reset), .b ({signal_2789, signal_1582}), .a ({plaintext_s1[67], plaintext_s0[67]}), .c ({signal_2921, signal_548}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_364 ( .s (reset), .b ({signal_2790, signal_1581}), .a ({plaintext_s1[68], plaintext_s0[68]}), .c ({signal_2923, signal_550}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_367 ( .s (reset), .b ({signal_2791, signal_1580}), .a ({plaintext_s1[69], plaintext_s0[69]}), .c ({signal_2925, signal_552}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_370 ( .s (reset), .b ({signal_2792, signal_1579}), .a ({plaintext_s1[70], plaintext_s0[70]}), .c ({signal_2927, signal_554}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_373 ( .s (reset), .b ({signal_2793, signal_1578}), .a ({plaintext_s1[71], plaintext_s0[71]}), .c ({signal_2929, signal_556}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_376 ( .s (reset), .b ({signal_2794, signal_1577}), .a ({plaintext_s1[72], plaintext_s0[72]}), .c ({signal_2931, signal_558}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_379 ( .s (reset), .b ({signal_2795, signal_1576}), .a ({plaintext_s1[73], plaintext_s0[73]}), .c ({signal_2933, signal_560}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_382 ( .s (reset), .b ({signal_2796, signal_1575}), .a ({plaintext_s1[74], plaintext_s0[74]}), .c ({signal_2935, signal_562}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_385 ( .s (reset), .b ({signal_2797, signal_1574}), .a ({plaintext_s1[75], plaintext_s0[75]}), .c ({signal_2937, signal_564}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_388 ( .s (reset), .b ({signal_2798, signal_1573}), .a ({plaintext_s1[76], plaintext_s0[76]}), .c ({signal_2939, signal_566}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_391 ( .s (reset), .b ({signal_2799, signal_1572}), .a ({plaintext_s1[77], plaintext_s0[77]}), .c ({signal_2941, signal_568}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_394 ( .s (reset), .b ({signal_2800, signal_1571}), .a ({plaintext_s1[78], plaintext_s0[78]}), .c ({signal_2943, signal_570}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_397 ( .s (reset), .b ({signal_2801, signal_1570}), .a ({plaintext_s1[79], plaintext_s0[79]}), .c ({signal_2945, signal_572}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_400 ( .s (reset), .b ({signal_2802, signal_1569}), .a ({plaintext_s1[80], plaintext_s0[80]}), .c ({signal_2947, signal_574}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_403 ( .s (reset), .b ({signal_2803, signal_1568}), .a ({plaintext_s1[81], plaintext_s0[81]}), .c ({signal_2949, signal_576}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_406 ( .s (reset), .b ({signal_2804, signal_1567}), .a ({plaintext_s1[82], plaintext_s0[82]}), .c ({signal_2951, signal_578}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_409 ( .s (reset), .b ({signal_2805, signal_1566}), .a ({plaintext_s1[83], plaintext_s0[83]}), .c ({signal_2953, signal_580}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_412 ( .s (reset), .b ({signal_2806, signal_1565}), .a ({plaintext_s1[84], plaintext_s0[84]}), .c ({signal_2955, signal_582}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_415 ( .s (reset), .b ({signal_2807, signal_1564}), .a ({plaintext_s1[85], plaintext_s0[85]}), .c ({signal_2957, signal_584}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_418 ( .s (reset), .b ({signal_2808, signal_1563}), .a ({plaintext_s1[86], plaintext_s0[86]}), .c ({signal_2959, signal_586}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_421 ( .s (reset), .b ({signal_2809, signal_1562}), .a ({plaintext_s1[87], plaintext_s0[87]}), .c ({signal_2961, signal_588}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_424 ( .s (reset), .b ({signal_2810, signal_1561}), .a ({plaintext_s1[88], plaintext_s0[88]}), .c ({signal_2963, signal_590}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_427 ( .s (reset), .b ({signal_2811, signal_1560}), .a ({plaintext_s1[89], plaintext_s0[89]}), .c ({signal_2965, signal_592}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_430 ( .s (reset), .b ({signal_2812, signal_1559}), .a ({plaintext_s1[90], plaintext_s0[90]}), .c ({signal_2967, signal_594}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_433 ( .s (reset), .b ({signal_2813, signal_1558}), .a ({plaintext_s1[91], plaintext_s0[91]}), .c ({signal_2969, signal_596}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_436 ( .s (reset), .b ({signal_2814, signal_1557}), .a ({plaintext_s1[92], plaintext_s0[92]}), .c ({signal_2971, signal_598}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_439 ( .s (reset), .b ({signal_2815, signal_1556}), .a ({plaintext_s1[93], plaintext_s0[93]}), .c ({signal_2973, signal_600}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_442 ( .s (reset), .b ({signal_2816, signal_1555}), .a ({plaintext_s1[94], plaintext_s0[94]}), .c ({signal_2975, signal_602}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_445 ( .s (reset), .b ({signal_2817, signal_1554}), .a ({plaintext_s1[95], plaintext_s0[95]}), .c ({signal_2977, signal_604}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_448 ( .s (reset), .b ({signal_2818, signal_1553}), .a ({plaintext_s1[96], plaintext_s0[96]}), .c ({signal_2979, signal_606}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_451 ( .s (reset), .b ({signal_2819, signal_1552}), .a ({plaintext_s1[97], plaintext_s0[97]}), .c ({signal_2981, signal_608}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_454 ( .s (reset), .b ({signal_2820, signal_1551}), .a ({plaintext_s1[98], plaintext_s0[98]}), .c ({signal_2983, signal_610}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_457 ( .s (reset), .b ({signal_2821, signal_1550}), .a ({plaintext_s1[99], plaintext_s0[99]}), .c ({signal_2985, signal_612}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_460 ( .s (reset), .b ({signal_2822, signal_1549}), .a ({plaintext_s1[100], plaintext_s0[100]}), .c ({signal_2987, signal_614}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_463 ( .s (reset), .b ({signal_2823, signal_1548}), .a ({plaintext_s1[101], plaintext_s0[101]}), .c ({signal_2989, signal_616}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_466 ( .s (reset), .b ({signal_2824, signal_1547}), .a ({plaintext_s1[102], plaintext_s0[102]}), .c ({signal_2991, signal_618}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_469 ( .s (reset), .b ({signal_2825, signal_1546}), .a ({plaintext_s1[103], plaintext_s0[103]}), .c ({signal_2993, signal_620}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_472 ( .s (reset), .b ({signal_2826, signal_1545}), .a ({plaintext_s1[104], plaintext_s0[104]}), .c ({signal_2995, signal_622}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_475 ( .s (reset), .b ({signal_2827, signal_1544}), .a ({plaintext_s1[105], plaintext_s0[105]}), .c ({signal_2997, signal_624}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_478 ( .s (reset), .b ({signal_2828, signal_1543}), .a ({plaintext_s1[106], plaintext_s0[106]}), .c ({signal_2999, signal_626}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_481 ( .s (reset), .b ({signal_2829, signal_1542}), .a ({plaintext_s1[107], plaintext_s0[107]}), .c ({signal_3001, signal_628}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_484 ( .s (reset), .b ({signal_2830, signal_1541}), .a ({plaintext_s1[108], plaintext_s0[108]}), .c ({signal_3003, signal_630}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_487 ( .s (reset), .b ({signal_2831, signal_1540}), .a ({plaintext_s1[109], plaintext_s0[109]}), .c ({signal_3005, signal_632}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_490 ( .s (reset), .b ({signal_2832, signal_1539}), .a ({plaintext_s1[110], plaintext_s0[110]}), .c ({signal_3007, signal_634}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_493 ( .s (reset), .b ({signal_2833, signal_1538}), .a ({plaintext_s1[111], plaintext_s0[111]}), .c ({signal_3009, signal_636}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_496 ( .s (reset), .b ({signal_2834, signal_1537}), .a ({plaintext_s1[112], plaintext_s0[112]}), .c ({signal_3011, signal_638}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_499 ( .s (reset), .b ({signal_2835, signal_1536}), .a ({plaintext_s1[113], plaintext_s0[113]}), .c ({signal_3013, signal_640}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_502 ( .s (reset), .b ({signal_2836, signal_1535}), .a ({plaintext_s1[114], plaintext_s0[114]}), .c ({signal_3015, signal_642}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_505 ( .s (reset), .b ({signal_2837, signal_1534}), .a ({plaintext_s1[115], plaintext_s0[115]}), .c ({signal_3017, signal_644}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_508 ( .s (reset), .b ({signal_2838, signal_1533}), .a ({plaintext_s1[116], plaintext_s0[116]}), .c ({signal_3019, signal_646}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_511 ( .s (reset), .b ({signal_2839, signal_1532}), .a ({plaintext_s1[117], plaintext_s0[117]}), .c ({signal_3021, signal_648}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_514 ( .s (reset), .b ({signal_2840, signal_1531}), .a ({plaintext_s1[118], plaintext_s0[118]}), .c ({signal_3023, signal_650}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_517 ( .s (reset), .b ({signal_2841, signal_1530}), .a ({plaintext_s1[119], plaintext_s0[119]}), .c ({signal_3025, signal_652}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_520 ( .s (reset), .b ({signal_2842, signal_1529}), .a ({plaintext_s1[120], plaintext_s0[120]}), .c ({signal_3027, signal_654}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_523 ( .s (reset), .b ({signal_2843, signal_1528}), .a ({plaintext_s1[121], plaintext_s0[121]}), .c ({signal_3029, signal_656}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_526 ( .s (reset), .b ({signal_2844, signal_1527}), .a ({plaintext_s1[122], plaintext_s0[122]}), .c ({signal_3031, signal_658}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_529 ( .s (reset), .b ({signal_2845, signal_1526}), .a ({plaintext_s1[123], plaintext_s0[123]}), .c ({signal_3033, signal_660}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_532 ( .s (reset), .b ({signal_2846, signal_1525}), .a ({plaintext_s1[124], plaintext_s0[124]}), .c ({signal_3035, signal_662}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_535 ( .s (reset), .b ({signal_2847, signal_1524}), .a ({plaintext_s1[125], plaintext_s0[125]}), .c ({signal_3037, signal_664}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_538 ( .s (reset), .b ({signal_2848, signal_1523}), .a ({plaintext_s1[126], plaintext_s0[126]}), .c ({signal_3039, signal_666}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_541 ( .s (reset), .b ({signal_2849, signal_1522}), .a ({plaintext_s1[127], plaintext_s0[127]}), .c ({signal_3041, signal_668}) ) ;
    INV_X1 cell_542 ( .A (signal_393), .ZN (signal_670) ) ;
    INV_X1 cell_543 ( .A (signal_670), .ZN (signal_672) ) ;
    INV_X1 cell_544 ( .A (signal_670), .ZN (signal_671) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_545 ( .s (signal_671), .b ({ciphertext_s1[0], ciphertext_s0[0]}), .a ({signal_2444, signal_1809}), .c ({signal_2723, signal_1841}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_546 ( .s (signal_671), .b ({ciphertext_s1[1], ciphertext_s0[1]}), .a ({signal_2447, signal_1808}), .c ({signal_2724, signal_1840}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_547 ( .s (signal_671), .b ({ciphertext_s1[2], ciphertext_s0[2]}), .a ({signal_2450, signal_1807}), .c ({signal_2725, signal_1839}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_548 ( .s (signal_671), .b ({ciphertext_s1[3], ciphertext_s0[3]}), .a ({signal_2453, signal_1806}), .c ({signal_2726, signal_1838}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_549 ( .s (signal_671), .b ({ciphertext_s1[4], ciphertext_s0[4]}), .a ({signal_2459, signal_1805}), .c ({signal_2727, signal_1837}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_550 ( .s (signal_671), .b ({ciphertext_s1[5], ciphertext_s0[5]}), .a ({signal_2462, signal_1804}), .c ({signal_2728, signal_1836}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_551 ( .s (signal_671), .b ({ciphertext_s1[6], ciphertext_s0[6]}), .a ({signal_2465, signal_1803}), .c ({signal_2729, signal_1835}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_552 ( .s (signal_671), .b ({ciphertext_s1[7], ciphertext_s0[7]}), .a ({signal_2468, signal_1802}), .c ({signal_2730, signal_1834}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_553 ( .s (signal_393), .b ({ciphertext_s1[40], ciphertext_s0[40]}), .a ({signal_2687, signal_1801}), .c ({signal_2722, signal_1833}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_554 ( .s (signal_672), .b ({ciphertext_s1[41], ciphertext_s0[41]}), .a ({signal_2720, signal_1800}), .c ({signal_2731, signal_1832}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_555 ( .s (signal_672), .b ({ciphertext_s1[42], ciphertext_s0[42]}), .a ({signal_2372, signal_1799}), .c ({signal_2732, signal_1831}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_556 ( .s (signal_672), .b ({ciphertext_s1[43], ciphertext_s0[43]}), .a ({signal_2405, signal_1798}), .c ({signal_2733, signal_1830}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_557 ( .s (signal_672), .b ({ciphertext_s1[44], ciphertext_s0[44]}), .a ({signal_2432, signal_1797}), .c ({signal_2734, signal_1829}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_558 ( .s (signal_671), .b ({ciphertext_s1[45], ciphertext_s0[45]}), .a ({signal_2435, signal_1796}), .c ({signal_2735, signal_1828}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_559 ( .s (signal_671), .b ({ciphertext_s1[46], ciphertext_s0[46]}), .a ({signal_2438, signal_1795}), .c ({signal_2736, signal_1827}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_560 ( .s (signal_672), .b ({ciphertext_s1[47], ciphertext_s0[47]}), .a ({signal_2441, signal_1794}), .c ({signal_2737, signal_1826}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_561 ( .s (signal_671), .b ({ciphertext_s1[80], ciphertext_s0[80]}), .a ({signal_2339, signal_1793}), .c ({signal_2738, signal_1825}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_562 ( .s (signal_672), .b ({ciphertext_s1[81], ciphertext_s0[81]}), .a ({signal_2456, signal_1792}), .c ({signal_2739, signal_1824}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_563 ( .s (signal_672), .b ({ciphertext_s1[82], ciphertext_s0[82]}), .a ({signal_2489, signal_1791}), .c ({signal_2740, signal_1823}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_564 ( .s (signal_672), .b ({ciphertext_s1[83], ciphertext_s0[83]}), .a ({signal_2522, signal_1790}), .c ({signal_2741, signal_1822}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_565 ( .s (signal_672), .b ({ciphertext_s1[84], ciphertext_s0[84]}), .a ({signal_2555, signal_1789}), .c ({signal_2742, signal_1821}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_566 ( .s (signal_672), .b ({ciphertext_s1[85], ciphertext_s0[85]}), .a ({signal_2588, signal_1788}), .c ({signal_2743, signal_1820}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_567 ( .s (signal_672), .b ({ciphertext_s1[86], ciphertext_s0[86]}), .a ({signal_2621, signal_1787}), .c ({signal_2744, signal_1819}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_568 ( .s (signal_672), .b ({ciphertext_s1[87], ciphertext_s0[87]}), .a ({signal_2654, signal_1786}), .c ({signal_2745, signal_1818}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_569 ( .s (signal_672), .b ({ciphertext_s1[120], ciphertext_s0[120]}), .a ({signal_2471, signal_1785}), .c ({signal_2746, signal_1817}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_570 ( .s (signal_672), .b ({ciphertext_s1[121], ciphertext_s0[121]}), .a ({signal_2474, signal_1784}), .c ({signal_2747, signal_1816}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_571 ( .s (signal_672), .b ({ciphertext_s1[122], ciphertext_s0[122]}), .a ({signal_2477, signal_1783}), .c ({signal_2748, signal_1815}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_572 ( .s (signal_672), .b ({ciphertext_s1[123], ciphertext_s0[123]}), .a ({signal_2480, signal_1782}), .c ({signal_2749, signal_1814}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_573 ( .s (signal_672), .b ({ciphertext_s1[124], ciphertext_s0[124]}), .a ({signal_2483, signal_1781}), .c ({signal_2750, signal_1813}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_574 ( .s (signal_672), .b ({ciphertext_s1[125], ciphertext_s0[125]}), .a ({signal_2486, signal_1780}), .c ({signal_2751, signal_1812}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_575 ( .s (signal_672), .b ({ciphertext_s1[126], ciphertext_s0[126]}), .a ({signal_2492, signal_1779}), .c ({signal_2752, signal_1811}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_576 ( .s (signal_672), .b ({ciphertext_s1[127], ciphertext_s0[127]}), .a ({signal_2495, signal_1778}), .c ({signal_2753, signal_1810}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_581 ( .a ({signal_2726, signal_1838}), .b ({signal_2724, signal_1840}), .c ({signal_3042, signal_788}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_709 ( .a ({signal_2733, signal_1830}), .b ({signal_2731, signal_1832}), .c ({signal_3043, signal_908}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_837 ( .a ({signal_2741, signal_1822}), .b ({signal_2739, signal_1824}), .c ({signal_3044, signal_1028}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_965 ( .a ({signal_2749, signal_1814}), .b ({signal_2747, signal_1816}), .c ({signal_3045, signal_1148}) ) ;
    INV_X1 cell_1197 ( .A (signal_394), .ZN (signal_1217) ) ;
    INV_X1 cell_1198 ( .A (signal_1217), .ZN (signal_1218) ) ;
    INV_X1 cell_1199 ( .A (signal_1217), .ZN (signal_1219) ) ;
    INV_X1 cell_1232 ( .A (signal_393), .ZN (signal_1220) ) ;
    INV_X1 cell_1233 ( .A (signal_1220), .ZN (signal_1223) ) ;
    INV_X1 cell_1234 ( .A (signal_1220), .ZN (signal_1225) ) ;
    INV_X1 cell_1235 ( .A (signal_1220), .ZN (signal_1226) ) ;
    INV_X1 cell_1236 ( .A (signal_1220), .ZN (signal_1224) ) ;
    INV_X1 cell_1237 ( .A (signal_1220), .ZN (signal_1221) ) ;
    INV_X1 cell_1238 ( .A (signal_1220), .ZN (signal_1222) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1271 ( .s (signal_1221), .b ({ciphertext_s1[32], ciphertext_s0[32]}), .a ({signal_2604, signal_1745}), .c ({signal_2754, signal_1617}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1272 ( .s (signal_1222), .b ({ciphertext_s1[33], ciphertext_s0[33]}), .a ({signal_2607, signal_1744}), .c ({signal_2755, signal_1616}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1273 ( .s (signal_1226), .b ({ciphertext_s1[34], ciphertext_s0[34]}), .a ({signal_2610, signal_1743}), .c ({signal_2756, signal_1615}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1274 ( .s (signal_1225), .b ({ciphertext_s1[35], ciphertext_s0[35]}), .a ({signal_2613, signal_1742}), .c ({signal_2757, signal_1614}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1275 ( .s (signal_1224), .b ({ciphertext_s1[36], ciphertext_s0[36]}), .a ({signal_2616, signal_1741}), .c ({signal_2758, signal_1613}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1276 ( .s (signal_1223), .b ({ciphertext_s1[37], ciphertext_s0[37]}), .a ({signal_2619, signal_1740}), .c ({signal_2759, signal_1612}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1277 ( .s (signal_1222), .b ({ciphertext_s1[38], ciphertext_s0[38]}), .a ({signal_2625, signal_1739}), .c ({signal_2760, signal_1611}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1278 ( .s (signal_1221), .b ({ciphertext_s1[39], ciphertext_s0[39]}), .a ({signal_2628, signal_1738}), .c ({signal_2761, signal_1610}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1279 ( .s (signal_1221), .b ({ciphertext_s1[72], ciphertext_s0[72]}), .a ({signal_2355, signal_1737}), .c ({signal_2762, signal_1609}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1280 ( .s (signal_1226), .b ({ciphertext_s1[73], ciphertext_s0[73]}), .a ({signal_2358, signal_1736}), .c ({signal_2763, signal_1608}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1281 ( .s (signal_1225), .b ({ciphertext_s1[74], ciphertext_s0[74]}), .a ({signal_2361, signal_1735}), .c ({signal_2764, signal_1607}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1282 ( .s (signal_1224), .b ({ciphertext_s1[75], ciphertext_s0[75]}), .a ({signal_2364, signal_1734}), .c ({signal_2765, signal_1606}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1283 ( .s (signal_1226), .b ({ciphertext_s1[76], ciphertext_s0[76]}), .a ({signal_2367, signal_1733}), .c ({signal_2766, signal_1605}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1284 ( .s (signal_1225), .b ({ciphertext_s1[77], ciphertext_s0[77]}), .a ({signal_2370, signal_1732}), .c ({signal_2767, signal_1604}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1285 ( .s (signal_1224), .b ({ciphertext_s1[78], ciphertext_s0[78]}), .a ({signal_2376, signal_1731}), .c ({signal_2768, signal_1603}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1286 ( .s (signal_1223), .b ({ciphertext_s1[79], ciphertext_s0[79]}), .a ({signal_2379, signal_1730}), .c ({signal_2769, signal_1602}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1287 ( .s (signal_1222), .b ({ciphertext_s1[112], ciphertext_s0[112]}), .a ({signal_2445, signal_1729}), .c ({signal_2770, signal_1601}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1288 ( .s (signal_1221), .b ({ciphertext_s1[113], ciphertext_s0[113]}), .a ({signal_2448, signal_1728}), .c ({signal_2771, signal_1600}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1289 ( .s (signal_1226), .b ({ciphertext_s1[114], ciphertext_s0[114]}), .a ({signal_2451, signal_1727}), .c ({signal_2772, signal_1599}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1290 ( .s (signal_1225), .b ({ciphertext_s1[115], ciphertext_s0[115]}), .a ({signal_2454, signal_1726}), .c ({signal_2773, signal_1598}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1291 ( .s (signal_1224), .b ({ciphertext_s1[116], ciphertext_s0[116]}), .a ({signal_2460, signal_1725}), .c ({signal_2774, signal_1597}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1292 ( .s (signal_1223), .b ({ciphertext_s1[117], ciphertext_s0[117]}), .a ({signal_2463, signal_1724}), .c ({signal_2775, signal_1596}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1293 ( .s (signal_1222), .b ({ciphertext_s1[118], ciphertext_s0[118]}), .a ({signal_2466, signal_1723}), .c ({signal_2776, signal_1595}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1294 ( .s (signal_1221), .b ({ciphertext_s1[119], ciphertext_s0[119]}), .a ({signal_2469, signal_1722}), .c ({signal_2777, signal_1594}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1295 ( .s (signal_1221), .b ({ciphertext_s1[24], ciphertext_s0[24]}), .a ({signal_2577, signal_1721}), .c ({signal_2778, signal_1593}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1296 ( .s (signal_1221), .b ({ciphertext_s1[25], ciphertext_s0[25]}), .a ({signal_2580, signal_1720}), .c ({signal_2779, signal_1592}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1297 ( .s (signal_1221), .b ({ciphertext_s1[26], ciphertext_s0[26]}), .a ({signal_2583, signal_1719}), .c ({signal_2780, signal_1591}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1298 ( .s (signal_1221), .b ({ciphertext_s1[27], ciphertext_s0[27]}), .a ({signal_2586, signal_1718}), .c ({signal_2781, signal_1590}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1299 ( .s (signal_1221), .b ({ciphertext_s1[28], ciphertext_s0[28]}), .a ({signal_2592, signal_1717}), .c ({signal_2782, signal_1589}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1300 ( .s (signal_1221), .b ({ciphertext_s1[29], ciphertext_s0[29]}), .a ({signal_2595, signal_1716}), .c ({signal_2783, signal_1588}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1301 ( .s (signal_1221), .b ({ciphertext_s1[30], ciphertext_s0[30]}), .a ({signal_2598, signal_1715}), .c ({signal_2784, signal_1587}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1302 ( .s (signal_1221), .b ({ciphertext_s1[31], ciphertext_s0[31]}), .a ({signal_2601, signal_1714}), .c ({signal_2785, signal_1586}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1303 ( .s (signal_1221), .b ({ciphertext_s1[64], ciphertext_s0[64]}), .a ({signal_2709, signal_1713}), .c ({signal_2786, signal_1585}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1304 ( .s (signal_1221), .b ({ciphertext_s1[65], ciphertext_s0[65]}), .a ({signal_2712, signal_1712}), .c ({signal_2787, signal_1584}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1305 ( .s (signal_1221), .b ({ciphertext_s1[66], ciphertext_s0[66]}), .a ({signal_2715, signal_1711}), .c ({signal_2788, signal_1583}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1306 ( .s (signal_1221), .b ({ciphertext_s1[67], ciphertext_s0[67]}), .a ({signal_2718, signal_1710}), .c ({signal_2789, signal_1582}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1307 ( .s (signal_1222), .b ({ciphertext_s1[68], ciphertext_s0[68]}), .a ({signal_2343, signal_1709}), .c ({signal_2790, signal_1581}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1308 ( .s (signal_1222), .b ({ciphertext_s1[69], ciphertext_s0[69]}), .a ({signal_2346, signal_1708}), .c ({signal_2791, signal_1580}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1309 ( .s (signal_1222), .b ({ciphertext_s1[70], ciphertext_s0[70]}), .a ({signal_2349, signal_1707}), .c ({signal_2792, signal_1579}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1310 ( .s (signal_1222), .b ({ciphertext_s1[71], ciphertext_s0[71]}), .a ({signal_2352, signal_1706}), .c ({signal_2793, signal_1578}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1311 ( .s (signal_1222), .b ({ciphertext_s1[104], ciphertext_s0[104]}), .a ({signal_2688, signal_1705}), .c ({signal_2794, signal_1577}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1312 ( .s (signal_1222), .b ({ciphertext_s1[105], ciphertext_s0[105]}), .a ({signal_2721, signal_1704}), .c ({signal_2795, signal_1576}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1313 ( .s (signal_1222), .b ({ciphertext_s1[106], ciphertext_s0[106]}), .a ({signal_2373, signal_1703}), .c ({signal_2796, signal_1575}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1314 ( .s (signal_1222), .b ({ciphertext_s1[107], ciphertext_s0[107]}), .a ({signal_2406, signal_1702}), .c ({signal_2797, signal_1574}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1315 ( .s (signal_1222), .b ({ciphertext_s1[108], ciphertext_s0[108]}), .a ({signal_2433, signal_1701}), .c ({signal_2798, signal_1573}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1316 ( .s (signal_1222), .b ({ciphertext_s1[109], ciphertext_s0[109]}), .a ({signal_2436, signal_1700}), .c ({signal_2799, signal_1572}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1317 ( .s (signal_1222), .b ({ciphertext_s1[110], ciphertext_s0[110]}), .a ({signal_2439, signal_1699}), .c ({signal_2800, signal_1571}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1318 ( .s (signal_1222), .b ({ciphertext_s1[111], ciphertext_s0[111]}), .a ({signal_2442, signal_1698}), .c ({signal_2801, signal_1570}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1319 ( .s (signal_1223), .b ({ciphertext_s1[16], ciphertext_s0[16]}), .a ({signal_2550, signal_1697}), .c ({signal_2802, signal_1569}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1320 ( .s (signal_1223), .b ({ciphertext_s1[17], ciphertext_s0[17]}), .a ({signal_2553, signal_1696}), .c ({signal_2803, signal_1568}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1321 ( .s (signal_1223), .b ({ciphertext_s1[18], ciphertext_s0[18]}), .a ({signal_2559, signal_1695}), .c ({signal_2804, signal_1567}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1322 ( .s (signal_1223), .b ({ciphertext_s1[19], ciphertext_s0[19]}), .a ({signal_2562, signal_1694}), .c ({signal_2805, signal_1566}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1323 ( .s (signal_1223), .b ({ciphertext_s1[20], ciphertext_s0[20]}), .a ({signal_2565, signal_1693}), .c ({signal_2806, signal_1565}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1324 ( .s (signal_1223), .b ({ciphertext_s1[21], ciphertext_s0[21]}), .a ({signal_2568, signal_1692}), .c ({signal_2807, signal_1564}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1325 ( .s (signal_1223), .b ({ciphertext_s1[22], ciphertext_s0[22]}), .a ({signal_2571, signal_1691}), .c ({signal_2808, signal_1563}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1326 ( .s (signal_1223), .b ({ciphertext_s1[23], ciphertext_s0[23]}), .a ({signal_2574, signal_1690}), .c ({signal_2809, signal_1562}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1327 ( .s (signal_1223), .b ({ciphertext_s1[56], ciphertext_s0[56]}), .a ({signal_2682, signal_1689}), .c ({signal_2810, signal_1561}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1328 ( .s (signal_1223), .b ({ciphertext_s1[57], ciphertext_s0[57]}), .a ({signal_2685, signal_1688}), .c ({signal_2811, signal_1560}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1329 ( .s (signal_1223), .b ({ciphertext_s1[58], ciphertext_s0[58]}), .a ({signal_2691, signal_1687}), .c ({signal_2812, signal_1559}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1330 ( .s (signal_1223), .b ({ciphertext_s1[59], ciphertext_s0[59]}), .a ({signal_2694, signal_1686}), .c ({signal_2813, signal_1558}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1331 ( .s (signal_1224), .b ({ciphertext_s1[60], ciphertext_s0[60]}), .a ({signal_2697, signal_1685}), .c ({signal_2814, signal_1557}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1332 ( .s (signal_1224), .b ({ciphertext_s1[61], ciphertext_s0[61]}), .a ({signal_2700, signal_1684}), .c ({signal_2815, signal_1556}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1333 ( .s (signal_1224), .b ({ciphertext_s1[62], ciphertext_s0[62]}), .a ({signal_2703, signal_1683}), .c ({signal_2816, signal_1555}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1334 ( .s (signal_1224), .b ({ciphertext_s1[63], ciphertext_s0[63]}), .a ({signal_2706, signal_1682}), .c ({signal_2817, signal_1554}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1335 ( .s (signal_1224), .b ({ciphertext_s1[96], ciphertext_s0[96]}), .a ({signal_2340, signal_1681}), .c ({signal_2818, signal_1553}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1336 ( .s (signal_1224), .b ({ciphertext_s1[97], ciphertext_s0[97]}), .a ({signal_2457, signal_1680}), .c ({signal_2819, signal_1552}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1337 ( .s (signal_1224), .b ({ciphertext_s1[98], ciphertext_s0[98]}), .a ({signal_2490, signal_1679}), .c ({signal_2820, signal_1551}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1338 ( .s (signal_1224), .b ({ciphertext_s1[99], ciphertext_s0[99]}), .a ({signal_2523, signal_1678}), .c ({signal_2821, signal_1550}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1339 ( .s (signal_1224), .b ({ciphertext_s1[100], ciphertext_s0[100]}), .a ({signal_2556, signal_1677}), .c ({signal_2822, signal_1549}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1340 ( .s (signal_1224), .b ({ciphertext_s1[101], ciphertext_s0[101]}), .a ({signal_2589, signal_1676}), .c ({signal_2823, signal_1548}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1341 ( .s (signal_1224), .b ({ciphertext_s1[102], ciphertext_s0[102]}), .a ({signal_2622, signal_1675}), .c ({signal_2824, signal_1547}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1342 ( .s (signal_1224), .b ({ciphertext_s1[103], ciphertext_s0[103]}), .a ({signal_2655, signal_1674}), .c ({signal_2825, signal_1546}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1343 ( .s (signal_1225), .b ({ciphertext_s1[8], ciphertext_s0[8]}), .a ({signal_2526, signal_1673}), .c ({signal_2826, signal_1545}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1344 ( .s (signal_1225), .b ({ciphertext_s1[9], ciphertext_s0[9]}), .a ({signal_2529, signal_1672}), .c ({signal_2827, signal_1544}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1345 ( .s (signal_1225), .b ({ciphertext_s1[10], ciphertext_s0[10]}), .a ({signal_2532, signal_1671}), .c ({signal_2828, signal_1543}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1346 ( .s (signal_1225), .b ({ciphertext_s1[11], ciphertext_s0[11]}), .a ({signal_2535, signal_1670}), .c ({signal_2829, signal_1542}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1347 ( .s (signal_1225), .b ({ciphertext_s1[12], ciphertext_s0[12]}), .a ({signal_2538, signal_1669}), .c ({signal_2830, signal_1541}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1348 ( .s (signal_1225), .b ({ciphertext_s1[13], ciphertext_s0[13]}), .a ({signal_2541, signal_1668}), .c ({signal_2831, signal_1540}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1349 ( .s (signal_1225), .b ({ciphertext_s1[14], ciphertext_s0[14]}), .a ({signal_2544, signal_1667}), .c ({signal_2832, signal_1539}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1350 ( .s (signal_1225), .b ({ciphertext_s1[15], ciphertext_s0[15]}), .a ({signal_2547, signal_1666}), .c ({signal_2833, signal_1538}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1351 ( .s (signal_1225), .b ({ciphertext_s1[48], ciphertext_s0[48]}), .a ({signal_2658, signal_1665}), .c ({signal_2834, signal_1537}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1352 ( .s (signal_1225), .b ({ciphertext_s1[49], ciphertext_s0[49]}), .a ({signal_2661, signal_1664}), .c ({signal_2835, signal_1536}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1353 ( .s (signal_1225), .b ({ciphertext_s1[50], ciphertext_s0[50]}), .a ({signal_2664, signal_1663}), .c ({signal_2836, signal_1535}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1354 ( .s (signal_1225), .b ({ciphertext_s1[51], ciphertext_s0[51]}), .a ({signal_2667, signal_1662}), .c ({signal_2837, signal_1534}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1355 ( .s (signal_1226), .b ({ciphertext_s1[52], ciphertext_s0[52]}), .a ({signal_2670, signal_1661}), .c ({signal_2838, signal_1533}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1356 ( .s (signal_1226), .b ({ciphertext_s1[53], ciphertext_s0[53]}), .a ({signal_2673, signal_1660}), .c ({signal_2839, signal_1532}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1357 ( .s (signal_1226), .b ({ciphertext_s1[54], ciphertext_s0[54]}), .a ({signal_2676, signal_1659}), .c ({signal_2840, signal_1531}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1358 ( .s (signal_1226), .b ({ciphertext_s1[55], ciphertext_s0[55]}), .a ({signal_2679, signal_1658}), .c ({signal_2841, signal_1530}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1359 ( .s (signal_1226), .b ({ciphertext_s1[88], ciphertext_s0[88]}), .a ({signal_2409, signal_1657}), .c ({signal_2842, signal_1529}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1360 ( .s (signal_1226), .b ({ciphertext_s1[89], ciphertext_s0[89]}), .a ({signal_2412, signal_1656}), .c ({signal_2843, signal_1528}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1361 ( .s (signal_1226), .b ({ciphertext_s1[90], ciphertext_s0[90]}), .a ({signal_2415, signal_1655}), .c ({signal_2844, signal_1527}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1362 ( .s (signal_1226), .b ({ciphertext_s1[91], ciphertext_s0[91]}), .a ({signal_2418, signal_1654}), .c ({signal_2845, signal_1526}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1363 ( .s (signal_1226), .b ({ciphertext_s1[92], ciphertext_s0[92]}), .a ({signal_2421, signal_1653}), .c ({signal_2846, signal_1525}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1364 ( .s (signal_1226), .b ({ciphertext_s1[93], ciphertext_s0[93]}), .a ({signal_2424, signal_1652}), .c ({signal_2847, signal_1524}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1365 ( .s (signal_1226), .b ({ciphertext_s1[94], ciphertext_s0[94]}), .a ({signal_2427, signal_1651}), .c ({signal_2848, signal_1523}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1366 ( .s (signal_1226), .b ({ciphertext_s1[95], ciphertext_s0[95]}), .a ({signal_2430, signal_1650}), .c ({signal_2849, signal_1522}) ) ;
    INV_X1 cell_1887 ( .A (signal_1483), .ZN (signal_1490) ) ;
    INV_X1 cell_1888 ( .A (signal_393), .ZN (signal_1483) ) ;
    INV_X1 cell_1889 ( .A (signal_1483), .ZN (signal_1488) ) ;
    INV_X1 cell_1890 ( .A (signal_1483), .ZN (signal_1487) ) ;
    INV_X1 cell_1891 ( .A (signal_1483), .ZN (signal_1486) ) ;
    INV_X1 cell_1892 ( .A (signal_1483), .ZN (signal_1485) ) ;
    INV_X1 cell_1893 ( .A (signal_1483), .ZN (signal_1484) ) ;
    INV_X1 cell_1894 ( .A (signal_1483), .ZN (signal_1489) ) ;
    NOR2_X1 cell_2023 ( .A1 (reset), .A2 (signal_1491), .ZN (signal_1502) ) ;
    XNOR2_X1 cell_2024 ( .A (signal_2273), .B (signal_393), .ZN (signal_1491) ) ;
    NOR2_X1 cell_2025 ( .A1 (reset), .A2 (signal_1492), .ZN (signal_1501) ) ;
    XOR2_X1 cell_2026 ( .A (signal_2272), .B (signal_1493), .Z (signal_1492) ) ;
    NOR2_X1 cell_2027 ( .A1 (reset), .A2 (signal_1494), .ZN (signal_1498) ) ;
    XOR2_X1 cell_2028 ( .A (signal_2270), .B (signal_1495), .Z (signal_1494) ) ;
    NAND2_X1 cell_2029 ( .A1 (signal_1496), .A2 (signal_2271), .ZN (signal_1495) ) ;
    NOR2_X1 cell_2030 ( .A1 (reset), .A2 (signal_1497), .ZN (signal_1499) ) ;
    XNOR2_X1 cell_2031 ( .A (signal_2271), .B (signal_1496), .ZN (signal_1497) ) ;
    NOR2_X1 cell_2032 ( .A1 (signal_1500), .A2 (signal_1493), .ZN (signal_1496) ) ;
    NAND2_X1 cell_2033 ( .A1 (signal_393), .A2 (signal_2273), .ZN (signal_1493) ) ;
    INV_X1 cell_2036 ( .A (signal_2272), .ZN (signal_1500) ) ;
    NOR2_X1 cell_2042 ( .A1 (reset), .A2 (signal_1506), .ZN (signal_1520) ) ;
    XOR2_X1 cell_2043 ( .A (signal_2276), .B (signal_1507), .Z (signal_1506) ) ;
    NAND2_X1 cell_2044 ( .A1 (signal_1508), .A2 (1'b1), .ZN (signal_1507) ) ;
    NAND2_X1 cell_2045 ( .A1 (signal_1509), .A2 (signal_2274), .ZN (signal_1508) ) ;
    NAND2_X1 cell_2046 ( .A1 (signal_2276), .A2 (signal_2275), .ZN (signal_1509) ) ;
    NOR2_X1 cell_2047 ( .A1 (reset), .A2 (signal_1510), .ZN (signal_1519) ) ;
    MUX2_X1 cell_2048 ( .S (signal_2275), .A (signal_1511), .B (signal_1512), .Z (signal_1510) ) ;
    NOR2_X1 cell_2049 ( .A1 (reset), .A2 (signal_1513), .ZN (signal_1518) ) ;
    NOR2_X1 cell_2050 ( .A1 (signal_1514), .A2 (signal_1515), .ZN (signal_1513) ) ;
    NOR2_X1 cell_2051 ( .A1 (signal_1516), .A2 (signal_1511), .ZN (signal_1515) ) ;
    NAND2_X1 cell_2052 ( .A1 (signal_1512), .A2 (signal_1517), .ZN (signal_1511) ) ;
    AND2_X1 cell_2053 ( .A1 (signal_2276), .A2 (1'b1), .ZN (signal_1512) ) ;
    NOR2_X1 cell_2054 ( .A1 (1'b1), .A2 (signal_1517), .ZN (signal_1514) ) ;
    INV_X1 cell_2057 ( .A (signal_2275), .ZN (signal_1516) ) ;
    INV_X1 cell_2059 ( .A (signal_2274), .ZN (signal_1517) ) ;

    /* cells in depth 1 */
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_160 ( .s (signal_11952), .b ({signal_3322, signal_1649}), .a ({signal_11954, signal_11953}), .c ({signal_3437, signal_414}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_163 ( .s (signal_11952), .b ({signal_3176, signal_1648}), .a ({signal_11956, signal_11955}), .c ({signal_3263, signal_416}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_166 ( .s (signal_11952), .b ({signal_3177, signal_1647}), .a ({signal_11958, signal_11957}), .c ({signal_3265, signal_418}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_169 ( .s (signal_11952), .b ({signal_3178, signal_1646}), .a ({signal_11960, signal_11959}), .c ({signal_3267, signal_420}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_172 ( .s (signal_11952), .b ({signal_3179, signal_1645}), .a ({signal_11962, signal_11961}), .c ({signal_3269, signal_422}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_175 ( .s (signal_11952), .b ({signal_3180, signal_1644}), .a ({signal_11964, signal_11963}), .c ({signal_3271, signal_424}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_178 ( .s (signal_11952), .b ({signal_3181, signal_1643}), .a ({signal_11966, signal_11965}), .c ({signal_3273, signal_426}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_181 ( .s (signal_11952), .b ({signal_3182, signal_1642}), .a ({signal_11968, signal_11967}), .c ({signal_3275, signal_428}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_184 ( .s (signal_11952), .b ({signal_3183, signal_1641}), .a ({signal_11970, signal_11969}), .c ({signal_3277, signal_430}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_187 ( .s (signal_11952), .b ({signal_3323, signal_1640}), .a ({signal_11972, signal_11971}), .c ({signal_3439, signal_432}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_190 ( .s (signal_11952), .b ({signal_3184, signal_1639}), .a ({signal_11974, signal_11973}), .c ({signal_3279, signal_434}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_193 ( .s (signal_11952), .b ({signal_3185, signal_1638}), .a ({signal_11976, signal_11975}), .c ({signal_3281, signal_436}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_196 ( .s (signal_11952), .b ({signal_3186, signal_1637}), .a ({signal_11978, signal_11977}), .c ({signal_3283, signal_438}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_199 ( .s (signal_11952), .b ({signal_3187, signal_1636}), .a ({signal_11980, signal_11979}), .c ({signal_3285, signal_440}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_202 ( .s (signal_11952), .b ({signal_3188, signal_1635}), .a ({signal_11982, signal_11981}), .c ({signal_3287, signal_442}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_205 ( .s (signal_11952), .b ({signal_3189, signal_1634}), .a ({signal_11984, signal_11983}), .c ({signal_3289, signal_444}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_208 ( .s (signal_11952), .b ({signal_3190, signal_1633}), .a ({signal_11986, signal_11985}), .c ({signal_3291, signal_446}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_211 ( .s (signal_11952), .b ({signal_3191, signal_1632}), .a ({signal_11988, signal_11987}), .c ({signal_3293, signal_448}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_214 ( .s (signal_11952), .b ({signal_3192, signal_1631}), .a ({signal_11990, signal_11989}), .c ({signal_3295, signal_450}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_217 ( .s (signal_11952), .b ({signal_3193, signal_1630}), .a ({signal_11992, signal_11991}), .c ({signal_3297, signal_452}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_220 ( .s (signal_11952), .b ({signal_3194, signal_1629}), .a ({signal_11994, signal_11993}), .c ({signal_3299, signal_454}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_223 ( .s (signal_11952), .b ({signal_3195, signal_1628}), .a ({signal_11996, signal_11995}), .c ({signal_3301, signal_456}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_226 ( .s (signal_11952), .b ({signal_3196, signal_1627}), .a ({signal_11998, signal_11997}), .c ({signal_3303, signal_458}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_229 ( .s (signal_11952), .b ({signal_3197, signal_1626}), .a ({signal_12000, signal_11999}), .c ({signal_3305, signal_460}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_232 ( .s (signal_11952), .b ({signal_3198, signal_1625}), .a ({signal_12002, signal_12001}), .c ({signal_3307, signal_462}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_235 ( .s (signal_11952), .b ({signal_3199, signal_1624}), .a ({signal_12004, signal_12003}), .c ({signal_3309, signal_464}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_238 ( .s (signal_11952), .b ({signal_3200, signal_1623}), .a ({signal_12006, signal_12005}), .c ({signal_3311, signal_466}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_241 ( .s (signal_11952), .b ({signal_3201, signal_1622}), .a ({signal_12008, signal_12007}), .c ({signal_3313, signal_468}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_244 ( .s (signal_11952), .b ({signal_3202, signal_1621}), .a ({signal_12010, signal_12009}), .c ({signal_3315, signal_470}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_247 ( .s (signal_11952), .b ({signal_3203, signal_1620}), .a ({signal_12012, signal_12011}), .c ({signal_3317, signal_472}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_250 ( .s (signal_11952), .b ({signal_3204, signal_1619}), .a ({signal_12014, signal_12013}), .c ({signal_3319, signal_474}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_253 ( .s (signal_11952), .b ({signal_3205, signal_1618}), .a ({signal_12016, signal_12015}), .c ({signal_3321, signal_476}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_1089 ( .a ({signal_3046, signal_1153}), .b ({signal_3100, signal_2328}), .c ({signal_3110, signal_1868}) ) ;
    xnor_GHPC #(.low_latency(1), .pipeline(1)) cell_1181 ( .a ({signal_3047, signal_1216}), .b ({signal_3093, signal_2321}), .c ({signal_3111, signal_1877}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1200 ( .s (signal_12017), .b ({signal_3111, signal_1877}), .a ({signal_3050, signal_1845}), .c ({signal_3174, signal_1909}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1201 ( .s (signal_12018), .b ({signal_3080, signal_1876}), .a ({signal_3084, signal_2303}), .c ({signal_3112, signal_1908}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1202 ( .s (signal_12018), .b ({signal_3079, signal_1875}), .a ({signal_3049, signal_1843}), .c ({signal_3113, signal_1907}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1203 ( .s (signal_12018), .b ({signal_3078, signal_1874}), .a ({signal_3048, signal_1842}), .c ({signal_3114, signal_1906}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1204 ( .s (signal_12018), .b ({signal_3077, signal_1873}), .a ({signal_3083, signal_2300}), .c ({signal_3115, signal_1905}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1205 ( .s (signal_12018), .b ({signal_3076, signal_1872}), .a ({signal_3082, signal_2299}), .c ({signal_3116, signal_1904}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1206 ( .s (signal_12018), .b ({signal_3075, signal_1871}), .a ({signal_3081, signal_2298}), .c ({signal_3117, signal_1903}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1207 ( .s (signal_12019), .b ({signal_3074, signal_1870}), .a ({signal_3085, signal_2305}), .c ({signal_3118, signal_1902}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1208 ( .s (signal_12017), .b ({signal_3073, signal_1869}), .a ({signal_3093, signal_2321}), .c ({signal_3119, signal_1901}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1209 ( .s (signal_12017), .b ({signal_3110, signal_1868}), .a ({signal_3092, signal_2320}), .c ({signal_3175, signal_1900}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1210 ( .s (signal_12017), .b ({signal_3072, signal_1867}), .a ({signal_3091, signal_2319}), .c ({signal_3120, signal_1899}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1211 ( .s (signal_12017), .b ({signal_3071, signal_1866}), .a ({signal_3090, signal_2318}), .c ({signal_3121, signal_1898}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1212 ( .s (signal_12017), .b ({signal_3070, signal_1865}), .a ({signal_3089, signal_2317}), .c ({signal_3122, signal_1897}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1213 ( .s (signal_12017), .b ({signal_3069, signal_1864}), .a ({signal_3088, signal_2316}), .c ({signal_3123, signal_1896}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1214 ( .s (signal_12017), .b ({signal_3068, signal_1863}), .a ({signal_3087, signal_2315}), .c ({signal_3124, signal_1895}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1215 ( .s (signal_12017), .b ({signal_3067, signal_1862}), .a ({signal_3086, signal_2314}), .c ({signal_3125, signal_1894}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1216 ( .s (signal_12017), .b ({signal_3066, signal_1861}), .a ({signal_3101, signal_2329}), .c ({signal_3126, signal_1893}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1217 ( .s (signal_12017), .b ({signal_3065, signal_1860}), .a ({signal_3100, signal_2328}), .c ({signal_3127, signal_1892}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1218 ( .s (signal_12017), .b ({signal_3064, signal_1859}), .a ({signal_3099, signal_2327}), .c ({signal_3128, signal_1891}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1219 ( .s (signal_12017), .b ({signal_3063, signal_1858}), .a ({signal_3098, signal_2326}), .c ({signal_3129, signal_1890}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1220 ( .s (signal_12019), .b ({signal_3062, signal_1857}), .a ({signal_3097, signal_2325}), .c ({signal_3130, signal_1889}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1221 ( .s (signal_12019), .b ({signal_3061, signal_1856}), .a ({signal_3096, signal_2324}), .c ({signal_3131, signal_1888}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1222 ( .s (signal_12019), .b ({signal_3060, signal_1855}), .a ({signal_3095, signal_2323}), .c ({signal_3132, signal_1887}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1223 ( .s (signal_12019), .b ({signal_3059, signal_1854}), .a ({signal_3094, signal_2322}), .c ({signal_3133, signal_1886}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1224 ( .s (signal_12019), .b ({signal_3058, signal_1853}), .a ({signal_3109, signal_2337}), .c ({signal_3134, signal_1885}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1225 ( .s (signal_12019), .b ({signal_3057, signal_1852}), .a ({signal_3108, signal_2336}), .c ({signal_3135, signal_1884}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1226 ( .s (signal_12019), .b ({signal_3056, signal_1851}), .a ({signal_3107, signal_2335}), .c ({signal_3136, signal_1883}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1227 ( .s (signal_12019), .b ({signal_3055, signal_1850}), .a ({signal_3106, signal_2334}), .c ({signal_3137, signal_1882}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1228 ( .s (signal_12019), .b ({signal_3054, signal_1849}), .a ({signal_3105, signal_2333}), .c ({signal_3138, signal_1881}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1229 ( .s (signal_12019), .b ({signal_3053, signal_1848}), .a ({signal_3104, signal_2332}), .c ({signal_3139, signal_1880}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1230 ( .s (signal_12019), .b ({signal_3052, signal_1847}), .a ({signal_3103, signal_2331}), .c ({signal_3140, signal_1879}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1231 ( .s (signal_12019), .b ({signal_3051, signal_1846}), .a ({signal_3102, signal_2330}), .c ({signal_3141, signal_1878}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1239 ( .s (signal_12020), .b ({signal_3174, signal_1909}), .a ({signal_12022, signal_12021}), .c ({signal_3322, signal_1649}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1240 ( .s (signal_12023), .b ({signal_3112, signal_1908}), .a ({signal_12025, signal_12024}), .c ({signal_3176, signal_1648}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1241 ( .s (signal_12026), .b ({signal_3113, signal_1907}), .a ({signal_12028, signal_12027}), .c ({signal_3177, signal_1647}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1242 ( .s (signal_12029), .b ({signal_3114, signal_1906}), .a ({signal_12031, signal_12030}), .c ({signal_3178, signal_1646}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1243 ( .s (signal_12032), .b ({signal_3115, signal_1905}), .a ({signal_12034, signal_12033}), .c ({signal_3179, signal_1645}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1244 ( .s (signal_12035), .b ({signal_3116, signal_1904}), .a ({signal_12037, signal_12036}), .c ({signal_3180, signal_1644}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1245 ( .s (signal_12038), .b ({signal_3117, signal_1903}), .a ({signal_12040, signal_12039}), .c ({signal_3181, signal_1643}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1246 ( .s (signal_12023), .b ({signal_3118, signal_1902}), .a ({signal_12042, signal_12041}), .c ({signal_3182, signal_1642}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1247 ( .s (signal_12032), .b ({signal_3119, signal_1901}), .a ({signal_12044, signal_12043}), .c ({signal_3183, signal_1641}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1248 ( .s (signal_12023), .b ({signal_3175, signal_1900}), .a ({signal_12046, signal_12045}), .c ({signal_3323, signal_1640}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1249 ( .s (signal_12020), .b ({signal_3120, signal_1899}), .a ({signal_12048, signal_12047}), .c ({signal_3184, signal_1639}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1250 ( .s (signal_12020), .b ({signal_3121, signal_1898}), .a ({signal_12050, signal_12049}), .c ({signal_3185, signal_1638}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1251 ( .s (signal_12020), .b ({signal_3122, signal_1897}), .a ({signal_12052, signal_12051}), .c ({signal_3186, signal_1637}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1252 ( .s (signal_12020), .b ({signal_3123, signal_1896}), .a ({signal_12054, signal_12053}), .c ({signal_3187, signal_1636}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1253 ( .s (signal_12020), .b ({signal_3124, signal_1895}), .a ({signal_12056, signal_12055}), .c ({signal_3188, signal_1635}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1254 ( .s (signal_12020), .b ({signal_3125, signal_1894}), .a ({signal_12058, signal_12057}), .c ({signal_3189, signal_1634}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1255 ( .s (signal_12020), .b ({signal_3126, signal_1893}), .a ({signal_12060, signal_12059}), .c ({signal_3190, signal_1633}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1256 ( .s (signal_12020), .b ({signal_3127, signal_1892}), .a ({signal_12062, signal_12061}), .c ({signal_3191, signal_1632}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1257 ( .s (signal_12020), .b ({signal_3128, signal_1891}), .a ({signal_12064, signal_12063}), .c ({signal_3192, signal_1631}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1258 ( .s (signal_12020), .b ({signal_3129, signal_1890}), .a ({signal_12066, signal_12065}), .c ({signal_3193, signal_1630}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1259 ( .s (signal_12026), .b ({signal_3130, signal_1889}), .a ({signal_12068, signal_12067}), .c ({signal_3194, signal_1629}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1260 ( .s (signal_12029), .b ({signal_3131, signal_1888}), .a ({signal_12070, signal_12069}), .c ({signal_3195, signal_1628}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1261 ( .s (signal_12032), .b ({signal_3132, signal_1887}), .a ({signal_12072, signal_12071}), .c ({signal_3196, signal_1627}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1262 ( .s (signal_12035), .b ({signal_3133, signal_1886}), .a ({signal_12074, signal_12073}), .c ({signal_3197, signal_1626}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1263 ( .s (signal_12038), .b ({signal_3134, signal_1885}), .a ({signal_12076, signal_12075}), .c ({signal_3198, signal_1625}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1264 ( .s (signal_12032), .b ({signal_3135, signal_1884}), .a ({signal_12078, signal_12077}), .c ({signal_3199, signal_1624}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1265 ( .s (signal_12035), .b ({signal_3136, signal_1883}), .a ({signal_12080, signal_12079}), .c ({signal_3200, signal_1623}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1266 ( .s (signal_12020), .b ({signal_3137, signal_1882}), .a ({signal_12082, signal_12081}), .c ({signal_3201, signal_1622}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1267 ( .s (signal_12020), .b ({signal_3138, signal_1881}), .a ({signal_12084, signal_12083}), .c ({signal_3202, signal_1621}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1268 ( .s (signal_12023), .b ({signal_3139, signal_1880}), .a ({signal_12086, signal_12085}), .c ({signal_3203, signal_1620}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1269 ( .s (signal_12026), .b ({signal_3140, signal_1879}), .a ({signal_12088, signal_12087}), .c ({signal_3204, signal_1619}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1270 ( .s (signal_12029), .b ({signal_3141, signal_1878}), .a ({signal_12090, signal_12089}), .c ({signal_3205, signal_1618}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1369 ( .s (signal_11952), .b ({signal_3640, signal_2037}), .a ({signal_12092, signal_12091}), .c ({signal_3673, signal_1227}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1372 ( .s (signal_11952), .b ({signal_3641, signal_2036}), .a ({signal_12094, signal_12093}), .c ({signal_3675, signal_1229}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1375 ( .s (signal_11952), .b ({signal_3642, signal_2035}), .a ({signal_12096, signal_12095}), .c ({signal_3677, signal_1231}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1378 ( .s (signal_11952), .b ({signal_3643, signal_2034}), .a ({signal_12098, signal_12097}), .c ({signal_3679, signal_1233}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1381 ( .s (signal_11952), .b ({signal_3644, signal_2033}), .a ({signal_12100, signal_12099}), .c ({signal_3681, signal_1235}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1384 ( .s (signal_11952), .b ({signal_3645, signal_2032}), .a ({signal_12102, signal_12101}), .c ({signal_3683, signal_1237}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1387 ( .s (signal_11952), .b ({signal_3646, signal_2031}), .a ({signal_12104, signal_12103}), .c ({signal_3685, signal_1239}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1390 ( .s (signal_11952), .b ({signal_3647, signal_2030}), .a ({signal_12106, signal_12105}), .c ({signal_3687, signal_1241}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1393 ( .s (signal_11952), .b ({signal_3648, signal_2029}), .a ({signal_12108, signal_12107}), .c ({signal_3689, signal_1243}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1396 ( .s (signal_11952), .b ({signal_3649, signal_2028}), .a ({signal_12110, signal_12109}), .c ({signal_3691, signal_1245}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1399 ( .s (signal_11952), .b ({signal_3650, signal_2027}), .a ({signal_12112, signal_12111}), .c ({signal_3693, signal_1247}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1402 ( .s (signal_11952), .b ({signal_3651, signal_2026}), .a ({signal_12114, signal_12113}), .c ({signal_3695, signal_1249}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1405 ( .s (signal_11952), .b ({signal_3652, signal_2025}), .a ({signal_12116, signal_12115}), .c ({signal_3697, signal_1251}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1408 ( .s (signal_11952), .b ({signal_3653, signal_2024}), .a ({signal_12118, signal_12117}), .c ({signal_3699, signal_1253}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1411 ( .s (signal_11952), .b ({signal_3654, signal_2023}), .a ({signal_12120, signal_12119}), .c ({signal_3701, signal_1255}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1414 ( .s (signal_11952), .b ({signal_3655, signal_2022}), .a ({signal_12122, signal_12121}), .c ({signal_3703, signal_1257}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1417 ( .s (signal_11952), .b ({signal_3656, signal_2021}), .a ({signal_12124, signal_12123}), .c ({signal_3705, signal_1259}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1420 ( .s (signal_11952), .b ({signal_3657, signal_2020}), .a ({signal_12126, signal_12125}), .c ({signal_3707, signal_1261}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1423 ( .s (signal_11952), .b ({signal_3658, signal_2019}), .a ({signal_12128, signal_12127}), .c ({signal_3709, signal_1263}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1426 ( .s (signal_11952), .b ({signal_3659, signal_2018}), .a ({signal_12130, signal_12129}), .c ({signal_3711, signal_1265}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1429 ( .s (signal_11952), .b ({signal_3660, signal_2017}), .a ({signal_12132, signal_12131}), .c ({signal_3713, signal_1267}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1432 ( .s (signal_11952), .b ({signal_3661, signal_2016}), .a ({signal_12134, signal_12133}), .c ({signal_3715, signal_1269}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1435 ( .s (signal_11952), .b ({signal_3662, signal_2015}), .a ({signal_12136, signal_12135}), .c ({signal_3717, signal_1271}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1438 ( .s (signal_11952), .b ({signal_3663, signal_2014}), .a ({signal_12138, signal_12137}), .c ({signal_3719, signal_1273}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1441 ( .s (signal_11952), .b ({signal_3736, signal_2013}), .a ({signal_12140, signal_12139}), .c ({signal_3745, signal_1275}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1444 ( .s (signal_11952), .b ({signal_3737, signal_2012}), .a ({signal_12142, signal_12141}), .c ({signal_3747, signal_1277}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1447 ( .s (signal_11952), .b ({signal_3738, signal_2011}), .a ({signal_12144, signal_12143}), .c ({signal_3749, signal_1279}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1450 ( .s (signal_11952), .b ({signal_3739, signal_2010}), .a ({signal_12146, signal_12145}), .c ({signal_3751, signal_1281}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1453 ( .s (signal_11952), .b ({signal_3740, signal_2009}), .a ({signal_12148, signal_12147}), .c ({signal_3753, signal_1283}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1456 ( .s (signal_11952), .b ({signal_3741, signal_2008}), .a ({signal_12150, signal_12149}), .c ({signal_3755, signal_1285}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1459 ( .s (signal_11952), .b ({signal_3742, signal_2007}), .a ({signal_12152, signal_12151}), .c ({signal_3757, signal_1287}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1462 ( .s (signal_11952), .b ({signal_3743, signal_2006}), .a ({signal_12154, signal_12153}), .c ({signal_3759, signal_1289}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1465 ( .s (signal_11952), .b ({signal_3536, signal_2005}), .a ({signal_12156, signal_12155}), .c ({signal_3569, signal_1291}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1468 ( .s (signal_11952), .b ({signal_3537, signal_2004}), .a ({signal_12158, signal_12157}), .c ({signal_3571, signal_1293}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1471 ( .s (signal_11952), .b ({signal_3538, signal_2003}), .a ({signal_12160, signal_12159}), .c ({signal_3573, signal_1295}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1474 ( .s (signal_11952), .b ({signal_3539, signal_2002}), .a ({signal_12162, signal_12161}), .c ({signal_3575, signal_1297}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1477 ( .s (signal_11952), .b ({signal_3540, signal_2001}), .a ({signal_12164, signal_12163}), .c ({signal_3577, signal_1299}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1480 ( .s (signal_11952), .b ({signal_3541, signal_2000}), .a ({signal_12166, signal_12165}), .c ({signal_3579, signal_1301}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1483 ( .s (signal_11952), .b ({signal_3542, signal_1999}), .a ({signal_12168, signal_12167}), .c ({signal_3581, signal_1303}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1486 ( .s (signal_11952), .b ({signal_3543, signal_1998}), .a ({signal_12170, signal_12169}), .c ({signal_3583, signal_1305}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1489 ( .s (signal_11952), .b ({signal_3544, signal_1997}), .a ({signal_12172, signal_12171}), .c ({signal_3585, signal_1307}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1492 ( .s (signal_11952), .b ({signal_3545, signal_1996}), .a ({signal_12174, signal_12173}), .c ({signal_3587, signal_1309}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1495 ( .s (signal_11952), .b ({signal_3546, signal_1995}), .a ({signal_12176, signal_12175}), .c ({signal_3589, signal_1311}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1498 ( .s (signal_11952), .b ({signal_3547, signal_1994}), .a ({signal_12178, signal_12177}), .c ({signal_3591, signal_1313}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1501 ( .s (signal_11952), .b ({signal_3548, signal_1993}), .a ({signal_12180, signal_12179}), .c ({signal_3593, signal_1315}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1504 ( .s (signal_11952), .b ({signal_3549, signal_1992}), .a ({signal_12182, signal_12181}), .c ({signal_3595, signal_1317}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1507 ( .s (signal_11952), .b ({signal_3550, signal_1991}), .a ({signal_12184, signal_12183}), .c ({signal_3597, signal_1319}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1510 ( .s (signal_11952), .b ({signal_3551, signal_1990}), .a ({signal_12186, signal_12185}), .c ({signal_3599, signal_1321}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1513 ( .s (signal_11952), .b ({signal_3552, signal_1989}), .a ({signal_12188, signal_12187}), .c ({signal_3601, signal_1323}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1516 ( .s (signal_11952), .b ({signal_3553, signal_1988}), .a ({signal_12190, signal_12189}), .c ({signal_3603, signal_1325}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1519 ( .s (signal_11952), .b ({signal_3554, signal_1987}), .a ({signal_12192, signal_12191}), .c ({signal_3605, signal_1327}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1522 ( .s (signal_11952), .b ({signal_3555, signal_1986}), .a ({signal_12194, signal_12193}), .c ({signal_3607, signal_1329}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1525 ( .s (signal_11952), .b ({signal_3556, signal_1985}), .a ({signal_12196, signal_12195}), .c ({signal_3609, signal_1331}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1528 ( .s (signal_11952), .b ({signal_3557, signal_1984}), .a ({signal_12198, signal_12197}), .c ({signal_3611, signal_1333}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1531 ( .s (signal_11952), .b ({signal_3558, signal_1983}), .a ({signal_12200, signal_12199}), .c ({signal_3613, signal_1335}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1534 ( .s (signal_11952), .b ({signal_3559, signal_1982}), .a ({signal_12202, signal_12201}), .c ({signal_3615, signal_1337}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1537 ( .s (signal_11952), .b ({signal_3664, signal_1981}), .a ({signal_12204, signal_12203}), .c ({signal_3721, signal_1339}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1540 ( .s (signal_11952), .b ({signal_3665, signal_1980}), .a ({signal_12206, signal_12205}), .c ({signal_3723, signal_1341}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1543 ( .s (signal_11952), .b ({signal_3666, signal_1979}), .a ({signal_12208, signal_12207}), .c ({signal_3725, signal_1343}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1546 ( .s (signal_11952), .b ({signal_3667, signal_1978}), .a ({signal_12210, signal_12209}), .c ({signal_3727, signal_1345}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1549 ( .s (signal_11952), .b ({signal_3668, signal_1977}), .a ({signal_12212, signal_12211}), .c ({signal_3729, signal_1347}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1552 ( .s (signal_11952), .b ({signal_3669, signal_1976}), .a ({signal_12214, signal_12213}), .c ({signal_3731, signal_1349}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1555 ( .s (signal_11952), .b ({signal_3670, signal_1975}), .a ({signal_12216, signal_12215}), .c ({signal_3733, signal_1351}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1558 ( .s (signal_11952), .b ({signal_3671, signal_1974}), .a ({signal_12218, signal_12217}), .c ({signal_3735, signal_1353}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1561 ( .s (signal_11952), .b ({signal_3404, signal_1973}), .a ({signal_12220, signal_12219}), .c ({signal_3441, signal_1355}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1564 ( .s (signal_11952), .b ({signal_3405, signal_1972}), .a ({signal_12222, signal_12221}), .c ({signal_3443, signal_1357}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1567 ( .s (signal_11952), .b ({signal_3406, signal_1971}), .a ({signal_12224, signal_12223}), .c ({signal_3445, signal_1359}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1570 ( .s (signal_11952), .b ({signal_3407, signal_1970}), .a ({signal_12226, signal_12225}), .c ({signal_3447, signal_1361}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1573 ( .s (signal_11952), .b ({signal_3408, signal_1969}), .a ({signal_12228, signal_12227}), .c ({signal_3449, signal_1363}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1576 ( .s (signal_11952), .b ({signal_3409, signal_1968}), .a ({signal_12230, signal_12229}), .c ({signal_3451, signal_1365}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1579 ( .s (signal_11952), .b ({signal_3410, signal_1967}), .a ({signal_12232, signal_12231}), .c ({signal_3453, signal_1367}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1582 ( .s (signal_11952), .b ({signal_3411, signal_1966}), .a ({signal_12234, signal_12233}), .c ({signal_3455, signal_1369}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1585 ( .s (signal_11952), .b ({signal_3412, signal_1965}), .a ({signal_12236, signal_12235}), .c ({signal_3457, signal_1371}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1588 ( .s (signal_11952), .b ({signal_3413, signal_1964}), .a ({signal_12238, signal_12237}), .c ({signal_3459, signal_1373}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1591 ( .s (signal_11952), .b ({signal_3414, signal_1963}), .a ({signal_12240, signal_12239}), .c ({signal_3461, signal_1375}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1594 ( .s (signal_11952), .b ({signal_3415, signal_1962}), .a ({signal_12242, signal_12241}), .c ({signal_3463, signal_1377}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1597 ( .s (signal_11952), .b ({signal_3416, signal_1961}), .a ({signal_12244, signal_12243}), .c ({signal_3465, signal_1379}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1600 ( .s (signal_11952), .b ({signal_3417, signal_1960}), .a ({signal_12246, signal_12245}), .c ({signal_3467, signal_1381}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1603 ( .s (signal_11952), .b ({signal_3418, signal_1959}), .a ({signal_12248, signal_12247}), .c ({signal_3469, signal_1383}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1606 ( .s (signal_11952), .b ({signal_3419, signal_1958}), .a ({signal_12250, signal_12249}), .c ({signal_3471, signal_1385}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1609 ( .s (signal_11952), .b ({signal_3420, signal_1957}), .a ({signal_12252, signal_12251}), .c ({signal_3473, signal_1387}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1612 ( .s (signal_11952), .b ({signal_3421, signal_1956}), .a ({signal_12254, signal_12253}), .c ({signal_3475, signal_1389}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1615 ( .s (signal_11952), .b ({signal_3422, signal_1955}), .a ({signal_12256, signal_12255}), .c ({signal_3477, signal_1391}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1618 ( .s (signal_11952), .b ({signal_3423, signal_1954}), .a ({signal_12258, signal_12257}), .c ({signal_3479, signal_1393}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1621 ( .s (signal_11952), .b ({signal_3424, signal_1953}), .a ({signal_12260, signal_12259}), .c ({signal_3481, signal_1395}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1624 ( .s (signal_11952), .b ({signal_3425, signal_1952}), .a ({signal_12262, signal_12261}), .c ({signal_3483, signal_1397}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1627 ( .s (signal_11952), .b ({signal_3426, signal_1951}), .a ({signal_12264, signal_12263}), .c ({signal_3485, signal_1399}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1630 ( .s (signal_11952), .b ({signal_3427, signal_1950}), .a ({signal_12266, signal_12265}), .c ({signal_3487, signal_1401}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1633 ( .s (signal_11952), .b ({signal_3560, signal_1949}), .a ({signal_12268, signal_12267}), .c ({signal_3617, signal_1403}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1636 ( .s (signal_11952), .b ({signal_3561, signal_1948}), .a ({signal_12270, signal_12269}), .c ({signal_3619, signal_1405}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1639 ( .s (signal_11952), .b ({signal_3562, signal_1947}), .a ({signal_12272, signal_12271}), .c ({signal_3621, signal_1407}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1642 ( .s (signal_11952), .b ({signal_3563, signal_1946}), .a ({signal_12274, signal_12273}), .c ({signal_3623, signal_1409}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1645 ( .s (signal_11952), .b ({signal_3564, signal_1945}), .a ({signal_12276, signal_12275}), .c ({signal_3625, signal_1411}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1648 ( .s (signal_11952), .b ({signal_3565, signal_1944}), .a ({signal_12278, signal_12277}), .c ({signal_3627, signal_1413}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1651 ( .s (signal_11952), .b ({signal_3566, signal_1943}), .a ({signal_12280, signal_12279}), .c ({signal_3629, signal_1415}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1654 ( .s (signal_11952), .b ({signal_3567, signal_1942}), .a ({signal_12282, signal_12281}), .c ({signal_3631, signal_1417}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1657 ( .s (signal_11952), .b ({signal_3238, signal_1941}), .a ({signal_12284, signal_12283}), .c ({signal_3325, signal_1419}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1660 ( .s (signal_11952), .b ({signal_3239, signal_1940}), .a ({signal_12286, signal_12285}), .c ({signal_3327, signal_1421}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1663 ( .s (signal_11952), .b ({signal_3240, signal_1939}), .a ({signal_12288, signal_12287}), .c ({signal_3329, signal_1423}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1666 ( .s (signal_11952), .b ({signal_3241, signal_1938}), .a ({signal_12290, signal_12289}), .c ({signal_3331, signal_1425}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1669 ( .s (signal_11952), .b ({signal_3242, signal_1937}), .a ({signal_12292, signal_12291}), .c ({signal_3333, signal_1427}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1672 ( .s (signal_11952), .b ({signal_3243, signal_1936}), .a ({signal_12294, signal_12293}), .c ({signal_3335, signal_1429}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1675 ( .s (signal_11952), .b ({signal_3244, signal_1935}), .a ({signal_12296, signal_12295}), .c ({signal_3337, signal_1431}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1678 ( .s (signal_11952), .b ({signal_3245, signal_1934}), .a ({signal_12298, signal_12297}), .c ({signal_3339, signal_1433}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1681 ( .s (signal_11952), .b ({signal_3246, signal_1933}), .a ({signal_12300, signal_12299}), .c ({signal_3341, signal_1435}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1684 ( .s (signal_11952), .b ({signal_3247, signal_1932}), .a ({signal_12302, signal_12301}), .c ({signal_3343, signal_1437}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1687 ( .s (signal_11952), .b ({signal_3248, signal_1931}), .a ({signal_12304, signal_12303}), .c ({signal_3345, signal_1439}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1690 ( .s (signal_11952), .b ({signal_3249, signal_1930}), .a ({signal_12306, signal_12305}), .c ({signal_3347, signal_1441}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1693 ( .s (signal_11952), .b ({signal_3250, signal_1929}), .a ({signal_12308, signal_12307}), .c ({signal_3349, signal_1443}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1696 ( .s (signal_11952), .b ({signal_3251, signal_1928}), .a ({signal_12310, signal_12309}), .c ({signal_3351, signal_1445}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1699 ( .s (signal_11952), .b ({signal_3252, signal_1927}), .a ({signal_12312, signal_12311}), .c ({signal_3353, signal_1447}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1702 ( .s (signal_11952), .b ({signal_3253, signal_1926}), .a ({signal_12314, signal_12313}), .c ({signal_3355, signal_1449}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1705 ( .s (signal_11952), .b ({signal_3254, signal_1925}), .a ({signal_12316, signal_12315}), .c ({signal_3357, signal_1451}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1708 ( .s (signal_11952), .b ({signal_3255, signal_1924}), .a ({signal_12318, signal_12317}), .c ({signal_3359, signal_1453}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1711 ( .s (signal_11952), .b ({signal_3256, signal_1923}), .a ({signal_12320, signal_12319}), .c ({signal_3361, signal_1455}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1714 ( .s (signal_11952), .b ({signal_3257, signal_1922}), .a ({signal_12322, signal_12321}), .c ({signal_3363, signal_1457}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1717 ( .s (signal_11952), .b ({signal_3258, signal_1921}), .a ({signal_12324, signal_12323}), .c ({signal_3365, signal_1459}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1720 ( .s (signal_11952), .b ({signal_3259, signal_1920}), .a ({signal_12326, signal_12325}), .c ({signal_3367, signal_1461}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1723 ( .s (signal_11952), .b ({signal_3260, signal_1919}), .a ({signal_12328, signal_12327}), .c ({signal_3369, signal_1463}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1726 ( .s (signal_11952), .b ({signal_3261, signal_1918}), .a ({signal_12330, signal_12329}), .c ({signal_3371, signal_1465}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1729 ( .s (signal_11952), .b ({signal_3428, signal_1917}), .a ({signal_12332, signal_12331}), .c ({signal_3489, signal_1467}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1732 ( .s (signal_11952), .b ({signal_3429, signal_1916}), .a ({signal_12334, signal_12333}), .c ({signal_3491, signal_1469}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1735 ( .s (signal_11952), .b ({signal_3430, signal_1915}), .a ({signal_12336, signal_12335}), .c ({signal_3493, signal_1471}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1738 ( .s (signal_11952), .b ({signal_3431, signal_1914}), .a ({signal_12338, signal_12337}), .c ({signal_3495, signal_1473}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1741 ( .s (signal_11952), .b ({signal_3432, signal_1913}), .a ({signal_12340, signal_12339}), .c ({signal_3497, signal_1475}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1744 ( .s (signal_11952), .b ({signal_3433, signal_1912}), .a ({signal_12342, signal_12341}), .c ({signal_3499, signal_1477}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1747 ( .s (signal_11952), .b ({signal_3434, signal_1911}), .a ({signal_12344, signal_12343}), .c ({signal_3501, signal_1479}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1750 ( .s (signal_11952), .b ({signal_3435, signal_1910}), .a ({signal_12346, signal_12345}), .c ({signal_3503, signal_1481}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1751 ( .a ({signal_12348, signal_12347}), .b ({signal_3372, signal_2228}), .c ({signal_3504, signal_2260}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1752 ( .a ({signal_12350, signal_12349}), .b ({signal_3373, signal_2229}), .c ({signal_3505, signal_2261}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1753 ( .a ({signal_12352, signal_12351}), .b ({signal_3374, signal_2230}), .c ({signal_3506, signal_2262}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1754 ( .a ({signal_12354, signal_12353}), .b ({signal_3375, signal_2231}), .c ({signal_3507, signal_2263}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1755 ( .a ({signal_12356, signal_12355}), .b ({signal_3376, signal_2232}), .c ({signal_3508, signal_2264}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1756 ( .a ({signal_12358, signal_12357}), .b ({signal_3377, signal_2233}), .c ({signal_3509, signal_2265}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1757 ( .a ({signal_12360, signal_12359}), .b ({signal_3206, signal_2196}), .c ({signal_3372, signal_2228}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1758 ( .a ({signal_12362, signal_12361}), .b ({signal_3159, signal_2164}), .c ({signal_3206, signal_2196}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1759 ( .a ({signal_12364, signal_12363}), .b ({signal_3207, signal_2197}), .c ({signal_3373, signal_2229}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1760 ( .a ({signal_12366, signal_12365}), .b ({signal_3160, signal_2165}), .c ({signal_3207, signal_2197}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1761 ( .a ({signal_12368, signal_12367}), .b ({signal_3378, signal_2234}), .c ({signal_3510, signal_2266}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1762 ( .a ({signal_12370, signal_12369}), .b ({signal_3208, signal_2198}), .c ({signal_3374, signal_2230}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1763 ( .a ({signal_12372, signal_12371}), .b ({signal_3161, signal_2166}), .c ({signal_3208, signal_2198}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1764 ( .a ({signal_12374, signal_12373}), .b ({signal_3209, signal_2199}), .c ({signal_3375, signal_2231}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1765 ( .a ({signal_12376, signal_12375}), .b ({signal_3162, signal_2167}), .c ({signal_3209, signal_2199}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1766 ( .a ({signal_12378, signal_12377}), .b ({signal_3210, signal_2200}), .c ({signal_3376, signal_2232}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1767 ( .a ({signal_12380, signal_12379}), .b ({signal_3163, signal_2168}), .c ({signal_3210, signal_2200}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1768 ( .a ({signal_12382, signal_12381}), .b ({signal_3211, signal_2201}), .c ({signal_3377, signal_2233}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1769 ( .a ({signal_12384, signal_12383}), .b ({signal_3164, signal_2169}), .c ({signal_3211, signal_2201}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1770 ( .a ({signal_12386, signal_12385}), .b ({signal_3212, signal_2202}), .c ({signal_3378, signal_2234}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1771 ( .a ({signal_12388, signal_12387}), .b ({signal_3142, signal_2170}), .c ({signal_3212, signal_2202}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1772 ( .a ({signal_12390, signal_12389}), .b ({signal_3106, signal_2334}), .c ({signal_3142, signal_2170}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1773 ( .a ({signal_12392, signal_12391}), .b ({signal_3511, signal_2206}), .c ({signal_3632, signal_2238}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1774 ( .a ({signal_12394, signal_12393}), .b ({signal_3379, signal_2174}), .c ({signal_3511, signal_2206}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1775 ( .a ({signal_12396, signal_12395}), .b ({signal_3227, signal_2142}), .c ({signal_3379, signal_2174}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1776 ( .a ({signal_12398, signal_12397}), .b ({signal_3512, signal_2207}), .c ({signal_3633, signal_2239}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1777 ( .a ({signal_12400, signal_12399}), .b ({signal_3380, signal_2175}), .c ({signal_3512, signal_2207}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1778 ( .a ({signal_12402, signal_12401}), .b ({signal_3228, signal_2143}), .c ({signal_3380, signal_2175}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1779 ( .a ({signal_12404, signal_12403}), .b ({signal_3381, signal_2235}), .c ({signal_3513, signal_2267}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1780 ( .a ({signal_12406, signal_12405}), .b ({signal_3213, signal_2203}), .c ({signal_3381, signal_2235}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1781 ( .a ({signal_12408, signal_12407}), .b ({signal_3143, signal_2171}), .c ({signal_3213, signal_2203}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1782 ( .a ({signal_12410, signal_12409}), .b ({signal_3107, signal_2335}), .c ({signal_3143, signal_2171}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1783 ( .a ({signal_12412, signal_12411}), .b ({signal_3514, signal_2208}), .c ({signal_3634, signal_2240}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1784 ( .a ({signal_12414, signal_12413}), .b ({signal_3382, signal_2176}), .c ({signal_3514, signal_2208}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1785 ( .a ({signal_12416, signal_12415}), .b ({signal_3229, signal_2144}), .c ({signal_3382, signal_2176}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1786 ( .a ({signal_12418, signal_12417}), .b ({signal_3515, signal_2209}), .c ({signal_3635, signal_2241}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1787 ( .a ({signal_12420, signal_12419}), .b ({signal_3383, signal_2177}), .c ({signal_3515, signal_2209}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1788 ( .a ({signal_12422, signal_12421}), .b ({signal_3230, signal_2145}), .c ({signal_3383, signal_2177}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1789 ( .a ({signal_12424, signal_12423}), .b ({signal_3516, signal_2210}), .c ({signal_3636, signal_2242}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1790 ( .a ({signal_12426, signal_12425}), .b ({signal_3384, signal_2178}), .c ({signal_3516, signal_2210}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1791 ( .a ({signal_12428, signal_12427}), .b ({signal_3231, signal_2146}), .c ({signal_3384, signal_2178}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1792 ( .a ({signal_12430, signal_12429}), .b ({signal_3517, signal_2211}), .c ({signal_3637, signal_2243}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1793 ( .a ({signal_12432, signal_12431}), .b ({signal_3385, signal_2179}), .c ({signal_3517, signal_2211}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1794 ( .a ({signal_12434, signal_12433}), .b ({signal_3232, signal_2147}), .c ({signal_3385, signal_2179}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1795 ( .a ({signal_12436, signal_12435}), .b ({signal_3518, signal_2212}), .c ({signal_3638, signal_2244}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1796 ( .a ({signal_12438, signal_12437}), .b ({signal_3386, signal_2180}), .c ({signal_3518, signal_2212}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1797 ( .a ({signal_12440, signal_12439}), .b ({signal_3233, signal_2148}), .c ({signal_3386, signal_2180}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1798 ( .a ({signal_12442, signal_12441}), .b ({signal_3519, signal_2213}), .c ({signal_3639, signal_2245}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1799 ( .a ({signal_12444, signal_12443}), .b ({signal_3387, signal_2181}), .c ({signal_3519, signal_2213}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1800 ( .a ({signal_12446, signal_12445}), .b ({signal_3234, signal_2149}), .c ({signal_3387, signal_2181}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1801 ( .a ({signal_12448, signal_12447}), .b ({signal_3388, signal_2214}), .c ({signal_3520, signal_2246}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1802 ( .a ({signal_12450, signal_12449}), .b ({signal_3214, signal_2182}), .c ({signal_3388, signal_2214}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1803 ( .a ({signal_12452, signal_12451}), .b ({signal_3145, signal_2150}), .c ({signal_3214, signal_2182}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1804 ( .a ({signal_12454, signal_12453}), .b ({signal_3389, signal_2215}), .c ({signal_3521, signal_2247}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1805 ( .a ({signal_12456, signal_12455}), .b ({signal_3215, signal_2183}), .c ({signal_3389, signal_2215}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1806 ( .a ({signal_12458, signal_12457}), .b ({signal_3146, signal_2151}), .c ({signal_3215, signal_2183}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1807 ( .a ({signal_12460, signal_12459}), .b ({signal_3390, signal_2216}), .c ({signal_3522, signal_2248}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1808 ( .a ({signal_12462, signal_12461}), .b ({signal_3216, signal_2184}), .c ({signal_3390, signal_2216}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1809 ( .a ({signal_12464, signal_12463}), .b ({signal_3147, signal_2152}), .c ({signal_3216, signal_2184}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1810 ( .a ({signal_12466, signal_12465}), .b ({signal_3391, signal_2217}), .c ({signal_3523, signal_2249}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1811 ( .a ({signal_12468, signal_12467}), .b ({signal_3217, signal_2185}), .c ({signal_3391, signal_2217}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1812 ( .a ({signal_12470, signal_12469}), .b ({signal_3148, signal_2153}), .c ({signal_3217, signal_2185}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1813 ( .a ({signal_12472, signal_12471}), .b ({signal_3392, signal_2236}), .c ({signal_3524, signal_2268}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1814 ( .a ({signal_12474, signal_12473}), .b ({signal_3218, signal_2204}), .c ({signal_3392, signal_2236}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1815 ( .a ({signal_12476, signal_12475}), .b ({signal_3144, signal_2172}), .c ({signal_3218, signal_2204}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1816 ( .a ({signal_12478, signal_12477}), .b ({signal_3108, signal_2336}), .c ({signal_3144, signal_2172}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1817 ( .a ({signal_12480, signal_12479}), .b ({signal_3393, signal_2218}), .c ({signal_3525, signal_2250}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1818 ( .a ({signal_12482, signal_12481}), .b ({signal_3219, signal_2186}), .c ({signal_3393, signal_2218}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1819 ( .a ({signal_12484, signal_12483}), .b ({signal_3149, signal_2154}), .c ({signal_3219, signal_2186}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1820 ( .a ({signal_12486, signal_12485}), .b ({signal_3394, signal_2219}), .c ({signal_3526, signal_2251}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1821 ( .a ({signal_12488, signal_12487}), .b ({signal_3220, signal_2187}), .c ({signal_3394, signal_2219}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1822 ( .a ({signal_12490, signal_12489}), .b ({signal_3150, signal_2155}), .c ({signal_3220, signal_2187}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1823 ( .a ({signal_12492, signal_12491}), .b ({signal_3395, signal_2220}), .c ({signal_3527, signal_2252}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1824 ( .a ({signal_12494, signal_12493}), .b ({signal_3221, signal_2188}), .c ({signal_3395, signal_2220}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1825 ( .a ({signal_12496, signal_12495}), .b ({signal_3151, signal_2156}), .c ({signal_3221, signal_2188}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1826 ( .a ({signal_12498, signal_12497}), .b ({signal_3396, signal_2221}), .c ({signal_3528, signal_2253}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1827 ( .a ({signal_12500, signal_12499}), .b ({signal_3222, signal_2189}), .c ({signal_3396, signal_2221}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1828 ( .a ({signal_12502, signal_12501}), .b ({signal_3152, signal_2157}), .c ({signal_3222, signal_2189}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1829 ( .a ({signal_12504, signal_12503}), .b ({signal_3397, signal_2222}), .c ({signal_3529, signal_2254}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1830 ( .a ({signal_12506, signal_12505}), .b ({signal_3223, signal_2190}), .c ({signal_3397, signal_2222}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1831 ( .a ({signal_12508, signal_12507}), .b ({signal_3153, signal_2158}), .c ({signal_3223, signal_2190}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1832 ( .a ({signal_12510, signal_12509}), .b ({signal_3398, signal_2223}), .c ({signal_3530, signal_2255}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1833 ( .a ({signal_12512, signal_12511}), .b ({signal_3224, signal_2191}), .c ({signal_3398, signal_2223}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1834 ( .a ({signal_12514, signal_12513}), .b ({signal_3154, signal_2159}), .c ({signal_3224, signal_2191}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1835 ( .a ({signal_12516, signal_12515}), .b ({signal_3399, signal_2224}), .c ({signal_3531, signal_2256}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1836 ( .a ({signal_12518, signal_12517}), .b ({signal_3225, signal_2192}), .c ({signal_3399, signal_2224}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1837 ( .a ({signal_12520, signal_12519}), .b ({signal_3155, signal_2160}), .c ({signal_3225, signal_2192}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1838 ( .a ({signal_12522, signal_12521}), .b ({signal_3400, signal_2225}), .c ({signal_3532, signal_2257}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1839 ( .a ({signal_12524, signal_12523}), .b ({signal_3226, signal_2193}), .c ({signal_3400, signal_2225}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1840 ( .a ({signal_12526, signal_12525}), .b ({signal_3156, signal_2161}), .c ({signal_3226, signal_2193}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1841 ( .a ({signal_12528, signal_12527}), .b ({signal_3166, signal_2306}), .c ({signal_3227, signal_2142}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1842 ( .a ({signal_12530, signal_12529}), .b ({signal_3167, signal_2307}), .c ({signal_3228, signal_2143}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1843 ( .a ({signal_12532, signal_12531}), .b ({signal_3168, signal_2308}), .c ({signal_3229, signal_2144}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1844 ( .a ({signal_12534, signal_12533}), .b ({signal_3169, signal_2309}), .c ({signal_3230, signal_2145}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1845 ( .a ({signal_12536, signal_12535}), .b ({signal_3170, signal_2310}), .c ({signal_3231, signal_2146}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1846 ( .a ({signal_12538, signal_12537}), .b ({signal_3171, signal_2311}), .c ({signal_3232, signal_2147}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1847 ( .a ({signal_12540, signal_12539}), .b ({signal_3172, signal_2312}), .c ({signal_3233, signal_2148}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1848 ( .a ({signal_12542, signal_12541}), .b ({signal_3173, signal_2313}), .c ({signal_3234, signal_2149}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1849 ( .a ({signal_12544, signal_12543}), .b ({signal_3401, signal_2226}), .c ({signal_3533, signal_2258}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1850 ( .a ({signal_12546, signal_12545}), .b ({signal_3235, signal_2194}), .c ({signal_3401, signal_2226}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1851 ( .a ({signal_12548, signal_12547}), .b ({signal_3157, signal_2162}), .c ({signal_3235, signal_2194}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1852 ( .a ({signal_12550, signal_12549}), .b ({signal_3086, signal_2314}), .c ({signal_3145, signal_2150}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1853 ( .a ({signal_12552, signal_12551}), .b ({signal_3087, signal_2315}), .c ({signal_3146, signal_2151}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1854 ( .a ({signal_12554, signal_12553}), .b ({signal_3088, signal_2316}), .c ({signal_3147, signal_2152}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1855 ( .a ({signal_12556, signal_12555}), .b ({signal_3089, signal_2317}), .c ({signal_3148, signal_2153}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1856 ( .a ({signal_12558, signal_12557}), .b ({signal_3090, signal_2318}), .c ({signal_3149, signal_2154}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1857 ( .a ({signal_12560, signal_12559}), .b ({signal_3091, signal_2319}), .c ({signal_3150, signal_2155}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1858 ( .a ({signal_12562, signal_12561}), .b ({signal_3092, signal_2320}), .c ({signal_3151, signal_2156}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1859 ( .a ({signal_12564, signal_12563}), .b ({signal_3093, signal_2321}), .c ({signal_3152, signal_2157}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1860 ( .a ({signal_12566, signal_12565}), .b ({signal_3094, signal_2322}), .c ({signal_3153, signal_2158}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1861 ( .a ({signal_12568, signal_12567}), .b ({signal_3095, signal_2323}), .c ({signal_3154, signal_2159}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1862 ( .a ({signal_12570, signal_12569}), .b ({signal_3402, signal_2227}), .c ({signal_3534, signal_2259}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1863 ( .a ({signal_12572, signal_12571}), .b ({signal_3236, signal_2195}), .c ({signal_3402, signal_2227}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1864 ( .a ({signal_12574, signal_12573}), .b ({signal_3158, signal_2163}), .c ({signal_3236, signal_2195}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1865 ( .a ({signal_12576, signal_12575}), .b ({signal_3096, signal_2324}), .c ({signal_3155, signal_2160}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1866 ( .a ({signal_12578, signal_12577}), .b ({signal_3097, signal_2325}), .c ({signal_3156, signal_2161}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1867 ( .a ({signal_12580, signal_12579}), .b ({signal_3098, signal_2326}), .c ({signal_3157, signal_2162}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1868 ( .a ({signal_12582, signal_12581}), .b ({signal_3099, signal_2327}), .c ({signal_3158, signal_2163}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1869 ( .a ({signal_12584, signal_12583}), .b ({signal_3100, signal_2328}), .c ({signal_3159, signal_2164}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1870 ( .a ({signal_12586, signal_12585}), .b ({signal_3101, signal_2329}), .c ({signal_3160, signal_2165}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1871 ( .a ({signal_12588, signal_12587}), .b ({signal_3102, signal_2330}), .c ({signal_3161, signal_2166}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1872 ( .a ({signal_12590, signal_12589}), .b ({signal_3103, signal_2331}), .c ({signal_3162, signal_2167}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1873 ( .a ({signal_12592, signal_12591}), .b ({signal_3104, signal_2332}), .c ({signal_3163, signal_2168}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1874 ( .a ({signal_12594, signal_12593}), .b ({signal_3105, signal_2333}), .c ({signal_3164, signal_2169}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1875 ( .a ({signal_12596, signal_12595}), .b ({signal_3403, signal_2237}), .c ({signal_3535, signal_2269}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1876 ( .a ({signal_12598, signal_12597}), .b ({signal_3237, signal_2205}), .c ({signal_3403, signal_2237}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1877 ( .a ({signal_12600, signal_12599}), .b ({signal_3165, signal_2173}), .c ({signal_3237, signal_2205}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1878 ( .a ({signal_12602, signal_12601}), .b ({signal_3109, signal_2337}), .c ({signal_3165, signal_2173}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1879 ( .a ({1'b0, signal_12603}), .b ({signal_3085, signal_2305}), .c ({signal_3166, signal_2306}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1880 ( .a ({1'b0, signal_12604}), .b ({signal_3081, signal_2298}), .c ({signal_3167, signal_2307}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1881 ( .a ({1'b0, signal_12605}), .b ({signal_3082, signal_2299}), .c ({signal_3168, signal_2308}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1882 ( .a ({1'b0, signal_12606}), .b ({signal_3083, signal_2300}), .c ({signal_3169, signal_2309}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1883 ( .a ({1'b0, signal_12607}), .b ({signal_3048, signal_1842}), .c ({signal_3170, signal_2310}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1884 ( .a ({1'b0, signal_12608}), .b ({signal_3049, signal_1843}), .c ({signal_3171, signal_2311}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1885 ( .a ({1'b0, signal_12609}), .b ({signal_3084, signal_2303}), .c ({signal_3172, signal_2312}) ) ;
    xor_GHPC #(.low_latency(1), .pipeline(1)) cell_1886 ( .a ({1'b0, signal_12610}), .b ({signal_3050, signal_1845}), .c ({signal_3173, signal_2313}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1895 ( .s (signal_12611), .b ({signal_12596, signal_12595}), .a ({signal_3535, signal_2269}), .c ({signal_3640, signal_2037}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1896 ( .s (signal_12612), .b ({signal_12472, signal_12471}), .a ({signal_3524, signal_2268}), .c ({signal_3641, signal_2036}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1897 ( .s (signal_12613), .b ({signal_12404, signal_12403}), .a ({signal_3513, signal_2267}), .c ({signal_3642, signal_2035}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1898 ( .s (signal_12614), .b ({signal_12368, signal_12367}), .a ({signal_3510, signal_2266}), .c ({signal_3643, signal_2034}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1899 ( .s (signal_12615), .b ({signal_12358, signal_12357}), .a ({signal_3509, signal_2265}), .c ({signal_3644, signal_2033}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1900 ( .s (signal_12616), .b ({signal_12356, signal_12355}), .a ({signal_3508, signal_2264}), .c ({signal_3645, signal_2032}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1901 ( .s (signal_12612), .b ({signal_12354, signal_12353}), .a ({signal_3507, signal_2263}), .c ({signal_3646, signal_2031}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1902 ( .s (signal_12614), .b ({signal_12352, signal_12351}), .a ({signal_3506, signal_2262}), .c ({signal_3647, signal_2030}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1903 ( .s (signal_12611), .b ({signal_12350, signal_12349}), .a ({signal_3505, signal_2261}), .c ({signal_3648, signal_2029}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1904 ( .s (signal_12612), .b ({signal_12348, signal_12347}), .a ({signal_3504, signal_2260}), .c ({signal_3649, signal_2028}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1905 ( .s (signal_12613), .b ({signal_12570, signal_12569}), .a ({signal_3534, signal_2259}), .c ({signal_3650, signal_2027}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1906 ( .s (signal_12614), .b ({signal_12544, signal_12543}), .a ({signal_3533, signal_2258}), .c ({signal_3651, signal_2026}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1907 ( .s (signal_12615), .b ({signal_12522, signal_12521}), .a ({signal_3532, signal_2257}), .c ({signal_3652, signal_2025}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1908 ( .s (signal_12616), .b ({signal_12516, signal_12515}), .a ({signal_3531, signal_2256}), .c ({signal_3653, signal_2024}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1909 ( .s (signal_12615), .b ({signal_12510, signal_12509}), .a ({signal_3530, signal_2255}), .c ({signal_3654, signal_2023}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1910 ( .s (signal_12615), .b ({signal_12504, signal_12503}), .a ({signal_3529, signal_2254}), .c ({signal_3655, signal_2022}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1911 ( .s (signal_12611), .b ({signal_12498, signal_12497}), .a ({signal_3528, signal_2253}), .c ({signal_3656, signal_2021}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1912 ( .s (signal_12612), .b ({signal_12492, signal_12491}), .a ({signal_3527, signal_2252}), .c ({signal_3657, signal_2020}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1913 ( .s (signal_12613), .b ({signal_12486, signal_12485}), .a ({signal_3526, signal_2251}), .c ({signal_3658, signal_2019}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1914 ( .s (signal_12614), .b ({signal_12480, signal_12479}), .a ({signal_3525, signal_2250}), .c ({signal_3659, signal_2018}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1915 ( .s (signal_12616), .b ({signal_12466, signal_12465}), .a ({signal_3523, signal_2249}), .c ({signal_3660, signal_2017}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1916 ( .s (signal_12616), .b ({signal_12460, signal_12459}), .a ({signal_3522, signal_2248}), .c ({signal_3661, signal_2016}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1917 ( .s (signal_12611), .b ({signal_12454, signal_12453}), .a ({signal_3521, signal_2247}), .c ({signal_3662, signal_2015}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1918 ( .s (signal_12612), .b ({signal_12448, signal_12447}), .a ({signal_3520, signal_2246}), .c ({signal_3663, signal_2014}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1919 ( .s (signal_12613), .b ({signal_12442, signal_12441}), .a ({signal_3639, signal_2245}), .c ({signal_3736, signal_2013}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1920 ( .s (signal_12614), .b ({signal_12436, signal_12435}), .a ({signal_3638, signal_2244}), .c ({signal_3737, signal_2012}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1921 ( .s (signal_12615), .b ({signal_12430, signal_12429}), .a ({signal_3637, signal_2243}), .c ({signal_3738, signal_2011}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1922 ( .s (signal_12616), .b ({signal_12424, signal_12423}), .a ({signal_3636, signal_2242}), .c ({signal_3739, signal_2010}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1923 ( .s (signal_12611), .b ({signal_12418, signal_12417}), .a ({signal_3635, signal_2241}), .c ({signal_3740, signal_2009}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1924 ( .s (signal_12611), .b ({signal_12412, signal_12411}), .a ({signal_3634, signal_2240}), .c ({signal_3741, signal_2008}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1925 ( .s (signal_12612), .b ({signal_12398, signal_12397}), .a ({signal_3633, signal_2239}), .c ({signal_3742, signal_2007}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1926 ( .s (signal_12613), .b ({signal_12392, signal_12391}), .a ({signal_3632, signal_2238}), .c ({signal_3743, signal_2006}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1927 ( .s (signal_12612), .b ({signal_12598, signal_12597}), .a ({signal_3403, signal_2237}), .c ({signal_3536, signal_2005}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1928 ( .s (signal_12613), .b ({signal_12474, signal_12473}), .a ({signal_3392, signal_2236}), .c ({signal_3537, signal_2004}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1929 ( .s (signal_12614), .b ({signal_12406, signal_12405}), .a ({signal_3381, signal_2235}), .c ({signal_3538, signal_2003}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1930 ( .s (signal_12615), .b ({signal_12386, signal_12385}), .a ({signal_3378, signal_2234}), .c ({signal_3539, signal_2002}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1931 ( .s (signal_12616), .b ({signal_12382, signal_12381}), .a ({signal_3377, signal_2233}), .c ({signal_3540, signal_2001}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1932 ( .s (signal_12611), .b ({signal_12378, signal_12377}), .a ({signal_3376, signal_2232}), .c ({signal_3541, signal_2000}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1933 ( .s (signal_12612), .b ({signal_12374, signal_12373}), .a ({signal_3375, signal_2231}), .c ({signal_3542, signal_1999}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1934 ( .s (signal_12613), .b ({signal_12370, signal_12369}), .a ({signal_3374, signal_2230}), .c ({signal_3543, signal_1998}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1935 ( .s (signal_12614), .b ({signal_12364, signal_12363}), .a ({signal_3373, signal_2229}), .c ({signal_3544, signal_1997}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1936 ( .s (signal_12615), .b ({signal_12360, signal_12359}), .a ({signal_3372, signal_2228}), .c ({signal_3545, signal_1996}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1937 ( .s (signal_12616), .b ({signal_12572, signal_12571}), .a ({signal_3402, signal_2227}), .c ({signal_3546, signal_1995}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1938 ( .s (signal_12611), .b ({signal_12546, signal_12545}), .a ({signal_3401, signal_2226}), .c ({signal_3547, signal_1994}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1939 ( .s (signal_12616), .b ({signal_12524, signal_12523}), .a ({signal_3400, signal_2225}), .c ({signal_3548, signal_1993}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1940 ( .s (signal_12616), .b ({signal_12518, signal_12517}), .a ({signal_3399, signal_2224}), .c ({signal_3549, signal_1992}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1941 ( .s (signal_12616), .b ({signal_12512, signal_12511}), .a ({signal_3398, signal_2223}), .c ({signal_3550, signal_1991}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1942 ( .s (signal_12616), .b ({signal_12506, signal_12505}), .a ({signal_3397, signal_2222}), .c ({signal_3551, signal_1990}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1943 ( .s (signal_12616), .b ({signal_12500, signal_12499}), .a ({signal_3396, signal_2221}), .c ({signal_3552, signal_1989}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1944 ( .s (signal_12616), .b ({signal_12494, signal_12493}), .a ({signal_3395, signal_2220}), .c ({signal_3553, signal_1988}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1945 ( .s (signal_12616), .b ({signal_12488, signal_12487}), .a ({signal_3394, signal_2219}), .c ({signal_3554, signal_1987}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1946 ( .s (signal_12616), .b ({signal_12482, signal_12481}), .a ({signal_3393, signal_2218}), .c ({signal_3555, signal_1986}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1947 ( .s (signal_12616), .b ({signal_12468, signal_12467}), .a ({signal_3391, signal_2217}), .c ({signal_3556, signal_1985}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1948 ( .s (signal_12616), .b ({signal_12462, signal_12461}), .a ({signal_3390, signal_2216}), .c ({signal_3557, signal_1984}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1949 ( .s (signal_12616), .b ({signal_12456, signal_12455}), .a ({signal_3389, signal_2215}), .c ({signal_3558, signal_1983}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1950 ( .s (signal_12616), .b ({signal_12450, signal_12449}), .a ({signal_3388, signal_2214}), .c ({signal_3559, signal_1982}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1951 ( .s (signal_12615), .b ({signal_12444, signal_12443}), .a ({signal_3519, signal_2213}), .c ({signal_3664, signal_1981}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1952 ( .s (signal_12615), .b ({signal_12438, signal_12437}), .a ({signal_3518, signal_2212}), .c ({signal_3665, signal_1980}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1953 ( .s (signal_12615), .b ({signal_12432, signal_12431}), .a ({signal_3517, signal_2211}), .c ({signal_3666, signal_1979}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1954 ( .s (signal_12615), .b ({signal_12426, signal_12425}), .a ({signal_3516, signal_2210}), .c ({signal_3667, signal_1978}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1955 ( .s (signal_12615), .b ({signal_12420, signal_12419}), .a ({signal_3515, signal_2209}), .c ({signal_3668, signal_1977}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1956 ( .s (signal_12615), .b ({signal_12414, signal_12413}), .a ({signal_3514, signal_2208}), .c ({signal_3669, signal_1976}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1957 ( .s (signal_12615), .b ({signal_12400, signal_12399}), .a ({signal_3512, signal_2207}), .c ({signal_3670, signal_1975}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1958 ( .s (signal_12615), .b ({signal_12394, signal_12393}), .a ({signal_3511, signal_2206}), .c ({signal_3671, signal_1974}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1959 ( .s (signal_12615), .b ({signal_12600, signal_12599}), .a ({signal_3237, signal_2205}), .c ({signal_3404, signal_1973}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1960 ( .s (signal_12615), .b ({signal_12476, signal_12475}), .a ({signal_3218, signal_2204}), .c ({signal_3405, signal_1972}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1961 ( .s (signal_12615), .b ({signal_12408, signal_12407}), .a ({signal_3213, signal_2203}), .c ({signal_3406, signal_1971}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1962 ( .s (signal_12615), .b ({signal_12388, signal_12387}), .a ({signal_3212, signal_2202}), .c ({signal_3407, signal_1970}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1963 ( .s (signal_12614), .b ({signal_12384, signal_12383}), .a ({signal_3211, signal_2201}), .c ({signal_3408, signal_1969}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1964 ( .s (signal_12614), .b ({signal_12380, signal_12379}), .a ({signal_3210, signal_2200}), .c ({signal_3409, signal_1968}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1965 ( .s (signal_12614), .b ({signal_12376, signal_12375}), .a ({signal_3209, signal_2199}), .c ({signal_3410, signal_1967}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1966 ( .s (signal_12614), .b ({signal_12372, signal_12371}), .a ({signal_3208, signal_2198}), .c ({signal_3411, signal_1966}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1967 ( .s (signal_12614), .b ({signal_12366, signal_12365}), .a ({signal_3207, signal_2197}), .c ({signal_3412, signal_1965}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1968 ( .s (signal_12614), .b ({signal_12362, signal_12361}), .a ({signal_3206, signal_2196}), .c ({signal_3413, signal_1964}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1969 ( .s (signal_12614), .b ({signal_12574, signal_12573}), .a ({signal_3236, signal_2195}), .c ({signal_3414, signal_1963}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1970 ( .s (signal_12614), .b ({signal_12548, signal_12547}), .a ({signal_3235, signal_2194}), .c ({signal_3415, signal_1962}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1971 ( .s (signal_12614), .b ({signal_12526, signal_12525}), .a ({signal_3226, signal_2193}), .c ({signal_3416, signal_1961}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1972 ( .s (signal_12614), .b ({signal_12520, signal_12519}), .a ({signal_3225, signal_2192}), .c ({signal_3417, signal_1960}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1973 ( .s (signal_12614), .b ({signal_12514, signal_12513}), .a ({signal_3224, signal_2191}), .c ({signal_3418, signal_1959}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1974 ( .s (signal_12614), .b ({signal_12508, signal_12507}), .a ({signal_3223, signal_2190}), .c ({signal_3419, signal_1958}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1975 ( .s (signal_12613), .b ({signal_12502, signal_12501}), .a ({signal_3222, signal_2189}), .c ({signal_3420, signal_1957}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1976 ( .s (signal_12613), .b ({signal_12496, signal_12495}), .a ({signal_3221, signal_2188}), .c ({signal_3421, signal_1956}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1977 ( .s (signal_12613), .b ({signal_12490, signal_12489}), .a ({signal_3220, signal_2187}), .c ({signal_3422, signal_1955}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1978 ( .s (signal_12613), .b ({signal_12484, signal_12483}), .a ({signal_3219, signal_2186}), .c ({signal_3423, signal_1954}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1979 ( .s (signal_12613), .b ({signal_12470, signal_12469}), .a ({signal_3217, signal_2185}), .c ({signal_3424, signal_1953}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1980 ( .s (signal_12613), .b ({signal_12464, signal_12463}), .a ({signal_3216, signal_2184}), .c ({signal_3425, signal_1952}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1981 ( .s (signal_12613), .b ({signal_12458, signal_12457}), .a ({signal_3215, signal_2183}), .c ({signal_3426, signal_1951}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1982 ( .s (signal_12613), .b ({signal_12452, signal_12451}), .a ({signal_3214, signal_2182}), .c ({signal_3427, signal_1950}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1983 ( .s (signal_12613), .b ({signal_12446, signal_12445}), .a ({signal_3387, signal_2181}), .c ({signal_3560, signal_1949}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1984 ( .s (signal_12613), .b ({signal_12440, signal_12439}), .a ({signal_3386, signal_2180}), .c ({signal_3561, signal_1948}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1985 ( .s (signal_12613), .b ({signal_12434, signal_12433}), .a ({signal_3385, signal_2179}), .c ({signal_3562, signal_1947}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1986 ( .s (signal_12613), .b ({signal_12428, signal_12427}), .a ({signal_3384, signal_2178}), .c ({signal_3563, signal_1946}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1987 ( .s (signal_12612), .b ({signal_12422, signal_12421}), .a ({signal_3383, signal_2177}), .c ({signal_3564, signal_1945}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1988 ( .s (signal_12612), .b ({signal_12416, signal_12415}), .a ({signal_3382, signal_2176}), .c ({signal_3565, signal_1944}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1989 ( .s (signal_12612), .b ({signal_12402, signal_12401}), .a ({signal_3380, signal_2175}), .c ({signal_3566, signal_1943}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1990 ( .s (signal_12612), .b ({signal_12396, signal_12395}), .a ({signal_3379, signal_2174}), .c ({signal_3567, signal_1942}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1991 ( .s (signal_12612), .b ({signal_12602, signal_12601}), .a ({signal_3165, signal_2173}), .c ({signal_3238, signal_1941}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1992 ( .s (signal_12612), .b ({signal_12478, signal_12477}), .a ({signal_3144, signal_2172}), .c ({signal_3239, signal_1940}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1993 ( .s (signal_12612), .b ({signal_12410, signal_12409}), .a ({signal_3143, signal_2171}), .c ({signal_3240, signal_1939}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1994 ( .s (signal_12612), .b ({signal_12390, signal_12389}), .a ({signal_3142, signal_2170}), .c ({signal_3241, signal_1938}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1995 ( .s (signal_12612), .b ({signal_12594, signal_12593}), .a ({signal_3164, signal_2169}), .c ({signal_3242, signal_1937}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1996 ( .s (signal_12612), .b ({signal_12592, signal_12591}), .a ({signal_3163, signal_2168}), .c ({signal_3243, signal_1936}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1997 ( .s (signal_12612), .b ({signal_12590, signal_12589}), .a ({signal_3162, signal_2167}), .c ({signal_3244, signal_1935}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1998 ( .s (signal_12612), .b ({signal_12588, signal_12587}), .a ({signal_3161, signal_2166}), .c ({signal_3245, signal_1934}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_1999 ( .s (signal_12611), .b ({signal_12586, signal_12585}), .a ({signal_3160, signal_2165}), .c ({signal_3246, signal_1933}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2000 ( .s (signal_12611), .b ({signal_12584, signal_12583}), .a ({signal_3159, signal_2164}), .c ({signal_3247, signal_1932}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2001 ( .s (signal_12611), .b ({signal_12582, signal_12581}), .a ({signal_3158, signal_2163}), .c ({signal_3248, signal_1931}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2002 ( .s (signal_12611), .b ({signal_12580, signal_12579}), .a ({signal_3157, signal_2162}), .c ({signal_3249, signal_1930}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2003 ( .s (signal_12611), .b ({signal_12578, signal_12577}), .a ({signal_3156, signal_2161}), .c ({signal_3250, signal_1929}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2004 ( .s (signal_12611), .b ({signal_12576, signal_12575}), .a ({signal_3155, signal_2160}), .c ({signal_3251, signal_1928}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2005 ( .s (signal_12611), .b ({signal_12568, signal_12567}), .a ({signal_3154, signal_2159}), .c ({signal_3252, signal_1927}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2006 ( .s (signal_12611), .b ({signal_12566, signal_12565}), .a ({signal_3153, signal_2158}), .c ({signal_3253, signal_1926}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2007 ( .s (signal_12611), .b ({signal_12564, signal_12563}), .a ({signal_3152, signal_2157}), .c ({signal_3254, signal_1925}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2008 ( .s (signal_12611), .b ({signal_12562, signal_12561}), .a ({signal_3151, signal_2156}), .c ({signal_3255, signal_1924}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2009 ( .s (signal_12611), .b ({signal_12560, signal_12559}), .a ({signal_3150, signal_2155}), .c ({signal_3256, signal_1923}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2010 ( .s (signal_12611), .b ({signal_12558, signal_12557}), .a ({signal_3149, signal_2154}), .c ({signal_3257, signal_1922}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2011 ( .s (signal_12617), .b ({signal_12556, signal_12555}), .a ({signal_3148, signal_2153}), .c ({signal_3258, signal_1921}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2012 ( .s (signal_12617), .b ({signal_12554, signal_12553}), .a ({signal_3147, signal_2152}), .c ({signal_3259, signal_1920}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2013 ( .s (signal_12617), .b ({signal_12552, signal_12551}), .a ({signal_3146, signal_2151}), .c ({signal_3260, signal_1919}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2014 ( .s (signal_12617), .b ({signal_12550, signal_12549}), .a ({signal_3145, signal_2150}), .c ({signal_3261, signal_1918}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2015 ( .s (signal_12617), .b ({signal_12542, signal_12541}), .a ({signal_3234, signal_2149}), .c ({signal_3428, signal_1917}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2016 ( .s (signal_12617), .b ({signal_12540, signal_12539}), .a ({signal_3233, signal_2148}), .c ({signal_3429, signal_1916}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2017 ( .s (signal_12617), .b ({signal_12538, signal_12537}), .a ({signal_3232, signal_2147}), .c ({signal_3430, signal_1915}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2018 ( .s (signal_12617), .b ({signal_12536, signal_12535}), .a ({signal_3231, signal_2146}), .c ({signal_3431, signal_1914}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2019 ( .s (signal_12617), .b ({signal_12534, signal_12533}), .a ({signal_3230, signal_2145}), .c ({signal_3432, signal_1913}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2020 ( .s (signal_12617), .b ({signal_12532, signal_12531}), .a ({signal_3229, signal_2144}), .c ({signal_3433, signal_1912}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2021 ( .s (signal_12617), .b ({signal_12530, signal_12529}), .a ({signal_3228, signal_2143}), .c ({signal_3434, signal_1911}) ) ;
    mux2_masked #(.low_latency(1), .pipeline(1)) cell_2022 ( .s (signal_12617), .b ({signal_12528, signal_12527}), .a ({signal_3227, signal_2142}), .c ({signal_3435, signal_1910}) ) ;
    AES_step2_ANF #(.low_latency(1), .pipeline(1)) cell_2061 ( .in0 ({signal_908, signal_788, signal_1841, signal_1840, signal_1839, signal_1837, signal_1836, signal_1835, signal_1834, signal_1833, signal_1832, signal_1831, signal_1829, signal_1828, signal_1827, signal_1826, signal_1825, signal_1824, signal_1823, signal_1821, signal_1820, signal_1819, signal_1818, signal_1817, signal_1816, signal_1815, signal_1813, signal_1812, signal_1811, signal_1810, signal_1148, signal_1028}), .in1 ({signal_3043, signal_3042, signal_2723, signal_2724, signal_2725, signal_2727, signal_2728, signal_2729, signal_2730, signal_2722, signal_2731, signal_2732, signal_2734, signal_2735, signal_2736, signal_2737, signal_2738, signal_2739, signal_2740, signal_2742, signal_2743, signal_2744, signal_2745, signal_2746, signal_2747, signal_2748, signal_2750, signal_2751, signal_2752, signal_2753, signal_3045, signal_3044}), .clk (clk), .r ({Fresh[8191], Fresh[8190], Fresh[8189], Fresh[8188], Fresh[8187], Fresh[8186], Fresh[8185], Fresh[8184], Fresh[8183], Fresh[8182], Fresh[8181], Fresh[8180], Fresh[8179], Fresh[8178], Fresh[8177], Fresh[8176], Fresh[8175], Fresh[8174], Fresh[8173], Fresh[8172], Fresh[8171], Fresh[8170], Fresh[8169], Fresh[8168], Fresh[8167], Fresh[8166], Fresh[8165], Fresh[8164], Fresh[8163], Fresh[8162], Fresh[8161], Fresh[8160], Fresh[8159], Fresh[8158], Fresh[8157], Fresh[8156], Fresh[8155], Fresh[8154], Fresh[8153], Fresh[8152], Fresh[8151], Fresh[8150], Fresh[8149], Fresh[8148], Fresh[8147], Fresh[8146], Fresh[8145], Fresh[8144], Fresh[8143], Fresh[8142], Fresh[8141], Fresh[8140], Fresh[8139], Fresh[8138], Fresh[8137], Fresh[8136], Fresh[8135], Fresh[8134], Fresh[8133], Fresh[8132], Fresh[8131], Fresh[8130], Fresh[8129], Fresh[8128], Fresh[8127], Fresh[8126], Fresh[8125], Fresh[8124], Fresh[8123], Fresh[8122], Fresh[8121], Fresh[8120], Fresh[8119], Fresh[8118], Fresh[8117], Fresh[8116], Fresh[8115], Fresh[8114], Fresh[8113], Fresh[8112], Fresh[8111], Fresh[8110], Fresh[8109], Fresh[8108], Fresh[8107], Fresh[8106], Fresh[8105], Fresh[8104], Fresh[8103], Fresh[8102], Fresh[8101], Fresh[8100], Fresh[8099], Fresh[8098], Fresh[8097], Fresh[8096], Fresh[8095], Fresh[8094], Fresh[8093], Fresh[8092], Fresh[8091], Fresh[8090], Fresh[8089], Fresh[8088], Fresh[8087], Fresh[8086], Fresh[8085], Fresh[8084], Fresh[8083], Fresh[8082], Fresh[8081], Fresh[8080], Fresh[8079], Fresh[8078], Fresh[8077], Fresh[8076], Fresh[8075], Fresh[8074], Fresh[8073], Fresh[8072], Fresh[8071], Fresh[8070], Fresh[8069], Fresh[8068], Fresh[8067], Fresh[8066], Fresh[8065], Fresh[8064], Fresh[8063], Fresh[8062], Fresh[8061], Fresh[8060], Fresh[8059], Fresh[8058], Fresh[8057], Fresh[8056], Fresh[8055], Fresh[8054], Fresh[8053], Fresh[8052], Fresh[8051], Fresh[8050], Fresh[8049], Fresh[8048], Fresh[8047], Fresh[8046], Fresh[8045], Fresh[8044], Fresh[8043], Fresh[8042], Fresh[8041], Fresh[8040], Fresh[8039], Fresh[8038], Fresh[8037], Fresh[8036], Fresh[8035], Fresh[8034], Fresh[8033], Fresh[8032], Fresh[8031], Fresh[8030], Fresh[8029], Fresh[8028], Fresh[8027], Fresh[8026], Fresh[8025], Fresh[8024], Fresh[8023], Fresh[8022], Fresh[8021], Fresh[8020], Fresh[8019], Fresh[8018], Fresh[8017], Fresh[8016], Fresh[8015], Fresh[8014], Fresh[8013], Fresh[8012], Fresh[8011], Fresh[8010], Fresh[8009], Fresh[8008], Fresh[8007], Fresh[8006], Fresh[8005], Fresh[8004], Fresh[8003], Fresh[8002], Fresh[8001], Fresh[8000], Fresh[7999], Fresh[7998], Fresh[7997], Fresh[7996], Fresh[7995], Fresh[7994], Fresh[7993], Fresh[7992], Fresh[7991], Fresh[7990], Fresh[7989], Fresh[7988], Fresh[7987], Fresh[7986], Fresh[7985], Fresh[7984], Fresh[7983], Fresh[7982], Fresh[7981], Fresh[7980], Fresh[7979], Fresh[7978], Fresh[7977], Fresh[7976], Fresh[7975], Fresh[7974], Fresh[7973], Fresh[7972], Fresh[7971], Fresh[7970], Fresh[7969], Fresh[7968], Fresh[7967], Fresh[7966], Fresh[7965], Fresh[7964], Fresh[7963], Fresh[7962], Fresh[7961], Fresh[7960], Fresh[7959], Fresh[7958], Fresh[7957], Fresh[7956], Fresh[7955], Fresh[7954], Fresh[7953], Fresh[7952], Fresh[7951], Fresh[7950], Fresh[7949], Fresh[7948], Fresh[7947], Fresh[7946], Fresh[7945], Fresh[7944], Fresh[7943], Fresh[7942], Fresh[7941], Fresh[7940], Fresh[7939], Fresh[7938], Fresh[7937], Fresh[7936], Fresh[7935], Fresh[7934], Fresh[7933], Fresh[7932], Fresh[7931], Fresh[7930], Fresh[7929], Fresh[7928], Fresh[7927], Fresh[7926], Fresh[7925], Fresh[7924], Fresh[7923], Fresh[7922], Fresh[7921], Fresh[7920], Fresh[7919], Fresh[7918], Fresh[7917], Fresh[7916], Fresh[7915], Fresh[7914], Fresh[7913], Fresh[7912], Fresh[7911], Fresh[7910], Fresh[7909], Fresh[7908], Fresh[7907], Fresh[7906], Fresh[7905], Fresh[7904], Fresh[7903], Fresh[7902], Fresh[7901], Fresh[7900], Fresh[7899], Fresh[7898], Fresh[7897], Fresh[7896], Fresh[7895], Fresh[7894], Fresh[7893], Fresh[7892], Fresh[7891], Fresh[7890], Fresh[7889], Fresh[7888], Fresh[7887], Fresh[7886], Fresh[7885], Fresh[7884], Fresh[7883], Fresh[7882], Fresh[7881], Fresh[7880], Fresh[7879], Fresh[7878], Fresh[7877], Fresh[7876], Fresh[7875], Fresh[7874], Fresh[7873], Fresh[7872], Fresh[7871], Fresh[7870], Fresh[7869], Fresh[7868], Fresh[7867], Fresh[7866], Fresh[7865], Fresh[7864], Fresh[7863], Fresh[7862], Fresh[7861], Fresh[7860], Fresh[7859], Fresh[7858], Fresh[7857], Fresh[7856], Fresh[7855], Fresh[7854], Fresh[7853], Fresh[7852], Fresh[7851], Fresh[7850], Fresh[7849], Fresh[7848], Fresh[7847], Fresh[7846], Fresh[7845], Fresh[7844], Fresh[7843], Fresh[7842], Fresh[7841], Fresh[7840], Fresh[7839], Fresh[7838], Fresh[7837], Fresh[7836], Fresh[7835], Fresh[7834], Fresh[7833], Fresh[7832], Fresh[7831], Fresh[7830], Fresh[7829], Fresh[7828], Fresh[7827], Fresh[7826], Fresh[7825], Fresh[7824], Fresh[7823], Fresh[7822], Fresh[7821], Fresh[7820], Fresh[7819], Fresh[7818], Fresh[7817], Fresh[7816], Fresh[7815], Fresh[7814], Fresh[7813], Fresh[7812], Fresh[7811], Fresh[7810], Fresh[7809], Fresh[7808], Fresh[7807], Fresh[7806], Fresh[7805], Fresh[7804], Fresh[7803], Fresh[7802], Fresh[7801], Fresh[7800], Fresh[7799], Fresh[7798], Fresh[7797], Fresh[7796], Fresh[7795], Fresh[7794], Fresh[7793], Fresh[7792], Fresh[7791], Fresh[7790], Fresh[7789], Fresh[7788], Fresh[7787], Fresh[7786], Fresh[7785], Fresh[7784], Fresh[7783], Fresh[7782], Fresh[7781], Fresh[7780], Fresh[7779], Fresh[7778], Fresh[7777], Fresh[7776], Fresh[7775], Fresh[7774], Fresh[7773], Fresh[7772], Fresh[7771], Fresh[7770], Fresh[7769], Fresh[7768], Fresh[7767], Fresh[7766], Fresh[7765], Fresh[7764], Fresh[7763], Fresh[7762], Fresh[7761], Fresh[7760], Fresh[7759], Fresh[7758], Fresh[7757], Fresh[7756], Fresh[7755], Fresh[7754], Fresh[7753], Fresh[7752], Fresh[7751], Fresh[7750], Fresh[7749], Fresh[7748], Fresh[7747], Fresh[7746], Fresh[7745], Fresh[7744], Fresh[7743], Fresh[7742], Fresh[7741], Fresh[7740], Fresh[7739], Fresh[7738], Fresh[7737], Fresh[7736], Fresh[7735], Fresh[7734], Fresh[7733], Fresh[7732], Fresh[7731], Fresh[7730], Fresh[7729], Fresh[7728], Fresh[7727], Fresh[7726], Fresh[7725], Fresh[7724], Fresh[7723], Fresh[7722], Fresh[7721], Fresh[7720], Fresh[7719], Fresh[7718], Fresh[7717], Fresh[7716], Fresh[7715], Fresh[7714], Fresh[7713], Fresh[7712], Fresh[7711], Fresh[7710], Fresh[7709], Fresh[7708], Fresh[7707], Fresh[7706], Fresh[7705], Fresh[7704], Fresh[7703], Fresh[7702], Fresh[7701], Fresh[7700], Fresh[7699], Fresh[7698], Fresh[7697], Fresh[7696], Fresh[7695], Fresh[7694], Fresh[7693], Fresh[7692], Fresh[7691], Fresh[7690], Fresh[7689], Fresh[7688], Fresh[7687], Fresh[7686], Fresh[7685], Fresh[7684], Fresh[7683], Fresh[7682], Fresh[7681], Fresh[7680], Fresh[7679], Fresh[7678], Fresh[7677], Fresh[7676], Fresh[7675], Fresh[7674], Fresh[7673], Fresh[7672], Fresh[7671], Fresh[7670], Fresh[7669], Fresh[7668], Fresh[7667], Fresh[7666], Fresh[7665], Fresh[7664], Fresh[7663], Fresh[7662], Fresh[7661], Fresh[7660], Fresh[7659], Fresh[7658], Fresh[7657], Fresh[7656], Fresh[7655], Fresh[7654], Fresh[7653], Fresh[7652], Fresh[7651], Fresh[7650], Fresh[7649], Fresh[7648], Fresh[7647], Fresh[7646], Fresh[7645], Fresh[7644], Fresh[7643], Fresh[7642], Fresh[7641], Fresh[7640], Fresh[7639], Fresh[7638], Fresh[7637], Fresh[7636], Fresh[7635], Fresh[7634], Fresh[7633], Fresh[7632], Fresh[7631], Fresh[7630], Fresh[7629], Fresh[7628], Fresh[7627], Fresh[7626], Fresh[7625], Fresh[7624], Fresh[7623], Fresh[7622], Fresh[7621], Fresh[7620], Fresh[7619], Fresh[7618], Fresh[7617], Fresh[7616], Fresh[7615], Fresh[7614], Fresh[7613], Fresh[7612], Fresh[7611], Fresh[7610], Fresh[7609], Fresh[7608], Fresh[7607], Fresh[7606], Fresh[7605], Fresh[7604], Fresh[7603], Fresh[7602], Fresh[7601], Fresh[7600], Fresh[7599], Fresh[7598], Fresh[7597], Fresh[7596], Fresh[7595], Fresh[7594], Fresh[7593], Fresh[7592], Fresh[7591], Fresh[7590], Fresh[7589], Fresh[7588], Fresh[7587], Fresh[7586], Fresh[7585], Fresh[7584], Fresh[7583], Fresh[7582], Fresh[7581], Fresh[7580], Fresh[7579], Fresh[7578], Fresh[7577], Fresh[7576], Fresh[7575], Fresh[7574], Fresh[7573], Fresh[7572], Fresh[7571], Fresh[7570], Fresh[7569], Fresh[7568], Fresh[7567], Fresh[7566], Fresh[7565], Fresh[7564], Fresh[7563], Fresh[7562], Fresh[7561], Fresh[7560], Fresh[7559], Fresh[7558], Fresh[7557], Fresh[7556], Fresh[7555], Fresh[7554], Fresh[7553], Fresh[7552], Fresh[7551], Fresh[7550], Fresh[7549], Fresh[7548], Fresh[7547], Fresh[7546], Fresh[7545], Fresh[7544], Fresh[7543], Fresh[7542], Fresh[7541], Fresh[7540], Fresh[7539], Fresh[7538], Fresh[7537], Fresh[7536], Fresh[7535], Fresh[7534], Fresh[7533], Fresh[7532], Fresh[7531], Fresh[7530], Fresh[7529], Fresh[7528], Fresh[7527], Fresh[7526], Fresh[7525], Fresh[7524], Fresh[7523], Fresh[7522], Fresh[7521], Fresh[7520], Fresh[7519], Fresh[7518], Fresh[7517], Fresh[7516], Fresh[7515], Fresh[7514], Fresh[7513], Fresh[7512], Fresh[7511], Fresh[7510], Fresh[7509], Fresh[7508], Fresh[7507], Fresh[7506], Fresh[7505], Fresh[7504], Fresh[7503], Fresh[7502], Fresh[7501], Fresh[7500], Fresh[7499], Fresh[7498], Fresh[7497], Fresh[7496], Fresh[7495], Fresh[7494], Fresh[7493], Fresh[7492], Fresh[7491], Fresh[7490], Fresh[7489], Fresh[7488], Fresh[7487], Fresh[7486], Fresh[7485], Fresh[7484], Fresh[7483], Fresh[7482], Fresh[7481], Fresh[7480], Fresh[7479], Fresh[7478], Fresh[7477], Fresh[7476], Fresh[7475], Fresh[7474], Fresh[7473], Fresh[7472], Fresh[7471], Fresh[7470], Fresh[7469], Fresh[7468], Fresh[7467], Fresh[7466], Fresh[7465], Fresh[7464], Fresh[7463], Fresh[7462], Fresh[7461], Fresh[7460], Fresh[7459], Fresh[7458], Fresh[7457], Fresh[7456], Fresh[7455], Fresh[7454], Fresh[7453], Fresh[7452], Fresh[7451], Fresh[7450], Fresh[7449], Fresh[7448], Fresh[7447], Fresh[7446], Fresh[7445], Fresh[7444], Fresh[7443], Fresh[7442], Fresh[7441], Fresh[7440], Fresh[7439], Fresh[7438], Fresh[7437], Fresh[7436], Fresh[7435], Fresh[7434], Fresh[7433], Fresh[7432], Fresh[7431], Fresh[7430], Fresh[7429], Fresh[7428], Fresh[7427], Fresh[7426], Fresh[7425], Fresh[7424], Fresh[7423], Fresh[7422], Fresh[7421], Fresh[7420], Fresh[7419], Fresh[7418], Fresh[7417], Fresh[7416], Fresh[7415], Fresh[7414], Fresh[7413], Fresh[7412], Fresh[7411], Fresh[7410], Fresh[7409], Fresh[7408], Fresh[7407], Fresh[7406], Fresh[7405], Fresh[7404], Fresh[7403], Fresh[7402], Fresh[7401], Fresh[7400], Fresh[7399], Fresh[7398], Fresh[7397], Fresh[7396], Fresh[7395], Fresh[7394], Fresh[7393], Fresh[7392], Fresh[7391], Fresh[7390], Fresh[7389], Fresh[7388], Fresh[7387], Fresh[7386], Fresh[7385], Fresh[7384], Fresh[7383], Fresh[7382], Fresh[7381], Fresh[7380], Fresh[7379], Fresh[7378], Fresh[7377], Fresh[7376], Fresh[7375], Fresh[7374], Fresh[7373], Fresh[7372], Fresh[7371], Fresh[7370], Fresh[7369], Fresh[7368], Fresh[7367], Fresh[7366], Fresh[7365], Fresh[7364], Fresh[7363], Fresh[7362], Fresh[7361], Fresh[7360], Fresh[7359], Fresh[7358], Fresh[7357], Fresh[7356], Fresh[7355], Fresh[7354], Fresh[7353], Fresh[7352], Fresh[7351], Fresh[7350], Fresh[7349], Fresh[7348], Fresh[7347], Fresh[7346], Fresh[7345], Fresh[7344], Fresh[7343], Fresh[7342], Fresh[7341], Fresh[7340], Fresh[7339], Fresh[7338], Fresh[7337], Fresh[7336], Fresh[7335], Fresh[7334], Fresh[7333], Fresh[7332], Fresh[7331], Fresh[7330], Fresh[7329], Fresh[7328], Fresh[7327], Fresh[7326], Fresh[7325], Fresh[7324], Fresh[7323], Fresh[7322], Fresh[7321], Fresh[7320], Fresh[7319], Fresh[7318], Fresh[7317], Fresh[7316], Fresh[7315], Fresh[7314], Fresh[7313], Fresh[7312], Fresh[7311], Fresh[7310], Fresh[7309], Fresh[7308], Fresh[7307], Fresh[7306], Fresh[7305], Fresh[7304], Fresh[7303], Fresh[7302], Fresh[7301], Fresh[7300], Fresh[7299], Fresh[7298], Fresh[7297], Fresh[7296], Fresh[7295], Fresh[7294], Fresh[7293], Fresh[7292], Fresh[7291], Fresh[7290], Fresh[7289], Fresh[7288], Fresh[7287], Fresh[7286], Fresh[7285], Fresh[7284], Fresh[7283], Fresh[7282], Fresh[7281], Fresh[7280], Fresh[7279], Fresh[7278], Fresh[7277], Fresh[7276], Fresh[7275], Fresh[7274], Fresh[7273], Fresh[7272], Fresh[7271], Fresh[7270], Fresh[7269], Fresh[7268], Fresh[7267], Fresh[7266], Fresh[7265], Fresh[7264], Fresh[7263], Fresh[7262], Fresh[7261], Fresh[7260], Fresh[7259], Fresh[7258], Fresh[7257], Fresh[7256], Fresh[7255], Fresh[7254], Fresh[7253], Fresh[7252], Fresh[7251], Fresh[7250], Fresh[7249], Fresh[7248], Fresh[7247], Fresh[7246], Fresh[7245], Fresh[7244], Fresh[7243], Fresh[7242], Fresh[7241], Fresh[7240], Fresh[7239], Fresh[7238], Fresh[7237], Fresh[7236], Fresh[7235], Fresh[7234], Fresh[7233], Fresh[7232], Fresh[7231], Fresh[7230], Fresh[7229], Fresh[7228], Fresh[7227], Fresh[7226], Fresh[7225], Fresh[7224], Fresh[7223], Fresh[7222], Fresh[7221], Fresh[7220], Fresh[7219], Fresh[7218], Fresh[7217], Fresh[7216], Fresh[7215], Fresh[7214], Fresh[7213], Fresh[7212], Fresh[7211], Fresh[7210], Fresh[7209], Fresh[7208], Fresh[7207], Fresh[7206], Fresh[7205], Fresh[7204], Fresh[7203], Fresh[7202], Fresh[7201], Fresh[7200], Fresh[7199], Fresh[7198], Fresh[7197], Fresh[7196], Fresh[7195], Fresh[7194], Fresh[7193], Fresh[7192], Fresh[7191], Fresh[7190], Fresh[7189], Fresh[7188], Fresh[7187], Fresh[7186], Fresh[7185], Fresh[7184], Fresh[7183], Fresh[7182], Fresh[7181], Fresh[7180], Fresh[7179], Fresh[7178], Fresh[7177], Fresh[7176], Fresh[7175], Fresh[7174], Fresh[7173], Fresh[7172], Fresh[7171], Fresh[7170], Fresh[7169], Fresh[7168], Fresh[7167], Fresh[7166], Fresh[7165], Fresh[7164], Fresh[7163], Fresh[7162], Fresh[7161], Fresh[7160], Fresh[7159], Fresh[7158], Fresh[7157], Fresh[7156], Fresh[7155], Fresh[7154], Fresh[7153], Fresh[7152], Fresh[7151], Fresh[7150], Fresh[7149], Fresh[7148], Fresh[7147], Fresh[7146], Fresh[7145], Fresh[7144], Fresh[7143], Fresh[7142], Fresh[7141], Fresh[7140], Fresh[7139], Fresh[7138], Fresh[7137], Fresh[7136], Fresh[7135], Fresh[7134], Fresh[7133], Fresh[7132], Fresh[7131], Fresh[7130], Fresh[7129], Fresh[7128], Fresh[7127], Fresh[7126], Fresh[7125], Fresh[7124], Fresh[7123], Fresh[7122], Fresh[7121], Fresh[7120], Fresh[7119], Fresh[7118], Fresh[7117], Fresh[7116], Fresh[7115], Fresh[7114], Fresh[7113], Fresh[7112], Fresh[7111], Fresh[7110], Fresh[7109], Fresh[7108], Fresh[7107], Fresh[7106], Fresh[7105], Fresh[7104], Fresh[7103], Fresh[7102], Fresh[7101], Fresh[7100], Fresh[7099], Fresh[7098], Fresh[7097], Fresh[7096], Fresh[7095], Fresh[7094], Fresh[7093], Fresh[7092], Fresh[7091], Fresh[7090], Fresh[7089], Fresh[7088], Fresh[7087], Fresh[7086], Fresh[7085], Fresh[7084], Fresh[7083], Fresh[7082], Fresh[7081], Fresh[7080], Fresh[7079], Fresh[7078], Fresh[7077], Fresh[7076], Fresh[7075], Fresh[7074], Fresh[7073], Fresh[7072], Fresh[7071], Fresh[7070], Fresh[7069], Fresh[7068], Fresh[7067], Fresh[7066], Fresh[7065], Fresh[7064], Fresh[7063], Fresh[7062], Fresh[7061], Fresh[7060], Fresh[7059], Fresh[7058], Fresh[7057], Fresh[7056], Fresh[7055], Fresh[7054], Fresh[7053], Fresh[7052], Fresh[7051], Fresh[7050], Fresh[7049], Fresh[7048], Fresh[7047], Fresh[7046], Fresh[7045], Fresh[7044], Fresh[7043], Fresh[7042], Fresh[7041], Fresh[7040], Fresh[7039], Fresh[7038], Fresh[7037], Fresh[7036], Fresh[7035], Fresh[7034], Fresh[7033], Fresh[7032], Fresh[7031], Fresh[7030], Fresh[7029], Fresh[7028], Fresh[7027], Fresh[7026], Fresh[7025], Fresh[7024], Fresh[7023], Fresh[7022], Fresh[7021], Fresh[7020], Fresh[7019], Fresh[7018], Fresh[7017], Fresh[7016], Fresh[7015], Fresh[7014], Fresh[7013], Fresh[7012], Fresh[7011], Fresh[7010], Fresh[7009], Fresh[7008], Fresh[7007], Fresh[7006], Fresh[7005], Fresh[7004], Fresh[7003], Fresh[7002], Fresh[7001], Fresh[7000], Fresh[6999], Fresh[6998], Fresh[6997], Fresh[6996], Fresh[6995], Fresh[6994], Fresh[6993], Fresh[6992], Fresh[6991], Fresh[6990], Fresh[6989], Fresh[6988], Fresh[6987], Fresh[6986], Fresh[6985], Fresh[6984], Fresh[6983], Fresh[6982], Fresh[6981], Fresh[6980], Fresh[6979], Fresh[6978], Fresh[6977], Fresh[6976], Fresh[6975], Fresh[6974], Fresh[6973], Fresh[6972], Fresh[6971], Fresh[6970], Fresh[6969], Fresh[6968], Fresh[6967], Fresh[6966], Fresh[6965], Fresh[6964], Fresh[6963], Fresh[6962], Fresh[6961], Fresh[6960], Fresh[6959], Fresh[6958], Fresh[6957], Fresh[6956], Fresh[6955], Fresh[6954], Fresh[6953], Fresh[6952], Fresh[6951], Fresh[6950], Fresh[6949], Fresh[6948], Fresh[6947], Fresh[6946], Fresh[6945], Fresh[6944], Fresh[6943], Fresh[6942], Fresh[6941], Fresh[6940], Fresh[6939], Fresh[6938], Fresh[6937], Fresh[6936], Fresh[6935], Fresh[6934], Fresh[6933], Fresh[6932], Fresh[6931], Fresh[6930], Fresh[6929], Fresh[6928], Fresh[6927], Fresh[6926], Fresh[6925], Fresh[6924], Fresh[6923], Fresh[6922], Fresh[6921], Fresh[6920], Fresh[6919], Fresh[6918], Fresh[6917], Fresh[6916], Fresh[6915], Fresh[6914], Fresh[6913], Fresh[6912], Fresh[6911], Fresh[6910], Fresh[6909], Fresh[6908], Fresh[6907], Fresh[6906], Fresh[6905], Fresh[6904], Fresh[6903], Fresh[6902], Fresh[6901], Fresh[6900], Fresh[6899], Fresh[6898], Fresh[6897], Fresh[6896], Fresh[6895], Fresh[6894], Fresh[6893], Fresh[6892], Fresh[6891], Fresh[6890], Fresh[6889], Fresh[6888], Fresh[6887], Fresh[6886], Fresh[6885], Fresh[6884], Fresh[6883], Fresh[6882], Fresh[6881], Fresh[6880], Fresh[6879], Fresh[6878], Fresh[6877], Fresh[6876], Fresh[6875], Fresh[6874], Fresh[6873], Fresh[6872], Fresh[6871], Fresh[6870], Fresh[6869], Fresh[6868], Fresh[6867], Fresh[6866], Fresh[6865], Fresh[6864], Fresh[6863], Fresh[6862], Fresh[6861], Fresh[6860], Fresh[6859], Fresh[6858], Fresh[6857], Fresh[6856], Fresh[6855], Fresh[6854], Fresh[6853], Fresh[6852], Fresh[6851], Fresh[6850], Fresh[6849], Fresh[6848], Fresh[6847], Fresh[6846], Fresh[6845], Fresh[6844], Fresh[6843], Fresh[6842], Fresh[6841], Fresh[6840], Fresh[6839], Fresh[6838], Fresh[6837], Fresh[6836], Fresh[6835], Fresh[6834], Fresh[6833], Fresh[6832], Fresh[6831], Fresh[6830], Fresh[6829], Fresh[6828], Fresh[6827], Fresh[6826], Fresh[6825], Fresh[6824], Fresh[6823], Fresh[6822], Fresh[6821], Fresh[6820], Fresh[6819], Fresh[6818], Fresh[6817], Fresh[6816], Fresh[6815], Fresh[6814], Fresh[6813], Fresh[6812], Fresh[6811], Fresh[6810], Fresh[6809], Fresh[6808], Fresh[6807], Fresh[6806], Fresh[6805], Fresh[6804], Fresh[6803], Fresh[6802], Fresh[6801], Fresh[6800], Fresh[6799], Fresh[6798], Fresh[6797], Fresh[6796], Fresh[6795], Fresh[6794], Fresh[6793], Fresh[6792], Fresh[6791], Fresh[6790], Fresh[6789], Fresh[6788], Fresh[6787], Fresh[6786], Fresh[6785], Fresh[6784], Fresh[6783], Fresh[6782], Fresh[6781], Fresh[6780], Fresh[6779], Fresh[6778], Fresh[6777], Fresh[6776], Fresh[6775], Fresh[6774], Fresh[6773], Fresh[6772], Fresh[6771], Fresh[6770], Fresh[6769], Fresh[6768], Fresh[6767], Fresh[6766], Fresh[6765], Fresh[6764], Fresh[6763], Fresh[6762], Fresh[6761], Fresh[6760], Fresh[6759], Fresh[6758], Fresh[6757], Fresh[6756], Fresh[6755], Fresh[6754], Fresh[6753], Fresh[6752], Fresh[6751], Fresh[6750], Fresh[6749], Fresh[6748], Fresh[6747], Fresh[6746], Fresh[6745], Fresh[6744], Fresh[6743], Fresh[6742], Fresh[6741], Fresh[6740], Fresh[6739], Fresh[6738], Fresh[6737], Fresh[6736], Fresh[6735], Fresh[6734], Fresh[6733], Fresh[6732], Fresh[6731], Fresh[6730], Fresh[6729], Fresh[6728], Fresh[6727], Fresh[6726], Fresh[6725], Fresh[6724], Fresh[6723], Fresh[6722], Fresh[6721], Fresh[6720], Fresh[6719], Fresh[6718], Fresh[6717], Fresh[6716], Fresh[6715], Fresh[6714], Fresh[6713], Fresh[6712], Fresh[6711], Fresh[6710], Fresh[6709], Fresh[6708], Fresh[6707], Fresh[6706], Fresh[6705], Fresh[6704], Fresh[6703], Fresh[6702], Fresh[6701], Fresh[6700], Fresh[6699], Fresh[6698], Fresh[6697], Fresh[6696], Fresh[6695], Fresh[6694], Fresh[6693], Fresh[6692], Fresh[6691], Fresh[6690], Fresh[6689], Fresh[6688], Fresh[6687], Fresh[6686], Fresh[6685], Fresh[6684], Fresh[6683], Fresh[6682], Fresh[6681], Fresh[6680], Fresh[6679], Fresh[6678], Fresh[6677], Fresh[6676], Fresh[6675], Fresh[6674], Fresh[6673], Fresh[6672], Fresh[6671], Fresh[6670], Fresh[6669], Fresh[6668], Fresh[6667], Fresh[6666], Fresh[6665], Fresh[6664], Fresh[6663], Fresh[6662], Fresh[6661], Fresh[6660], Fresh[6659], Fresh[6658], Fresh[6657], Fresh[6656], Fresh[6655], Fresh[6654], Fresh[6653], Fresh[6652], Fresh[6651], Fresh[6650], Fresh[6649], Fresh[6648], Fresh[6647], Fresh[6646], Fresh[6645], Fresh[6644], Fresh[6643], Fresh[6642], Fresh[6641], Fresh[6640], Fresh[6639], Fresh[6638], Fresh[6637], Fresh[6636], Fresh[6635], Fresh[6634], Fresh[6633], Fresh[6632], Fresh[6631], Fresh[6630], Fresh[6629], Fresh[6628], Fresh[6627], Fresh[6626], Fresh[6625], Fresh[6624], Fresh[6623], Fresh[6622], Fresh[6621], Fresh[6620], Fresh[6619], Fresh[6618], Fresh[6617], Fresh[6616], Fresh[6615], Fresh[6614], Fresh[6613], Fresh[6612], Fresh[6611], Fresh[6610], Fresh[6609], Fresh[6608], Fresh[6607], Fresh[6606], Fresh[6605], Fresh[6604], Fresh[6603], Fresh[6602], Fresh[6601], Fresh[6600], Fresh[6599], Fresh[6598], Fresh[6597], Fresh[6596], Fresh[6595], Fresh[6594], Fresh[6593], Fresh[6592], Fresh[6591], Fresh[6590], Fresh[6589], Fresh[6588], Fresh[6587], Fresh[6586], Fresh[6585], Fresh[6584], Fresh[6583], Fresh[6582], Fresh[6581], Fresh[6580], Fresh[6579], Fresh[6578], Fresh[6577], Fresh[6576], Fresh[6575], Fresh[6574], Fresh[6573], Fresh[6572], Fresh[6571], Fresh[6570], Fresh[6569], Fresh[6568], Fresh[6567], Fresh[6566], Fresh[6565], Fresh[6564], Fresh[6563], Fresh[6562], Fresh[6561], Fresh[6560], Fresh[6559], Fresh[6558], Fresh[6557], Fresh[6556], Fresh[6555], Fresh[6554], Fresh[6553], Fresh[6552], Fresh[6551], Fresh[6550], Fresh[6549], Fresh[6548], Fresh[6547], Fresh[6546], Fresh[6545], Fresh[6544], Fresh[6543], Fresh[6542], Fresh[6541], Fresh[6540], Fresh[6539], Fresh[6538], Fresh[6537], Fresh[6536], Fresh[6535], Fresh[6534], Fresh[6533], Fresh[6532], Fresh[6531], Fresh[6530], Fresh[6529], Fresh[6528], Fresh[6527], Fresh[6526], Fresh[6525], Fresh[6524], Fresh[6523], Fresh[6522], Fresh[6521], Fresh[6520], Fresh[6519], Fresh[6518], Fresh[6517], Fresh[6516], Fresh[6515], Fresh[6514], Fresh[6513], Fresh[6512], Fresh[6511], Fresh[6510], Fresh[6509], Fresh[6508], Fresh[6507], Fresh[6506], Fresh[6505], Fresh[6504], Fresh[6503], Fresh[6502], Fresh[6501], Fresh[6500], Fresh[6499], Fresh[6498], Fresh[6497], Fresh[6496], Fresh[6495], Fresh[6494], Fresh[6493], Fresh[6492], Fresh[6491], Fresh[6490], Fresh[6489], Fresh[6488], Fresh[6487], Fresh[6486], Fresh[6485], Fresh[6484], Fresh[6483], Fresh[6482], Fresh[6481], Fresh[6480], Fresh[6479], Fresh[6478], Fresh[6477], Fresh[6476], Fresh[6475], Fresh[6474], Fresh[6473], Fresh[6472], Fresh[6471], Fresh[6470], Fresh[6469], Fresh[6468], Fresh[6467], Fresh[6466], Fresh[6465], Fresh[6464], Fresh[6463], Fresh[6462], Fresh[6461], Fresh[6460], Fresh[6459], Fresh[6458], Fresh[6457], Fresh[6456], Fresh[6455], Fresh[6454], Fresh[6453], Fresh[6452], Fresh[6451], Fresh[6450], Fresh[6449], Fresh[6448], Fresh[6447], Fresh[6446], Fresh[6445], Fresh[6444], Fresh[6443], Fresh[6442], Fresh[6441], Fresh[6440], Fresh[6439], Fresh[6438], Fresh[6437], Fresh[6436], Fresh[6435], Fresh[6434], Fresh[6433], Fresh[6432], Fresh[6431], Fresh[6430], Fresh[6429], Fresh[6428], Fresh[6427], Fresh[6426], Fresh[6425], Fresh[6424], Fresh[6423], Fresh[6422], Fresh[6421], Fresh[6420], Fresh[6419], Fresh[6418], Fresh[6417], Fresh[6416], Fresh[6415], Fresh[6414], Fresh[6413], Fresh[6412], Fresh[6411], Fresh[6410], Fresh[6409], Fresh[6408], Fresh[6407], Fresh[6406], Fresh[6405], Fresh[6404], Fresh[6403], Fresh[6402], Fresh[6401], Fresh[6400], Fresh[6399], Fresh[6398], Fresh[6397], Fresh[6396], Fresh[6395], Fresh[6394], Fresh[6393], Fresh[6392], Fresh[6391], Fresh[6390], Fresh[6389], Fresh[6388], Fresh[6387], Fresh[6386], Fresh[6385], Fresh[6384], Fresh[6383], Fresh[6382], Fresh[6381], Fresh[6380], Fresh[6379], Fresh[6378], Fresh[6377], Fresh[6376], Fresh[6375], Fresh[6374], Fresh[6373], Fresh[6372], Fresh[6371], Fresh[6370], Fresh[6369], Fresh[6368], Fresh[6367], Fresh[6366], Fresh[6365], Fresh[6364], Fresh[6363], Fresh[6362], Fresh[6361], Fresh[6360], Fresh[6359], Fresh[6358], Fresh[6357], Fresh[6356], Fresh[6355], Fresh[6354], Fresh[6353], Fresh[6352], Fresh[6351], Fresh[6350], Fresh[6349], Fresh[6348], Fresh[6347], Fresh[6346], Fresh[6345], Fresh[6344], Fresh[6343], Fresh[6342], Fresh[6341], Fresh[6340], Fresh[6339], Fresh[6338], Fresh[6337], Fresh[6336], Fresh[6335], Fresh[6334], Fresh[6333], Fresh[6332], Fresh[6331], Fresh[6330], Fresh[6329], Fresh[6328], Fresh[6327], Fresh[6326], Fresh[6325], Fresh[6324], Fresh[6323], Fresh[6322], Fresh[6321], Fresh[6320], Fresh[6319], Fresh[6318], Fresh[6317], Fresh[6316], Fresh[6315], Fresh[6314], Fresh[6313], Fresh[6312], Fresh[6311], Fresh[6310], Fresh[6309], Fresh[6308], Fresh[6307], Fresh[6306], Fresh[6305], Fresh[6304], Fresh[6303], Fresh[6302], Fresh[6301], Fresh[6300], Fresh[6299], Fresh[6298], Fresh[6297], Fresh[6296], Fresh[6295], Fresh[6294], Fresh[6293], Fresh[6292], Fresh[6291], Fresh[6290], Fresh[6289], Fresh[6288], Fresh[6287], Fresh[6286], Fresh[6285], Fresh[6284], Fresh[6283], Fresh[6282], Fresh[6281], Fresh[6280], Fresh[6279], Fresh[6278], Fresh[6277], Fresh[6276], Fresh[6275], Fresh[6274], Fresh[6273], Fresh[6272], Fresh[6271], Fresh[6270], Fresh[6269], Fresh[6268], Fresh[6267], Fresh[6266], Fresh[6265], Fresh[6264], Fresh[6263], Fresh[6262], Fresh[6261], Fresh[6260], Fresh[6259], Fresh[6258], Fresh[6257], Fresh[6256], Fresh[6255], Fresh[6254], Fresh[6253], Fresh[6252], Fresh[6251], Fresh[6250], Fresh[6249], Fresh[6248], Fresh[6247], Fresh[6246], Fresh[6245], Fresh[6244], Fresh[6243], Fresh[6242], Fresh[6241], Fresh[6240], Fresh[6239], Fresh[6238], Fresh[6237], Fresh[6236], Fresh[6235], Fresh[6234], Fresh[6233], Fresh[6232], Fresh[6231], Fresh[6230], Fresh[6229], Fresh[6228], Fresh[6227], Fresh[6226], Fresh[6225], Fresh[6224], Fresh[6223], Fresh[6222], Fresh[6221], Fresh[6220], Fresh[6219], Fresh[6218], Fresh[6217], Fresh[6216], Fresh[6215], Fresh[6214], Fresh[6213], Fresh[6212], Fresh[6211], Fresh[6210], Fresh[6209], Fresh[6208], Fresh[6207], Fresh[6206], Fresh[6205], Fresh[6204], Fresh[6203], Fresh[6202], Fresh[6201], Fresh[6200], Fresh[6199], Fresh[6198], Fresh[6197], Fresh[6196], Fresh[6195], Fresh[6194], Fresh[6193], Fresh[6192], Fresh[6191], Fresh[6190], Fresh[6189], Fresh[6188], Fresh[6187], Fresh[6186], Fresh[6185], Fresh[6184], Fresh[6183], Fresh[6182], Fresh[6181], Fresh[6180], Fresh[6179], Fresh[6178], Fresh[6177], Fresh[6176], Fresh[6175], Fresh[6174], Fresh[6173], Fresh[6172], Fresh[6171], Fresh[6170], Fresh[6169], Fresh[6168], Fresh[6167], Fresh[6166], Fresh[6165], Fresh[6164], Fresh[6163], Fresh[6162], Fresh[6161], Fresh[6160], Fresh[6159], Fresh[6158], Fresh[6157], Fresh[6156], Fresh[6155], Fresh[6154], Fresh[6153], Fresh[6152], Fresh[6151], Fresh[6150], Fresh[6149], Fresh[6148], Fresh[6147], Fresh[6146], Fresh[6145], Fresh[6144], Fresh[6143], Fresh[6142], Fresh[6141], Fresh[6140], Fresh[6139], Fresh[6138], Fresh[6137], Fresh[6136], Fresh[6135], Fresh[6134], Fresh[6133], Fresh[6132], Fresh[6131], Fresh[6130], Fresh[6129], Fresh[6128], Fresh[6127], Fresh[6126], Fresh[6125], Fresh[6124], Fresh[6123], Fresh[6122], Fresh[6121], Fresh[6120], Fresh[6119], Fresh[6118], Fresh[6117], Fresh[6116], Fresh[6115], Fresh[6114], Fresh[6113], Fresh[6112], Fresh[6111], Fresh[6110], Fresh[6109], Fresh[6108], Fresh[6107], Fresh[6106], Fresh[6105], Fresh[6104], Fresh[6103], Fresh[6102], Fresh[6101], Fresh[6100], Fresh[6099], Fresh[6098], Fresh[6097], Fresh[6096], Fresh[6095], Fresh[6094], Fresh[6093], Fresh[6092], Fresh[6091], Fresh[6090], Fresh[6089], Fresh[6088], Fresh[6087], Fresh[6086], Fresh[6085], Fresh[6084], Fresh[6083], Fresh[6082], Fresh[6081], Fresh[6080], Fresh[6079], Fresh[6078], Fresh[6077], Fresh[6076], Fresh[6075], Fresh[6074], Fresh[6073], Fresh[6072], Fresh[6071], Fresh[6070], Fresh[6069], Fresh[6068], Fresh[6067], Fresh[6066], Fresh[6065], Fresh[6064], Fresh[6063], Fresh[6062], Fresh[6061], Fresh[6060], Fresh[6059], Fresh[6058], Fresh[6057], Fresh[6056], Fresh[6055], Fresh[6054], Fresh[6053], Fresh[6052], Fresh[6051], Fresh[6050], Fresh[6049], Fresh[6048], Fresh[6047], Fresh[6046], Fresh[6045], Fresh[6044], Fresh[6043], Fresh[6042], Fresh[6041], Fresh[6040], Fresh[6039], Fresh[6038], Fresh[6037], Fresh[6036], Fresh[6035], Fresh[6034], Fresh[6033], Fresh[6032], Fresh[6031], Fresh[6030], Fresh[6029], Fresh[6028], Fresh[6027], Fresh[6026], Fresh[6025], Fresh[6024], Fresh[6023], Fresh[6022], Fresh[6021], Fresh[6020], Fresh[6019], Fresh[6018], Fresh[6017], Fresh[6016], Fresh[6015], Fresh[6014], Fresh[6013], Fresh[6012], Fresh[6011], Fresh[6010], Fresh[6009], Fresh[6008], Fresh[6007], Fresh[6006], Fresh[6005], Fresh[6004], Fresh[6003], Fresh[6002], Fresh[6001], Fresh[6000], Fresh[5999], Fresh[5998], Fresh[5997], Fresh[5996], Fresh[5995], Fresh[5994], Fresh[5993], Fresh[5992], Fresh[5991], Fresh[5990], Fresh[5989], Fresh[5988], Fresh[5987], Fresh[5986], Fresh[5985], Fresh[5984], Fresh[5983], Fresh[5982], Fresh[5981], Fresh[5980], Fresh[5979], Fresh[5978], Fresh[5977], Fresh[5976], Fresh[5975], Fresh[5974], Fresh[5973], Fresh[5972], Fresh[5971], Fresh[5970], Fresh[5969], Fresh[5968], Fresh[5967], Fresh[5966], Fresh[5965], Fresh[5964], Fresh[5963], Fresh[5962], Fresh[5961], Fresh[5960], Fresh[5959], Fresh[5958], Fresh[5957], Fresh[5956], Fresh[5955], Fresh[5954], Fresh[5953], Fresh[5952], Fresh[5951], Fresh[5950], Fresh[5949], Fresh[5948], Fresh[5947], Fresh[5946], Fresh[5945], Fresh[5944], Fresh[5943], Fresh[5942], Fresh[5941], Fresh[5940], Fresh[5939], Fresh[5938], Fresh[5937], Fresh[5936], Fresh[5935], Fresh[5934], Fresh[5933], Fresh[5932], Fresh[5931], Fresh[5930], Fresh[5929], Fresh[5928], Fresh[5927], Fresh[5926], Fresh[5925], Fresh[5924], Fresh[5923], Fresh[5922], Fresh[5921], Fresh[5920], Fresh[5919], Fresh[5918], Fresh[5917], Fresh[5916], Fresh[5915], Fresh[5914], Fresh[5913], Fresh[5912], Fresh[5911], Fresh[5910], Fresh[5909], Fresh[5908], Fresh[5907], Fresh[5906], Fresh[5905], Fresh[5904], Fresh[5903], Fresh[5902], Fresh[5901], Fresh[5900], Fresh[5899], Fresh[5898], Fresh[5897], Fresh[5896], Fresh[5895], Fresh[5894], Fresh[5893], Fresh[5892], Fresh[5891], Fresh[5890], Fresh[5889], Fresh[5888], Fresh[5887], Fresh[5886], Fresh[5885], Fresh[5884], Fresh[5883], Fresh[5882], Fresh[5881], Fresh[5880], Fresh[5879], Fresh[5878], Fresh[5877], Fresh[5876], Fresh[5875], Fresh[5874], Fresh[5873], Fresh[5872], Fresh[5871], Fresh[5870], Fresh[5869], Fresh[5868], Fresh[5867], Fresh[5866], Fresh[5865], Fresh[5864], Fresh[5863], Fresh[5862], Fresh[5861], Fresh[5860], Fresh[5859], Fresh[5858], Fresh[5857], Fresh[5856], Fresh[5855], Fresh[5854], Fresh[5853], Fresh[5852], Fresh[5851], Fresh[5850], Fresh[5849], Fresh[5848], Fresh[5847], Fresh[5846], Fresh[5845], Fresh[5844], Fresh[5843], Fresh[5842], Fresh[5841], Fresh[5840], Fresh[5839], Fresh[5838], Fresh[5837], Fresh[5836], Fresh[5835], Fresh[5834], Fresh[5833], Fresh[5832], Fresh[5831], Fresh[5830], Fresh[5829], Fresh[5828], Fresh[5827], Fresh[5826], Fresh[5825], Fresh[5824], Fresh[5823], Fresh[5822], Fresh[5821], Fresh[5820], Fresh[5819], Fresh[5818], Fresh[5817], Fresh[5816], Fresh[5815], Fresh[5814], Fresh[5813], Fresh[5812], Fresh[5811], Fresh[5810], Fresh[5809], Fresh[5808], Fresh[5807], Fresh[5806], Fresh[5805], Fresh[5804], Fresh[5803], Fresh[5802], Fresh[5801], Fresh[5800], Fresh[5799], Fresh[5798], Fresh[5797], Fresh[5796], Fresh[5795], Fresh[5794], Fresh[5793], Fresh[5792], Fresh[5791], Fresh[5790], Fresh[5789], Fresh[5788], Fresh[5787], Fresh[5786], Fresh[5785], Fresh[5784], Fresh[5783], Fresh[5782], Fresh[5781], Fresh[5780], Fresh[5779], Fresh[5778], Fresh[5777], Fresh[5776], Fresh[5775], Fresh[5774], Fresh[5773], Fresh[5772], Fresh[5771], Fresh[5770], Fresh[5769], Fresh[5768], Fresh[5767], Fresh[5766], Fresh[5765], Fresh[5764], Fresh[5763], Fresh[5762], Fresh[5761], Fresh[5760], Fresh[5759], Fresh[5758], Fresh[5757], Fresh[5756], Fresh[5755], Fresh[5754], Fresh[5753], Fresh[5752], Fresh[5751], Fresh[5750], Fresh[5749], Fresh[5748], Fresh[5747], Fresh[5746], Fresh[5745], Fresh[5744], Fresh[5743], Fresh[5742], Fresh[5741], Fresh[5740], Fresh[5739], Fresh[5738], Fresh[5737], Fresh[5736], Fresh[5735], Fresh[5734], Fresh[5733], Fresh[5732], Fresh[5731], Fresh[5730], Fresh[5729], Fresh[5728], Fresh[5727], Fresh[5726], Fresh[5725], Fresh[5724], Fresh[5723], Fresh[5722], Fresh[5721], Fresh[5720], Fresh[5719], Fresh[5718], Fresh[5717], Fresh[5716], Fresh[5715], Fresh[5714], Fresh[5713], Fresh[5712], Fresh[5711], Fresh[5710], Fresh[5709], Fresh[5708], Fresh[5707], Fresh[5706], Fresh[5705], Fresh[5704], Fresh[5703], Fresh[5702], Fresh[5701], Fresh[5700], Fresh[5699], Fresh[5698], Fresh[5697], Fresh[5696], Fresh[5695], Fresh[5694], Fresh[5693], Fresh[5692], Fresh[5691], Fresh[5690], Fresh[5689], Fresh[5688], Fresh[5687], Fresh[5686], Fresh[5685], Fresh[5684], Fresh[5683], Fresh[5682], Fresh[5681], Fresh[5680], Fresh[5679], Fresh[5678], Fresh[5677], Fresh[5676], Fresh[5675], Fresh[5674], Fresh[5673], Fresh[5672], Fresh[5671], Fresh[5670], Fresh[5669], Fresh[5668], Fresh[5667], Fresh[5666], Fresh[5665], Fresh[5664], Fresh[5663], Fresh[5662], Fresh[5661], Fresh[5660], Fresh[5659], Fresh[5658], Fresh[5657], Fresh[5656], Fresh[5655], Fresh[5654], Fresh[5653], Fresh[5652], Fresh[5651], Fresh[5650], Fresh[5649], Fresh[5648], Fresh[5647], Fresh[5646], Fresh[5645], Fresh[5644], Fresh[5643], Fresh[5642], Fresh[5641], Fresh[5640], Fresh[5639], Fresh[5638], Fresh[5637], Fresh[5636], Fresh[5635], Fresh[5634], Fresh[5633], Fresh[5632], Fresh[5631], Fresh[5630], Fresh[5629], Fresh[5628], Fresh[5627], Fresh[5626], Fresh[5625], Fresh[5624], Fresh[5623], Fresh[5622], Fresh[5621], Fresh[5620], Fresh[5619], Fresh[5618], Fresh[5617], Fresh[5616], Fresh[5615], Fresh[5614], Fresh[5613], Fresh[5612], Fresh[5611], Fresh[5610], Fresh[5609], Fresh[5608], Fresh[5607], Fresh[5606], Fresh[5605], Fresh[5604], Fresh[5603], Fresh[5602], Fresh[5601], Fresh[5600], Fresh[5599], Fresh[5598], Fresh[5597], Fresh[5596], Fresh[5595], Fresh[5594], Fresh[5593], Fresh[5592], Fresh[5591], Fresh[5590], Fresh[5589], Fresh[5588], Fresh[5587], Fresh[5586], Fresh[5585], Fresh[5584], Fresh[5583], Fresh[5582], Fresh[5581], Fresh[5580], Fresh[5579], Fresh[5578], Fresh[5577], Fresh[5576], Fresh[5575], Fresh[5574], Fresh[5573], Fresh[5572], Fresh[5571], Fresh[5570], Fresh[5569], Fresh[5568], Fresh[5567], Fresh[5566], Fresh[5565], Fresh[5564], Fresh[5563], Fresh[5562], Fresh[5561], Fresh[5560], Fresh[5559], Fresh[5558], Fresh[5557], Fresh[5556], Fresh[5555], Fresh[5554], Fresh[5553], Fresh[5552], Fresh[5551], Fresh[5550], Fresh[5549], Fresh[5548], Fresh[5547], Fresh[5546], Fresh[5545], Fresh[5544], Fresh[5543], Fresh[5542], Fresh[5541], Fresh[5540], Fresh[5539], Fresh[5538], Fresh[5537], Fresh[5536], Fresh[5535], Fresh[5534], Fresh[5533], Fresh[5532], Fresh[5531], Fresh[5530], Fresh[5529], Fresh[5528], Fresh[5527], Fresh[5526], Fresh[5525], Fresh[5524], Fresh[5523], Fresh[5522], Fresh[5521], Fresh[5520], Fresh[5519], Fresh[5518], Fresh[5517], Fresh[5516], Fresh[5515], Fresh[5514], Fresh[5513], Fresh[5512], Fresh[5511], Fresh[5510], Fresh[5509], Fresh[5508], Fresh[5507], Fresh[5506], Fresh[5505], Fresh[5504], Fresh[5503], Fresh[5502], Fresh[5501], Fresh[5500], Fresh[5499], Fresh[5498], Fresh[5497], Fresh[5496], Fresh[5495], Fresh[5494], Fresh[5493], Fresh[5492], Fresh[5491], Fresh[5490], Fresh[5489], Fresh[5488], Fresh[5487], Fresh[5486], Fresh[5485], Fresh[5484], Fresh[5483], Fresh[5482], Fresh[5481], Fresh[5480], Fresh[5479], Fresh[5478], Fresh[5477], Fresh[5476], Fresh[5475], Fresh[5474], Fresh[5473], Fresh[5472], Fresh[5471], Fresh[5470], Fresh[5469], Fresh[5468], Fresh[5467], Fresh[5466], Fresh[5465], Fresh[5464], Fresh[5463], Fresh[5462], Fresh[5461], Fresh[5460], Fresh[5459], Fresh[5458], Fresh[5457], Fresh[5456], Fresh[5455], Fresh[5454], Fresh[5453], Fresh[5452], Fresh[5451], Fresh[5450], Fresh[5449], Fresh[5448], Fresh[5447], Fresh[5446], Fresh[5445], Fresh[5444], Fresh[5443], Fresh[5442], Fresh[5441], Fresh[5440], Fresh[5439], Fresh[5438], Fresh[5437], Fresh[5436], Fresh[5435], Fresh[5434], Fresh[5433], Fresh[5432], Fresh[5431], Fresh[5430], Fresh[5429], Fresh[5428], Fresh[5427], Fresh[5426], Fresh[5425], Fresh[5424], Fresh[5423], Fresh[5422], Fresh[5421], Fresh[5420], Fresh[5419], Fresh[5418], Fresh[5417], Fresh[5416], Fresh[5415], Fresh[5414], Fresh[5413], Fresh[5412], Fresh[5411], Fresh[5410], Fresh[5409], Fresh[5408], Fresh[5407], Fresh[5406], Fresh[5405], Fresh[5404], Fresh[5403], Fresh[5402], Fresh[5401], Fresh[5400], Fresh[5399], Fresh[5398], Fresh[5397], Fresh[5396], Fresh[5395], Fresh[5394], Fresh[5393], Fresh[5392], Fresh[5391], Fresh[5390], Fresh[5389], Fresh[5388], Fresh[5387], Fresh[5386], Fresh[5385], Fresh[5384], Fresh[5383], Fresh[5382], Fresh[5381], Fresh[5380], Fresh[5379], Fresh[5378], Fresh[5377], Fresh[5376], Fresh[5375], Fresh[5374], Fresh[5373], Fresh[5372], Fresh[5371], Fresh[5370], Fresh[5369], Fresh[5368], Fresh[5367], Fresh[5366], Fresh[5365], Fresh[5364], Fresh[5363], Fresh[5362], Fresh[5361], Fresh[5360], Fresh[5359], Fresh[5358], Fresh[5357], Fresh[5356], Fresh[5355], Fresh[5354], Fresh[5353], Fresh[5352], Fresh[5351], Fresh[5350], Fresh[5349], Fresh[5348], Fresh[5347], Fresh[5346], Fresh[5345], Fresh[5344], Fresh[5343], Fresh[5342], Fresh[5341], Fresh[5340], Fresh[5339], Fresh[5338], Fresh[5337], Fresh[5336], Fresh[5335], Fresh[5334], Fresh[5333], Fresh[5332], Fresh[5331], Fresh[5330], Fresh[5329], Fresh[5328], Fresh[5327], Fresh[5326], Fresh[5325], Fresh[5324], Fresh[5323], Fresh[5322], Fresh[5321], Fresh[5320], Fresh[5319], Fresh[5318], Fresh[5317], Fresh[5316], Fresh[5315], Fresh[5314], Fresh[5313], Fresh[5312], Fresh[5311], Fresh[5310], Fresh[5309], Fresh[5308], Fresh[5307], Fresh[5306], Fresh[5305], Fresh[5304], Fresh[5303], Fresh[5302], Fresh[5301], Fresh[5300], Fresh[5299], Fresh[5298], Fresh[5297], Fresh[5296], Fresh[5295], Fresh[5294], Fresh[5293], Fresh[5292], Fresh[5291], Fresh[5290], Fresh[5289], Fresh[5288], Fresh[5287], Fresh[5286], Fresh[5285], Fresh[5284], Fresh[5283], Fresh[5282], Fresh[5281], Fresh[5280], Fresh[5279], Fresh[5278], Fresh[5277], Fresh[5276], Fresh[5275], Fresh[5274], Fresh[5273], Fresh[5272], Fresh[5271], Fresh[5270], Fresh[5269], Fresh[5268], Fresh[5267], Fresh[5266], Fresh[5265], Fresh[5264], Fresh[5263], Fresh[5262], Fresh[5261], Fresh[5260], Fresh[5259], Fresh[5258], Fresh[5257], Fresh[5256], Fresh[5255], Fresh[5254], Fresh[5253], Fresh[5252], Fresh[5251], Fresh[5250], Fresh[5249], Fresh[5248], Fresh[5247], Fresh[5246], Fresh[5245], Fresh[5244], Fresh[5243], Fresh[5242], Fresh[5241], Fresh[5240], Fresh[5239], Fresh[5238], Fresh[5237], Fresh[5236], Fresh[5235], Fresh[5234], Fresh[5233], Fresh[5232], Fresh[5231], Fresh[5230], Fresh[5229], Fresh[5228], Fresh[5227], Fresh[5226], Fresh[5225], Fresh[5224], Fresh[5223], Fresh[5222], Fresh[5221], Fresh[5220], Fresh[5219], Fresh[5218], Fresh[5217], Fresh[5216], Fresh[5215], Fresh[5214], Fresh[5213], Fresh[5212], Fresh[5211], Fresh[5210], Fresh[5209], Fresh[5208], Fresh[5207], Fresh[5206], Fresh[5205], Fresh[5204], Fresh[5203], Fresh[5202], Fresh[5201], Fresh[5200], Fresh[5199], Fresh[5198], Fresh[5197], Fresh[5196], Fresh[5195], Fresh[5194], Fresh[5193], Fresh[5192], Fresh[5191], Fresh[5190], Fresh[5189], Fresh[5188], Fresh[5187], Fresh[5186], Fresh[5185], Fresh[5184], Fresh[5183], Fresh[5182], Fresh[5181], Fresh[5180], Fresh[5179], Fresh[5178], Fresh[5177], Fresh[5176], Fresh[5175], Fresh[5174], Fresh[5173], Fresh[5172], Fresh[5171], Fresh[5170], Fresh[5169], Fresh[5168], Fresh[5167], Fresh[5166], Fresh[5165], Fresh[5164], Fresh[5163], Fresh[5162], Fresh[5161], Fresh[5160], Fresh[5159], Fresh[5158], Fresh[5157], Fresh[5156], Fresh[5155], Fresh[5154], Fresh[5153], Fresh[5152], Fresh[5151], Fresh[5150], Fresh[5149], Fresh[5148], Fresh[5147], Fresh[5146], Fresh[5145], Fresh[5144], Fresh[5143], Fresh[5142], Fresh[5141], Fresh[5140], Fresh[5139], Fresh[5138], Fresh[5137], Fresh[5136], Fresh[5135], Fresh[5134], Fresh[5133], Fresh[5132], Fresh[5131], Fresh[5130], Fresh[5129], Fresh[5128], Fresh[5127], Fresh[5126], Fresh[5125], Fresh[5124], Fresh[5123], Fresh[5122], Fresh[5121], Fresh[5120], Fresh[5119], Fresh[5118], Fresh[5117], Fresh[5116], Fresh[5115], Fresh[5114], Fresh[5113], Fresh[5112], Fresh[5111], Fresh[5110], Fresh[5109], Fresh[5108], Fresh[5107], Fresh[5106], Fresh[5105], Fresh[5104], Fresh[5103], Fresh[5102], Fresh[5101], Fresh[5100], Fresh[5099], Fresh[5098], Fresh[5097], Fresh[5096], Fresh[5095], Fresh[5094], Fresh[5093], Fresh[5092], Fresh[5091], Fresh[5090], Fresh[5089], Fresh[5088], Fresh[5087], Fresh[5086], Fresh[5085], Fresh[5084], Fresh[5083], Fresh[5082], Fresh[5081], Fresh[5080], Fresh[5079], Fresh[5078], Fresh[5077], Fresh[5076], Fresh[5075], Fresh[5074], Fresh[5073], Fresh[5072], Fresh[5071], Fresh[5070], Fresh[5069], Fresh[5068], Fresh[5067], Fresh[5066], Fresh[5065], Fresh[5064], Fresh[5063], Fresh[5062], Fresh[5061], Fresh[5060], Fresh[5059], Fresh[5058], Fresh[5057], Fresh[5056], Fresh[5055], Fresh[5054], Fresh[5053], Fresh[5052], Fresh[5051], Fresh[5050], Fresh[5049], Fresh[5048], Fresh[5047], Fresh[5046], Fresh[5045], Fresh[5044], Fresh[5043], Fresh[5042], Fresh[5041], Fresh[5040], Fresh[5039], Fresh[5038], Fresh[5037], Fresh[5036], Fresh[5035], Fresh[5034], Fresh[5033], Fresh[5032], Fresh[5031], Fresh[5030], Fresh[5029], Fresh[5028], Fresh[5027], Fresh[5026], Fresh[5025], Fresh[5024], Fresh[5023], Fresh[5022], Fresh[5021], Fresh[5020], Fresh[5019], Fresh[5018], Fresh[5017], Fresh[5016], Fresh[5015], Fresh[5014], Fresh[5013], Fresh[5012], Fresh[5011], Fresh[5010], Fresh[5009], Fresh[5008], Fresh[5007], Fresh[5006], Fresh[5005], Fresh[5004], Fresh[5003], Fresh[5002], Fresh[5001], Fresh[5000], Fresh[4999], Fresh[4998], Fresh[4997], Fresh[4996], Fresh[4995], Fresh[4994], Fresh[4993], Fresh[4992], Fresh[4991], Fresh[4990], Fresh[4989], Fresh[4988], Fresh[4987], Fresh[4986], Fresh[4985], Fresh[4984], Fresh[4983], Fresh[4982], Fresh[4981], Fresh[4980], Fresh[4979], Fresh[4978], Fresh[4977], Fresh[4976], Fresh[4975], Fresh[4974], Fresh[4973], Fresh[4972], Fresh[4971], Fresh[4970], Fresh[4969], Fresh[4968], Fresh[4967], Fresh[4966], Fresh[4965], Fresh[4964], Fresh[4963], Fresh[4962], Fresh[4961], Fresh[4960], Fresh[4959], Fresh[4958], Fresh[4957], Fresh[4956], Fresh[4955], Fresh[4954], Fresh[4953], Fresh[4952], Fresh[4951], Fresh[4950], Fresh[4949], Fresh[4948], Fresh[4947], Fresh[4946], Fresh[4945], Fresh[4944], Fresh[4943], Fresh[4942], Fresh[4941], Fresh[4940], Fresh[4939], Fresh[4938], Fresh[4937], Fresh[4936], Fresh[4935], Fresh[4934], Fresh[4933], Fresh[4932], Fresh[4931], Fresh[4930], Fresh[4929], Fresh[4928], Fresh[4927], Fresh[4926], Fresh[4925], Fresh[4924], Fresh[4923], Fresh[4922], Fresh[4921], Fresh[4920], Fresh[4919], Fresh[4918], Fresh[4917], Fresh[4916], Fresh[4915], Fresh[4914], Fresh[4913], Fresh[4912], Fresh[4911], Fresh[4910], Fresh[4909], Fresh[4908], Fresh[4907], Fresh[4906], Fresh[4905], Fresh[4904], Fresh[4903], Fresh[4902], Fresh[4901], Fresh[4900], Fresh[4899], Fresh[4898], Fresh[4897], Fresh[4896], Fresh[4895], Fresh[4894], Fresh[4893], Fresh[4892], Fresh[4891], Fresh[4890], Fresh[4889], Fresh[4888], Fresh[4887], Fresh[4886], Fresh[4885], Fresh[4884], Fresh[4883], Fresh[4882], Fresh[4881], Fresh[4880], Fresh[4879], Fresh[4878], Fresh[4877], Fresh[4876], Fresh[4875], Fresh[4874], Fresh[4873], Fresh[4872], Fresh[4871], Fresh[4870], Fresh[4869], Fresh[4868], Fresh[4867], Fresh[4866], Fresh[4865], Fresh[4864], Fresh[4863], Fresh[4862], Fresh[4861], Fresh[4860], Fresh[4859], Fresh[4858], Fresh[4857], Fresh[4856], Fresh[4855], Fresh[4854], Fresh[4853], Fresh[4852], Fresh[4851], Fresh[4850], Fresh[4849], Fresh[4848], Fresh[4847], Fresh[4846], Fresh[4845], Fresh[4844], Fresh[4843], Fresh[4842], Fresh[4841], Fresh[4840], Fresh[4839], Fresh[4838], Fresh[4837], Fresh[4836], Fresh[4835], Fresh[4834], Fresh[4833], Fresh[4832], Fresh[4831], Fresh[4830], Fresh[4829], Fresh[4828], Fresh[4827], Fresh[4826], Fresh[4825], Fresh[4824], Fresh[4823], Fresh[4822], Fresh[4821], Fresh[4820], Fresh[4819], Fresh[4818], Fresh[4817], Fresh[4816], Fresh[4815], Fresh[4814], Fresh[4813], Fresh[4812], Fresh[4811], Fresh[4810], Fresh[4809], Fresh[4808], Fresh[4807], Fresh[4806], Fresh[4805], Fresh[4804], Fresh[4803], Fresh[4802], Fresh[4801], Fresh[4800], Fresh[4799], Fresh[4798], Fresh[4797], Fresh[4796], Fresh[4795], Fresh[4794], Fresh[4793], Fresh[4792], Fresh[4791], Fresh[4790], Fresh[4789], Fresh[4788], Fresh[4787], Fresh[4786], Fresh[4785], Fresh[4784], Fresh[4783], Fresh[4782], Fresh[4781], Fresh[4780], Fresh[4779], Fresh[4778], Fresh[4777], Fresh[4776], Fresh[4775], Fresh[4774], Fresh[4773], Fresh[4772], Fresh[4771], Fresh[4770], Fresh[4769], Fresh[4768], Fresh[4767], Fresh[4766], Fresh[4765], Fresh[4764], Fresh[4763], Fresh[4762], Fresh[4761], Fresh[4760], Fresh[4759], Fresh[4758], Fresh[4757], Fresh[4756], Fresh[4755], Fresh[4754], Fresh[4753], Fresh[4752], Fresh[4751], Fresh[4750], Fresh[4749], Fresh[4748], Fresh[4747], Fresh[4746], Fresh[4745], Fresh[4744], Fresh[4743], Fresh[4742], Fresh[4741], Fresh[4740], Fresh[4739], Fresh[4738], Fresh[4737], Fresh[4736], Fresh[4735], Fresh[4734], Fresh[4733], Fresh[4732], Fresh[4731], Fresh[4730], Fresh[4729], Fresh[4728], Fresh[4727], Fresh[4726], Fresh[4725], Fresh[4724], Fresh[4723], Fresh[4722], Fresh[4721], Fresh[4720], Fresh[4719], Fresh[4718], Fresh[4717], Fresh[4716], Fresh[4715], Fresh[4714], Fresh[4713], Fresh[4712], Fresh[4711], Fresh[4710], Fresh[4709], Fresh[4708], Fresh[4707], Fresh[4706], Fresh[4705], Fresh[4704], Fresh[4703], Fresh[4702], Fresh[4701], Fresh[4700], Fresh[4699], Fresh[4698], Fresh[4697], Fresh[4696], Fresh[4695], Fresh[4694], Fresh[4693], Fresh[4692], Fresh[4691], Fresh[4690], Fresh[4689], Fresh[4688], Fresh[4687], Fresh[4686], Fresh[4685], Fresh[4684], Fresh[4683], Fresh[4682], Fresh[4681], Fresh[4680], Fresh[4679], Fresh[4678], Fresh[4677], Fresh[4676], Fresh[4675], Fresh[4674], Fresh[4673], Fresh[4672], Fresh[4671], Fresh[4670], Fresh[4669], Fresh[4668], Fresh[4667], Fresh[4666], Fresh[4665], Fresh[4664], Fresh[4663], Fresh[4662], Fresh[4661], Fresh[4660], Fresh[4659], Fresh[4658], Fresh[4657], Fresh[4656], Fresh[4655], Fresh[4654], Fresh[4653], Fresh[4652], Fresh[4651], Fresh[4650], Fresh[4649], Fresh[4648], Fresh[4647], Fresh[4646], Fresh[4645], Fresh[4644], Fresh[4643], Fresh[4642], Fresh[4641], Fresh[4640], Fresh[4639], Fresh[4638], Fresh[4637], Fresh[4636], Fresh[4635], Fresh[4634], Fresh[4633], Fresh[4632], Fresh[4631], Fresh[4630], Fresh[4629], Fresh[4628], Fresh[4627], Fresh[4626], Fresh[4625], Fresh[4624], Fresh[4623], Fresh[4622], Fresh[4621], Fresh[4620], Fresh[4619], Fresh[4618], Fresh[4617], Fresh[4616], Fresh[4615], Fresh[4614], Fresh[4613], Fresh[4612], Fresh[4611], Fresh[4610], Fresh[4609], Fresh[4608], Fresh[4607], Fresh[4606], Fresh[4605], Fresh[4604], Fresh[4603], Fresh[4602], Fresh[4601], Fresh[4600], Fresh[4599], Fresh[4598], Fresh[4597], Fresh[4596], Fresh[4595], Fresh[4594], Fresh[4593], Fresh[4592], Fresh[4591], Fresh[4590], Fresh[4589], Fresh[4588], Fresh[4587], Fresh[4586], Fresh[4585], Fresh[4584], Fresh[4583], Fresh[4582], Fresh[4581], Fresh[4580], Fresh[4579], Fresh[4578], Fresh[4577], Fresh[4576], Fresh[4575], Fresh[4574], Fresh[4573], Fresh[4572], Fresh[4571], Fresh[4570], Fresh[4569], Fresh[4568], Fresh[4567], Fresh[4566], Fresh[4565], Fresh[4564], Fresh[4563], Fresh[4562], Fresh[4561], Fresh[4560], Fresh[4559], Fresh[4558], Fresh[4557], Fresh[4556], Fresh[4555], Fresh[4554], Fresh[4553], Fresh[4552], Fresh[4551], Fresh[4550], Fresh[4549], Fresh[4548], Fresh[4547], Fresh[4546], Fresh[4545], Fresh[4544], Fresh[4543], Fresh[4542], Fresh[4541], Fresh[4540], Fresh[4539], Fresh[4538], Fresh[4537], Fresh[4536], Fresh[4535], Fresh[4534], Fresh[4533], Fresh[4532], Fresh[4531], Fresh[4530], Fresh[4529], Fresh[4528], Fresh[4527], Fresh[4526], Fresh[4525], Fresh[4524], Fresh[4523], Fresh[4522], Fresh[4521], Fresh[4520], Fresh[4519], Fresh[4518], Fresh[4517], Fresh[4516], Fresh[4515], Fresh[4514], Fresh[4513], Fresh[4512], Fresh[4511], Fresh[4510], Fresh[4509], Fresh[4508], Fresh[4507], Fresh[4506], Fresh[4505], Fresh[4504], Fresh[4503], Fresh[4502], Fresh[4501], Fresh[4500], Fresh[4499], Fresh[4498], Fresh[4497], Fresh[4496], Fresh[4495], Fresh[4494], Fresh[4493], Fresh[4492], Fresh[4491], Fresh[4490], Fresh[4489], Fresh[4488], Fresh[4487], Fresh[4486], Fresh[4485], Fresh[4484], Fresh[4483], Fresh[4482], Fresh[4481], Fresh[4480], Fresh[4479], Fresh[4478], Fresh[4477], Fresh[4476], Fresh[4475], Fresh[4474], Fresh[4473], Fresh[4472], Fresh[4471], Fresh[4470], Fresh[4469], Fresh[4468], Fresh[4467], Fresh[4466], Fresh[4465], Fresh[4464], Fresh[4463], Fresh[4462], Fresh[4461], Fresh[4460], Fresh[4459], Fresh[4458], Fresh[4457], Fresh[4456], Fresh[4455], Fresh[4454], Fresh[4453], Fresh[4452], Fresh[4451], Fresh[4450], Fresh[4449], Fresh[4448], Fresh[4447], Fresh[4446], Fresh[4445], Fresh[4444], Fresh[4443], Fresh[4442], Fresh[4441], Fresh[4440], Fresh[4439], Fresh[4438], Fresh[4437], Fresh[4436], Fresh[4435], Fresh[4434], Fresh[4433], Fresh[4432], Fresh[4431], Fresh[4430], Fresh[4429], Fresh[4428], Fresh[4427], Fresh[4426], Fresh[4425], Fresh[4424], Fresh[4423], Fresh[4422], Fresh[4421], Fresh[4420], Fresh[4419], Fresh[4418], Fresh[4417], Fresh[4416], Fresh[4415], Fresh[4414], Fresh[4413], Fresh[4412], Fresh[4411], Fresh[4410], Fresh[4409], Fresh[4408], Fresh[4407], Fresh[4406], Fresh[4405], Fresh[4404], Fresh[4403], Fresh[4402], Fresh[4401], Fresh[4400], Fresh[4399], Fresh[4398], Fresh[4397], Fresh[4396], Fresh[4395], Fresh[4394], Fresh[4393], Fresh[4392], Fresh[4391], Fresh[4390], Fresh[4389], Fresh[4388], Fresh[4387], Fresh[4386], Fresh[4385], Fresh[4384], Fresh[4383], Fresh[4382], Fresh[4381], Fresh[4380], Fresh[4379], Fresh[4378], Fresh[4377], Fresh[4376], Fresh[4375], Fresh[4374], Fresh[4373], Fresh[4372], Fresh[4371], Fresh[4370], Fresh[4369], Fresh[4368], Fresh[4367], Fresh[4366], Fresh[4365], Fresh[4364], Fresh[4363], Fresh[4362], Fresh[4361], Fresh[4360], Fresh[4359], Fresh[4358], Fresh[4357], Fresh[4356], Fresh[4355], Fresh[4354], Fresh[4353], Fresh[4352], Fresh[4351], Fresh[4350], Fresh[4349], Fresh[4348], Fresh[4347], Fresh[4346], Fresh[4345], Fresh[4344], Fresh[4343], Fresh[4342], Fresh[4341], Fresh[4340], Fresh[4339], Fresh[4338], Fresh[4337], Fresh[4336], Fresh[4335], Fresh[4334], Fresh[4333], Fresh[4332], Fresh[4331], Fresh[4330], Fresh[4329], Fresh[4328], Fresh[4327], Fresh[4326], Fresh[4325], Fresh[4324], Fresh[4323], Fresh[4322], Fresh[4321], Fresh[4320], Fresh[4319], Fresh[4318], Fresh[4317], Fresh[4316], Fresh[4315], Fresh[4314], Fresh[4313], Fresh[4312], Fresh[4311], Fresh[4310], Fresh[4309], Fresh[4308], Fresh[4307], Fresh[4306], Fresh[4305], Fresh[4304], Fresh[4303], Fresh[4302], Fresh[4301], Fresh[4300], Fresh[4299], Fresh[4298], Fresh[4297], Fresh[4296], Fresh[4295], Fresh[4294], Fresh[4293], Fresh[4292], Fresh[4291], Fresh[4290], Fresh[4289], Fresh[4288], Fresh[4287], Fresh[4286], Fresh[4285], Fresh[4284], Fresh[4283], Fresh[4282], Fresh[4281], Fresh[4280], Fresh[4279], Fresh[4278], Fresh[4277], Fresh[4276], Fresh[4275], Fresh[4274], Fresh[4273], Fresh[4272], Fresh[4271], Fresh[4270], Fresh[4269], Fresh[4268], Fresh[4267], Fresh[4266], Fresh[4265], Fresh[4264], Fresh[4263], Fresh[4262], Fresh[4261], Fresh[4260], Fresh[4259], Fresh[4258], Fresh[4257], Fresh[4256], Fresh[4255], Fresh[4254], Fresh[4253], Fresh[4252], Fresh[4251], Fresh[4250], Fresh[4249], Fresh[4248], Fresh[4247], Fresh[4246], Fresh[4245], Fresh[4244], Fresh[4243], Fresh[4242], Fresh[4241], Fresh[4240], Fresh[4239], Fresh[4238], Fresh[4237], Fresh[4236], Fresh[4235], Fresh[4234], Fresh[4233], Fresh[4232], Fresh[4231], Fresh[4230], Fresh[4229], Fresh[4228], Fresh[4227], Fresh[4226], Fresh[4225], Fresh[4224], Fresh[4223], Fresh[4222], Fresh[4221], Fresh[4220], Fresh[4219], Fresh[4218], Fresh[4217], Fresh[4216], Fresh[4215], Fresh[4214], Fresh[4213], Fresh[4212], Fresh[4211], Fresh[4210], Fresh[4209], Fresh[4208], Fresh[4207], Fresh[4206], Fresh[4205], Fresh[4204], Fresh[4203], Fresh[4202], Fresh[4201], Fresh[4200], Fresh[4199], Fresh[4198], Fresh[4197], Fresh[4196], Fresh[4195], Fresh[4194], Fresh[4193], Fresh[4192], Fresh[4191], Fresh[4190], Fresh[4189], Fresh[4188], Fresh[4187], Fresh[4186], Fresh[4185], Fresh[4184], Fresh[4183], Fresh[4182], Fresh[4181], Fresh[4180], Fresh[4179], Fresh[4178], Fresh[4177], Fresh[4176], Fresh[4175], Fresh[4174], Fresh[4173], Fresh[4172], Fresh[4171], Fresh[4170], Fresh[4169], Fresh[4168], Fresh[4167], Fresh[4166], Fresh[4165], Fresh[4164], Fresh[4163], Fresh[4162], Fresh[4161], Fresh[4160], Fresh[4159], Fresh[4158], Fresh[4157], Fresh[4156], Fresh[4155], Fresh[4154], Fresh[4153], Fresh[4152], Fresh[4151], Fresh[4150], Fresh[4149], Fresh[4148], Fresh[4147], Fresh[4146], Fresh[4145], Fresh[4144], Fresh[4143], Fresh[4142], Fresh[4141], Fresh[4140], Fresh[4139], Fresh[4138], Fresh[4137], Fresh[4136], Fresh[4135], Fresh[4134], Fresh[4133], Fresh[4132], Fresh[4131], Fresh[4130], Fresh[4129], Fresh[4128], Fresh[4127], Fresh[4126], Fresh[4125], Fresh[4124], Fresh[4123], Fresh[4122], Fresh[4121], Fresh[4120], Fresh[4119], Fresh[4118], Fresh[4117], Fresh[4116], Fresh[4115], Fresh[4114], Fresh[4113], Fresh[4112], Fresh[4111], Fresh[4110], Fresh[4109], Fresh[4108], Fresh[4107], Fresh[4106], Fresh[4105], Fresh[4104], Fresh[4103], Fresh[4102], Fresh[4101], Fresh[4100], Fresh[4099], Fresh[4098], Fresh[4097], Fresh[4096], Fresh[4095], Fresh[4094], Fresh[4093], Fresh[4092], Fresh[4091], Fresh[4090], Fresh[4089], Fresh[4088], Fresh[4087], Fresh[4086], Fresh[4085], Fresh[4084], Fresh[4083], Fresh[4082], Fresh[4081], Fresh[4080], Fresh[4079], Fresh[4078], Fresh[4077], Fresh[4076], Fresh[4075], Fresh[4074], Fresh[4073], Fresh[4072], Fresh[4071], Fresh[4070], Fresh[4069], Fresh[4068], Fresh[4067], Fresh[4066], Fresh[4065], Fresh[4064], Fresh[4063], Fresh[4062], Fresh[4061], Fresh[4060], Fresh[4059], Fresh[4058], Fresh[4057], Fresh[4056], Fresh[4055], Fresh[4054], Fresh[4053], Fresh[4052], Fresh[4051], Fresh[4050], Fresh[4049], Fresh[4048], Fresh[4047], Fresh[4046], Fresh[4045], Fresh[4044], Fresh[4043], Fresh[4042], Fresh[4041], Fresh[4040], Fresh[4039], Fresh[4038], Fresh[4037], Fresh[4036], Fresh[4035], Fresh[4034], Fresh[4033], Fresh[4032], Fresh[4031], Fresh[4030], Fresh[4029], Fresh[4028], Fresh[4027], Fresh[4026], Fresh[4025], Fresh[4024], Fresh[4023], Fresh[4022], Fresh[4021], Fresh[4020], Fresh[4019], Fresh[4018], Fresh[4017], Fresh[4016], Fresh[4015], Fresh[4014], Fresh[4013], Fresh[4012], Fresh[4011], Fresh[4010], Fresh[4009], Fresh[4008], Fresh[4007], Fresh[4006], Fresh[4005], Fresh[4004], Fresh[4003], Fresh[4002], Fresh[4001], Fresh[4000], Fresh[3999], Fresh[3998], Fresh[3997], Fresh[3996], Fresh[3995], Fresh[3994], Fresh[3993], Fresh[3992], Fresh[3991], Fresh[3990], Fresh[3989], Fresh[3988], Fresh[3987], Fresh[3986], Fresh[3985], Fresh[3984], Fresh[3983], Fresh[3982], Fresh[3981], Fresh[3980], Fresh[3979], Fresh[3978], Fresh[3977], Fresh[3976], Fresh[3975], Fresh[3974], Fresh[3973], Fresh[3972], Fresh[3971], Fresh[3970], Fresh[3969], Fresh[3968], Fresh[3967], Fresh[3966], Fresh[3965], Fresh[3964], Fresh[3963], Fresh[3962], Fresh[3961], Fresh[3960], Fresh[3959], Fresh[3958], Fresh[3957], Fresh[3956], Fresh[3955], Fresh[3954], Fresh[3953], Fresh[3952], Fresh[3951], Fresh[3950], Fresh[3949], Fresh[3948], Fresh[3947], Fresh[3946], Fresh[3945], Fresh[3944], Fresh[3943], Fresh[3942], Fresh[3941], Fresh[3940], Fresh[3939], Fresh[3938], Fresh[3937], Fresh[3936], Fresh[3935], Fresh[3934], Fresh[3933], Fresh[3932], Fresh[3931], Fresh[3930], Fresh[3929], Fresh[3928], Fresh[3927], Fresh[3926], Fresh[3925], Fresh[3924], Fresh[3923], Fresh[3922], Fresh[3921], Fresh[3920], Fresh[3919], Fresh[3918], Fresh[3917], Fresh[3916], Fresh[3915], Fresh[3914], Fresh[3913], Fresh[3912], Fresh[3911], Fresh[3910], Fresh[3909], Fresh[3908], Fresh[3907], Fresh[3906], Fresh[3905], Fresh[3904], Fresh[3903], Fresh[3902], Fresh[3901], Fresh[3900], Fresh[3899], Fresh[3898], Fresh[3897], Fresh[3896], Fresh[3895], Fresh[3894], Fresh[3893], Fresh[3892], Fresh[3891], Fresh[3890], Fresh[3889], Fresh[3888], Fresh[3887], Fresh[3886], Fresh[3885], Fresh[3884], Fresh[3883], Fresh[3882], Fresh[3881], Fresh[3880], Fresh[3879], Fresh[3878], Fresh[3877], Fresh[3876], Fresh[3875], Fresh[3874], Fresh[3873], Fresh[3872], Fresh[3871], Fresh[3870], Fresh[3869], Fresh[3868], Fresh[3867], Fresh[3866], Fresh[3865], Fresh[3864], Fresh[3863], Fresh[3862], Fresh[3861], Fresh[3860], Fresh[3859], Fresh[3858], Fresh[3857], Fresh[3856], Fresh[3855], Fresh[3854], Fresh[3853], Fresh[3852], Fresh[3851], Fresh[3850], Fresh[3849], Fresh[3848], Fresh[3847], Fresh[3846], Fresh[3845], Fresh[3844], Fresh[3843], Fresh[3842], Fresh[3841], Fresh[3840], Fresh[3839], Fresh[3838], Fresh[3837], Fresh[3836], Fresh[3835], Fresh[3834], Fresh[3833], Fresh[3832], Fresh[3831], Fresh[3830], Fresh[3829], Fresh[3828], Fresh[3827], Fresh[3826], Fresh[3825], Fresh[3824], Fresh[3823], Fresh[3822], Fresh[3821], Fresh[3820], Fresh[3819], Fresh[3818], Fresh[3817], Fresh[3816], Fresh[3815], Fresh[3814], Fresh[3813], Fresh[3812], Fresh[3811], Fresh[3810], Fresh[3809], Fresh[3808], Fresh[3807], Fresh[3806], Fresh[3805], Fresh[3804], Fresh[3803], Fresh[3802], Fresh[3801], Fresh[3800], Fresh[3799], Fresh[3798], Fresh[3797], Fresh[3796], Fresh[3795], Fresh[3794], Fresh[3793], Fresh[3792], Fresh[3791], Fresh[3790], Fresh[3789], Fresh[3788], Fresh[3787], Fresh[3786], Fresh[3785], Fresh[3784], Fresh[3783], Fresh[3782], Fresh[3781], Fresh[3780], Fresh[3779], Fresh[3778], Fresh[3777], Fresh[3776], Fresh[3775], Fresh[3774], Fresh[3773], Fresh[3772], Fresh[3771], Fresh[3770], Fresh[3769], Fresh[3768], Fresh[3767], Fresh[3766], Fresh[3765], Fresh[3764], Fresh[3763], Fresh[3762], Fresh[3761], Fresh[3760], Fresh[3759], Fresh[3758], Fresh[3757], Fresh[3756], Fresh[3755], Fresh[3754], Fresh[3753], Fresh[3752], Fresh[3751], Fresh[3750], Fresh[3749], Fresh[3748], Fresh[3747], Fresh[3746], Fresh[3745], Fresh[3744], Fresh[3743], Fresh[3742], Fresh[3741], Fresh[3740], Fresh[3739], Fresh[3738], Fresh[3737], Fresh[3736], Fresh[3735], Fresh[3734], Fresh[3733], Fresh[3732], Fresh[3731], Fresh[3730], Fresh[3729], Fresh[3728], Fresh[3727], Fresh[3726], Fresh[3725], Fresh[3724], Fresh[3723], Fresh[3722], Fresh[3721], Fresh[3720], Fresh[3719], Fresh[3718], Fresh[3717], Fresh[3716], Fresh[3715], Fresh[3714], Fresh[3713], Fresh[3712], Fresh[3711], Fresh[3710], Fresh[3709], Fresh[3708], Fresh[3707], Fresh[3706], Fresh[3705], Fresh[3704], Fresh[3703], Fresh[3702], Fresh[3701], Fresh[3700], Fresh[3699], Fresh[3698], Fresh[3697], Fresh[3696], Fresh[3695], Fresh[3694], Fresh[3693], Fresh[3692], Fresh[3691], Fresh[3690], Fresh[3689], Fresh[3688], Fresh[3687], Fresh[3686], Fresh[3685], Fresh[3684], Fresh[3683], Fresh[3682], Fresh[3681], Fresh[3680], Fresh[3679], Fresh[3678], Fresh[3677], Fresh[3676], Fresh[3675], Fresh[3674], Fresh[3673], Fresh[3672], Fresh[3671], Fresh[3670], Fresh[3669], Fresh[3668], Fresh[3667], Fresh[3666], Fresh[3665], Fresh[3664], Fresh[3663], Fresh[3662], Fresh[3661], Fresh[3660], Fresh[3659], Fresh[3658], Fresh[3657], Fresh[3656], Fresh[3655], Fresh[3654], Fresh[3653], Fresh[3652], Fresh[3651], Fresh[3650], Fresh[3649], Fresh[3648], Fresh[3647], Fresh[3646], Fresh[3645], Fresh[3644], Fresh[3643], Fresh[3642], Fresh[3641], Fresh[3640], Fresh[3639], Fresh[3638], Fresh[3637], Fresh[3636], Fresh[3635], Fresh[3634], Fresh[3633], Fresh[3632], Fresh[3631], Fresh[3630], Fresh[3629], Fresh[3628], Fresh[3627], Fresh[3626], Fresh[3625], Fresh[3624], Fresh[3623], Fresh[3622], Fresh[3621], Fresh[3620], Fresh[3619], Fresh[3618], Fresh[3617], Fresh[3616], Fresh[3615], Fresh[3614], Fresh[3613], Fresh[3612], Fresh[3611], Fresh[3610], Fresh[3609], Fresh[3608], Fresh[3607], Fresh[3606], Fresh[3605], Fresh[3604], Fresh[3603], Fresh[3602], Fresh[3601], Fresh[3600], Fresh[3599], Fresh[3598], Fresh[3597], Fresh[3596], Fresh[3595], Fresh[3594], Fresh[3593], Fresh[3592], Fresh[3591], Fresh[3590], Fresh[3589], Fresh[3588], Fresh[3587], Fresh[3586], Fresh[3585], Fresh[3584], Fresh[3583], Fresh[3582], Fresh[3581], Fresh[3580], Fresh[3579], Fresh[3578], Fresh[3577], Fresh[3576], Fresh[3575], Fresh[3574], Fresh[3573], Fresh[3572], Fresh[3571], Fresh[3570], Fresh[3569], Fresh[3568], Fresh[3567], Fresh[3566], Fresh[3565], Fresh[3564], Fresh[3563], Fresh[3562], Fresh[3561], Fresh[3560], Fresh[3559], Fresh[3558], Fresh[3557], Fresh[3556], Fresh[3555], Fresh[3554], Fresh[3553], Fresh[3552], Fresh[3551], Fresh[3550], Fresh[3549], Fresh[3548], Fresh[3547], Fresh[3546], Fresh[3545], Fresh[3544], Fresh[3543], Fresh[3542], Fresh[3541], Fresh[3540], Fresh[3539], Fresh[3538], Fresh[3537], Fresh[3536], Fresh[3535], Fresh[3534], Fresh[3533], Fresh[3532], Fresh[3531], Fresh[3530], Fresh[3529], Fresh[3528], Fresh[3527], Fresh[3526], Fresh[3525], Fresh[3524], Fresh[3523], Fresh[3522], Fresh[3521], Fresh[3520], Fresh[3519], Fresh[3518], Fresh[3517], Fresh[3516], Fresh[3515], Fresh[3514], Fresh[3513], Fresh[3512], Fresh[3511], Fresh[3510], Fresh[3509], Fresh[3508], Fresh[3507], Fresh[3506], Fresh[3505], Fresh[3504], Fresh[3503], Fresh[3502], Fresh[3501], Fresh[3500], Fresh[3499], Fresh[3498], Fresh[3497], Fresh[3496], Fresh[3495], Fresh[3494], Fresh[3493], Fresh[3492], Fresh[3491], Fresh[3490], Fresh[3489], Fresh[3488], Fresh[3487], Fresh[3486], Fresh[3485], Fresh[3484], Fresh[3483], Fresh[3482], Fresh[3481], Fresh[3480], Fresh[3479], Fresh[3478], Fresh[3477], Fresh[3476], Fresh[3475], Fresh[3474], Fresh[3473], Fresh[3472], Fresh[3471], Fresh[3470], Fresh[3469], Fresh[3468], Fresh[3467], Fresh[3466], Fresh[3465], Fresh[3464], Fresh[3463], Fresh[3462], Fresh[3461], Fresh[3460], Fresh[3459], Fresh[3458], Fresh[3457], Fresh[3456], Fresh[3455], Fresh[3454], Fresh[3453], Fresh[3452], Fresh[3451], Fresh[3450], Fresh[3449], Fresh[3448], Fresh[3447], Fresh[3446], Fresh[3445], Fresh[3444], Fresh[3443], Fresh[3442], Fresh[3441], Fresh[3440], Fresh[3439], Fresh[3438], Fresh[3437], Fresh[3436], Fresh[3435], Fresh[3434], Fresh[3433], Fresh[3432], Fresh[3431], Fresh[3430], Fresh[3429], Fresh[3428], Fresh[3427], Fresh[3426], Fresh[3425], Fresh[3424], Fresh[3423], Fresh[3422], Fresh[3421], Fresh[3420], Fresh[3419], Fresh[3418], Fresh[3417], Fresh[3416], Fresh[3415], Fresh[3414], Fresh[3413], Fresh[3412], Fresh[3411], Fresh[3410], Fresh[3409], Fresh[3408], Fresh[3407], Fresh[3406], Fresh[3405], Fresh[3404], Fresh[3403], Fresh[3402], Fresh[3401], Fresh[3400], Fresh[3399], Fresh[3398], Fresh[3397], Fresh[3396], Fresh[3395], Fresh[3394], Fresh[3393], Fresh[3392], Fresh[3391], Fresh[3390], Fresh[3389], Fresh[3388], Fresh[3387], Fresh[3386], Fresh[3385], Fresh[3384], Fresh[3383], Fresh[3382], Fresh[3381], Fresh[3380], Fresh[3379], Fresh[3378], Fresh[3377], Fresh[3376], Fresh[3375], Fresh[3374], Fresh[3373], Fresh[3372], Fresh[3371], Fresh[3370], Fresh[3369], Fresh[3368], Fresh[3367], Fresh[3366], Fresh[3365], Fresh[3364], Fresh[3363], Fresh[3362], Fresh[3361], Fresh[3360], Fresh[3359], Fresh[3358], Fresh[3357], Fresh[3356], Fresh[3355], Fresh[3354], Fresh[3353], Fresh[3352], Fresh[3351], Fresh[3350], Fresh[3349], Fresh[3348], Fresh[3347], Fresh[3346], Fresh[3345], Fresh[3344], Fresh[3343], Fresh[3342], Fresh[3341], Fresh[3340], Fresh[3339], Fresh[3338], Fresh[3337], Fresh[3336], Fresh[3335], Fresh[3334], Fresh[3333], Fresh[3332], Fresh[3331], Fresh[3330], Fresh[3329], Fresh[3328], Fresh[3327], Fresh[3326], Fresh[3325], Fresh[3324], Fresh[3323], Fresh[3322], Fresh[3321], Fresh[3320], Fresh[3319], Fresh[3318], Fresh[3317], Fresh[3316], Fresh[3315], Fresh[3314], Fresh[3313], Fresh[3312], Fresh[3311], Fresh[3310], Fresh[3309], Fresh[3308], Fresh[3307], Fresh[3306], Fresh[3305], Fresh[3304], Fresh[3303], Fresh[3302], Fresh[3301], Fresh[3300], Fresh[3299], Fresh[3298], Fresh[3297], Fresh[3296], Fresh[3295], Fresh[3294], Fresh[3293], Fresh[3292], Fresh[3291], Fresh[3290], Fresh[3289], Fresh[3288], Fresh[3287], Fresh[3286], Fresh[3285], Fresh[3284], Fresh[3283], Fresh[3282], Fresh[3281], Fresh[3280], Fresh[3279], Fresh[3278], Fresh[3277], Fresh[3276], Fresh[3275], Fresh[3274], Fresh[3273], Fresh[3272], Fresh[3271], Fresh[3270], Fresh[3269], Fresh[3268], Fresh[3267], Fresh[3266], Fresh[3265], Fresh[3264], Fresh[3263], Fresh[3262], Fresh[3261], Fresh[3260], Fresh[3259], Fresh[3258], Fresh[3257], Fresh[3256], Fresh[3255], Fresh[3254], Fresh[3253], Fresh[3252], Fresh[3251], Fresh[3250], Fresh[3249], Fresh[3248], Fresh[3247], Fresh[3246], Fresh[3245], Fresh[3244], Fresh[3243], Fresh[3242], Fresh[3241], Fresh[3240], Fresh[3239], Fresh[3238], Fresh[3237], Fresh[3236], Fresh[3235], Fresh[3234], Fresh[3233], Fresh[3232], Fresh[3231], Fresh[3230], Fresh[3229], Fresh[3228], Fresh[3227], Fresh[3226], Fresh[3225], Fresh[3224], Fresh[3223], Fresh[3222], Fresh[3221], Fresh[3220], Fresh[3219], Fresh[3218], Fresh[3217], Fresh[3216], Fresh[3215], Fresh[3214], Fresh[3213], Fresh[3212], Fresh[3211], Fresh[3210], Fresh[3209], Fresh[3208], Fresh[3207], Fresh[3206], Fresh[3205], Fresh[3204], Fresh[3203], Fresh[3202], Fresh[3201], Fresh[3200], Fresh[3199], Fresh[3198], Fresh[3197], Fresh[3196], Fresh[3195], Fresh[3194], Fresh[3193], Fresh[3192], Fresh[3191], Fresh[3190], Fresh[3189], Fresh[3188], Fresh[3187], Fresh[3186], Fresh[3185], Fresh[3184], Fresh[3183], Fresh[3182], Fresh[3181], Fresh[3180], Fresh[3179], Fresh[3178], Fresh[3177], Fresh[3176], Fresh[3175], Fresh[3174], Fresh[3173], Fresh[3172], Fresh[3171], Fresh[3170], Fresh[3169], Fresh[3168], Fresh[3167], Fresh[3166], Fresh[3165], Fresh[3164], Fresh[3163], Fresh[3162], Fresh[3161], Fresh[3160], Fresh[3159], Fresh[3158], Fresh[3157], Fresh[3156], Fresh[3155], Fresh[3154], Fresh[3153], Fresh[3152], Fresh[3151], Fresh[3150], Fresh[3149], Fresh[3148], Fresh[3147], Fresh[3146], Fresh[3145], Fresh[3144], Fresh[3143], Fresh[3142], Fresh[3141], Fresh[3140], Fresh[3139], Fresh[3138], Fresh[3137], Fresh[3136], Fresh[3135], Fresh[3134], Fresh[3133], Fresh[3132], Fresh[3131], Fresh[3130], Fresh[3129], Fresh[3128], Fresh[3127], Fresh[3126], Fresh[3125], Fresh[3124], Fresh[3123], Fresh[3122], Fresh[3121], Fresh[3120], Fresh[3119], Fresh[3118], Fresh[3117], Fresh[3116], Fresh[3115], Fresh[3114], Fresh[3113], Fresh[3112], Fresh[3111], Fresh[3110], Fresh[3109], Fresh[3108], Fresh[3107], Fresh[3106], Fresh[3105], Fresh[3104], Fresh[3103], Fresh[3102], Fresh[3101], Fresh[3100], Fresh[3099], Fresh[3098], Fresh[3097], Fresh[3096], Fresh[3095], Fresh[3094], Fresh[3093], Fresh[3092], Fresh[3091], Fresh[3090], Fresh[3089], Fresh[3088], Fresh[3087], Fresh[3086], Fresh[3085], Fresh[3084], Fresh[3083], Fresh[3082], Fresh[3081], Fresh[3080], Fresh[3079], Fresh[3078], Fresh[3077], Fresh[3076], Fresh[3075], Fresh[3074], Fresh[3073], Fresh[3072], Fresh[3071], Fresh[3070], Fresh[3069], Fresh[3068], Fresh[3067], Fresh[3066], Fresh[3065], Fresh[3064], Fresh[3063], Fresh[3062], Fresh[3061], Fresh[3060], Fresh[3059], Fresh[3058], Fresh[3057], Fresh[3056], Fresh[3055], Fresh[3054], Fresh[3053], Fresh[3052], Fresh[3051], Fresh[3050], Fresh[3049], Fresh[3048], Fresh[3047], Fresh[3046], Fresh[3045], Fresh[3044], Fresh[3043], Fresh[3042], Fresh[3041], Fresh[3040], Fresh[3039], Fresh[3038], Fresh[3037], Fresh[3036], Fresh[3035], Fresh[3034], Fresh[3033], Fresh[3032], Fresh[3031], Fresh[3030], Fresh[3029], Fresh[3028], Fresh[3027], Fresh[3026], Fresh[3025], Fresh[3024], Fresh[3023], Fresh[3022], Fresh[3021], Fresh[3020], Fresh[3019], Fresh[3018], Fresh[3017], Fresh[3016], Fresh[3015], Fresh[3014], Fresh[3013], Fresh[3012], Fresh[3011], Fresh[3010], Fresh[3009], Fresh[3008], Fresh[3007], Fresh[3006], Fresh[3005], Fresh[3004], Fresh[3003], Fresh[3002], Fresh[3001], Fresh[3000], Fresh[2999], Fresh[2998], Fresh[2997], Fresh[2996], Fresh[2995], Fresh[2994], Fresh[2993], Fresh[2992], Fresh[2991], Fresh[2990], Fresh[2989], Fresh[2988], Fresh[2987], Fresh[2986], Fresh[2985], Fresh[2984], Fresh[2983], Fresh[2982], Fresh[2981], Fresh[2980], Fresh[2979], Fresh[2978], Fresh[2977], Fresh[2976], Fresh[2975], Fresh[2974], Fresh[2973], Fresh[2972], Fresh[2971], Fresh[2970], Fresh[2969], Fresh[2968], Fresh[2967], Fresh[2966], Fresh[2965], Fresh[2964], Fresh[2963], Fresh[2962], Fresh[2961], Fresh[2960], Fresh[2959], Fresh[2958], Fresh[2957], Fresh[2956], Fresh[2955], Fresh[2954], Fresh[2953], Fresh[2952], Fresh[2951], Fresh[2950], Fresh[2949], Fresh[2948], Fresh[2947], Fresh[2946], Fresh[2945], Fresh[2944], Fresh[2943], Fresh[2942], Fresh[2941], Fresh[2940], Fresh[2939], Fresh[2938], Fresh[2937], Fresh[2936], Fresh[2935], Fresh[2934], Fresh[2933], Fresh[2932], Fresh[2931], Fresh[2930], Fresh[2929], Fresh[2928], Fresh[2927], Fresh[2926], Fresh[2925], Fresh[2924], Fresh[2923], Fresh[2922], Fresh[2921], Fresh[2920], Fresh[2919], Fresh[2918], Fresh[2917], Fresh[2916], Fresh[2915], Fresh[2914], Fresh[2913], Fresh[2912], Fresh[2911], Fresh[2910], Fresh[2909], Fresh[2908], Fresh[2907], Fresh[2906], Fresh[2905], Fresh[2904], Fresh[2903], Fresh[2902], Fresh[2901], Fresh[2900], Fresh[2899], Fresh[2898], Fresh[2897], Fresh[2896], Fresh[2895], Fresh[2894], Fresh[2893], Fresh[2892], Fresh[2891], Fresh[2890], Fresh[2889], Fresh[2888], Fresh[2887], Fresh[2886], Fresh[2885], Fresh[2884], Fresh[2883], Fresh[2882], Fresh[2881], Fresh[2880], Fresh[2879], Fresh[2878], Fresh[2877], Fresh[2876], Fresh[2875], Fresh[2874], Fresh[2873], Fresh[2872], Fresh[2871], Fresh[2870], Fresh[2869], Fresh[2868], Fresh[2867], Fresh[2866], Fresh[2865], Fresh[2864], Fresh[2863], Fresh[2862], Fresh[2861], Fresh[2860], Fresh[2859], Fresh[2858], Fresh[2857], Fresh[2856], Fresh[2855], Fresh[2854], Fresh[2853], Fresh[2852], Fresh[2851], Fresh[2850], Fresh[2849], Fresh[2848], Fresh[2847], Fresh[2846], Fresh[2845], Fresh[2844], Fresh[2843], Fresh[2842], Fresh[2841], Fresh[2840], Fresh[2839], Fresh[2838], Fresh[2837], Fresh[2836], Fresh[2835], Fresh[2834], Fresh[2833], Fresh[2832], Fresh[2831], Fresh[2830], Fresh[2829], Fresh[2828], Fresh[2827], Fresh[2826], Fresh[2825], Fresh[2824], Fresh[2823], Fresh[2822], Fresh[2821], Fresh[2820], Fresh[2819], Fresh[2818], Fresh[2817], Fresh[2816], Fresh[2815], Fresh[2814], Fresh[2813], Fresh[2812], Fresh[2811], Fresh[2810], Fresh[2809], Fresh[2808], Fresh[2807], Fresh[2806], Fresh[2805], Fresh[2804], Fresh[2803], Fresh[2802], Fresh[2801], Fresh[2800], Fresh[2799], Fresh[2798], Fresh[2797], Fresh[2796], Fresh[2795], Fresh[2794], Fresh[2793], Fresh[2792], Fresh[2791], Fresh[2790], Fresh[2789], Fresh[2788], Fresh[2787], Fresh[2786], Fresh[2785], Fresh[2784], Fresh[2783], Fresh[2782], Fresh[2781], Fresh[2780], Fresh[2779], Fresh[2778], Fresh[2777], Fresh[2776], Fresh[2775], Fresh[2774], Fresh[2773], Fresh[2772], Fresh[2771], Fresh[2770], Fresh[2769], Fresh[2768], Fresh[2767], Fresh[2766], Fresh[2765], Fresh[2764], Fresh[2763], Fresh[2762], Fresh[2761], Fresh[2760], Fresh[2759], Fresh[2758], Fresh[2757], Fresh[2756], Fresh[2755], Fresh[2754], Fresh[2753], Fresh[2752], Fresh[2751], Fresh[2750], Fresh[2749], Fresh[2748], Fresh[2747], Fresh[2746], Fresh[2745], Fresh[2744], Fresh[2743], Fresh[2742], Fresh[2741], Fresh[2740], Fresh[2739], Fresh[2738], Fresh[2737], Fresh[2736], Fresh[2735], Fresh[2734], Fresh[2733], Fresh[2732], Fresh[2731], Fresh[2730], Fresh[2729], Fresh[2728], Fresh[2727], Fresh[2726], Fresh[2725], Fresh[2724], Fresh[2723], Fresh[2722], Fresh[2721], Fresh[2720], Fresh[2719], Fresh[2718], Fresh[2717], Fresh[2716], Fresh[2715], Fresh[2714], Fresh[2713], Fresh[2712], Fresh[2711], Fresh[2710], Fresh[2709], Fresh[2708], Fresh[2707], Fresh[2706], Fresh[2705], Fresh[2704], Fresh[2703], Fresh[2702], Fresh[2701], Fresh[2700], Fresh[2699], Fresh[2698], Fresh[2697], Fresh[2696], Fresh[2695], Fresh[2694], Fresh[2693], Fresh[2692], Fresh[2691], Fresh[2690], Fresh[2689], Fresh[2688], Fresh[2687], Fresh[2686], Fresh[2685], Fresh[2684], Fresh[2683], Fresh[2682], Fresh[2681], Fresh[2680], Fresh[2679], Fresh[2678], Fresh[2677], Fresh[2676], Fresh[2675], Fresh[2674], Fresh[2673], Fresh[2672], Fresh[2671], Fresh[2670], Fresh[2669], Fresh[2668], Fresh[2667], Fresh[2666], Fresh[2665], Fresh[2664], Fresh[2663], Fresh[2662], Fresh[2661], Fresh[2660], Fresh[2659], Fresh[2658], Fresh[2657], Fresh[2656], Fresh[2655], Fresh[2654], Fresh[2653], Fresh[2652], Fresh[2651], Fresh[2650], Fresh[2649], Fresh[2648], Fresh[2647], Fresh[2646], Fresh[2645], Fresh[2644], Fresh[2643], Fresh[2642], Fresh[2641], Fresh[2640], Fresh[2639], Fresh[2638], Fresh[2637], Fresh[2636], Fresh[2635], Fresh[2634], Fresh[2633], Fresh[2632], Fresh[2631], Fresh[2630], Fresh[2629], Fresh[2628], Fresh[2627], Fresh[2626], Fresh[2625], Fresh[2624], Fresh[2623], Fresh[2622], Fresh[2621], Fresh[2620], Fresh[2619], Fresh[2618], Fresh[2617], Fresh[2616], Fresh[2615], Fresh[2614], Fresh[2613], Fresh[2612], Fresh[2611], Fresh[2610], Fresh[2609], Fresh[2608], Fresh[2607], Fresh[2606], Fresh[2605], Fresh[2604], Fresh[2603], Fresh[2602], Fresh[2601], Fresh[2600], Fresh[2599], Fresh[2598], Fresh[2597], Fresh[2596], Fresh[2595], Fresh[2594], Fresh[2593], Fresh[2592], Fresh[2591], Fresh[2590], Fresh[2589], Fresh[2588], Fresh[2587], Fresh[2586], Fresh[2585], Fresh[2584], Fresh[2583], Fresh[2582], Fresh[2581], Fresh[2580], Fresh[2579], Fresh[2578], Fresh[2577], Fresh[2576], Fresh[2575], Fresh[2574], Fresh[2573], Fresh[2572], Fresh[2571], Fresh[2570], Fresh[2569], Fresh[2568], Fresh[2567], Fresh[2566], Fresh[2565], Fresh[2564], Fresh[2563], Fresh[2562], Fresh[2561], Fresh[2560], Fresh[2559], Fresh[2558], Fresh[2557], Fresh[2556], Fresh[2555], Fresh[2554], Fresh[2553], Fresh[2552], Fresh[2551], Fresh[2550], Fresh[2549], Fresh[2548], Fresh[2547], Fresh[2546], Fresh[2545], Fresh[2544], Fresh[2543], Fresh[2542], Fresh[2541], Fresh[2540], Fresh[2539], Fresh[2538], Fresh[2537], Fresh[2536], Fresh[2535], Fresh[2534], Fresh[2533], Fresh[2532], Fresh[2531], Fresh[2530], Fresh[2529], Fresh[2528], Fresh[2527], Fresh[2526], Fresh[2525], Fresh[2524], Fresh[2523], Fresh[2522], Fresh[2521], Fresh[2520], Fresh[2519], Fresh[2518], Fresh[2517], Fresh[2516], Fresh[2515], Fresh[2514], Fresh[2513], Fresh[2512], Fresh[2511], Fresh[2510], Fresh[2509], Fresh[2508], Fresh[2507], Fresh[2506], Fresh[2505], Fresh[2504], Fresh[2503], Fresh[2502], Fresh[2501], Fresh[2500], Fresh[2499], Fresh[2498], Fresh[2497], Fresh[2496], Fresh[2495], Fresh[2494], Fresh[2493], Fresh[2492], Fresh[2491], Fresh[2490], Fresh[2489], Fresh[2488], Fresh[2487], Fresh[2486], Fresh[2485], Fresh[2484], Fresh[2483], Fresh[2482], Fresh[2481], Fresh[2480], Fresh[2479], Fresh[2478], Fresh[2477], Fresh[2476], Fresh[2475], Fresh[2474], Fresh[2473], Fresh[2472], Fresh[2471], Fresh[2470], Fresh[2469], Fresh[2468], Fresh[2467], Fresh[2466], Fresh[2465], Fresh[2464], Fresh[2463], Fresh[2462], Fresh[2461], Fresh[2460], Fresh[2459], Fresh[2458], Fresh[2457], Fresh[2456], Fresh[2455], Fresh[2454], Fresh[2453], Fresh[2452], Fresh[2451], Fresh[2450], Fresh[2449], Fresh[2448], Fresh[2447], Fresh[2446], Fresh[2445], Fresh[2444], Fresh[2443], Fresh[2442], Fresh[2441], Fresh[2440], Fresh[2439], Fresh[2438], Fresh[2437], Fresh[2436], Fresh[2435], Fresh[2434], Fresh[2433], Fresh[2432], Fresh[2431], Fresh[2430], Fresh[2429], Fresh[2428], Fresh[2427], Fresh[2426], Fresh[2425], Fresh[2424], Fresh[2423], Fresh[2422], Fresh[2421], Fresh[2420], Fresh[2419], Fresh[2418], Fresh[2417], Fresh[2416], Fresh[2415], Fresh[2414], Fresh[2413], Fresh[2412], Fresh[2411], Fresh[2410], Fresh[2409], Fresh[2408], Fresh[2407], Fresh[2406], Fresh[2405], Fresh[2404], Fresh[2403], Fresh[2402], Fresh[2401], Fresh[2400], Fresh[2399], Fresh[2398], Fresh[2397], Fresh[2396], Fresh[2395], Fresh[2394], Fresh[2393], Fresh[2392], Fresh[2391], Fresh[2390], Fresh[2389], Fresh[2388], Fresh[2387], Fresh[2386], Fresh[2385], Fresh[2384], Fresh[2383], Fresh[2382], Fresh[2381], Fresh[2380], Fresh[2379], Fresh[2378], Fresh[2377], Fresh[2376], Fresh[2375], Fresh[2374], Fresh[2373], Fresh[2372], Fresh[2371], Fresh[2370], Fresh[2369], Fresh[2368], Fresh[2367], Fresh[2366], Fresh[2365], Fresh[2364], Fresh[2363], Fresh[2362], Fresh[2361], Fresh[2360], Fresh[2359], Fresh[2358], Fresh[2357], Fresh[2356], Fresh[2355], Fresh[2354], Fresh[2353], Fresh[2352], Fresh[2351], Fresh[2350], Fresh[2349], Fresh[2348], Fresh[2347], Fresh[2346], Fresh[2345], Fresh[2344], Fresh[2343], Fresh[2342], Fresh[2341], Fresh[2340], Fresh[2339], Fresh[2338], Fresh[2337], Fresh[2336], Fresh[2335], Fresh[2334], Fresh[2333], Fresh[2332], Fresh[2331], Fresh[2330], Fresh[2329], Fresh[2328], Fresh[2327], Fresh[2326], Fresh[2325], Fresh[2324], Fresh[2323], Fresh[2322], Fresh[2321], Fresh[2320], Fresh[2319], Fresh[2318], Fresh[2317], Fresh[2316], Fresh[2315], Fresh[2314], Fresh[2313], Fresh[2312], Fresh[2311], Fresh[2310], Fresh[2309], Fresh[2308], Fresh[2307], Fresh[2306], Fresh[2305], Fresh[2304], Fresh[2303], Fresh[2302], Fresh[2301], Fresh[2300], Fresh[2299], Fresh[2298], Fresh[2297], Fresh[2296], Fresh[2295], Fresh[2294], Fresh[2293], Fresh[2292], Fresh[2291], Fresh[2290], Fresh[2289], Fresh[2288], Fresh[2287], Fresh[2286], Fresh[2285], Fresh[2284], Fresh[2283], Fresh[2282], Fresh[2281], Fresh[2280], Fresh[2279], Fresh[2278], Fresh[2277], Fresh[2276], Fresh[2275], Fresh[2274], Fresh[2273], Fresh[2272], Fresh[2271], Fresh[2270], Fresh[2269], Fresh[2268], Fresh[2267], Fresh[2266], Fresh[2265], Fresh[2264], Fresh[2263], Fresh[2262], Fresh[2261], Fresh[2260], Fresh[2259], Fresh[2258], Fresh[2257], Fresh[2256], Fresh[2255], Fresh[2254], Fresh[2253], Fresh[2252], Fresh[2251], Fresh[2250], Fresh[2249], Fresh[2248], Fresh[2247], Fresh[2246], Fresh[2245], Fresh[2244], Fresh[2243], Fresh[2242], Fresh[2241], Fresh[2240], Fresh[2239], Fresh[2238], Fresh[2237], Fresh[2236], Fresh[2235], Fresh[2234], Fresh[2233], Fresh[2232], Fresh[2231], Fresh[2230], Fresh[2229], Fresh[2228], Fresh[2227], Fresh[2226], Fresh[2225], Fresh[2224], Fresh[2223], Fresh[2222], Fresh[2221], Fresh[2220], Fresh[2219], Fresh[2218], Fresh[2217], Fresh[2216], Fresh[2215], Fresh[2214], Fresh[2213], Fresh[2212], Fresh[2211], Fresh[2210], Fresh[2209], Fresh[2208], Fresh[2207], Fresh[2206], Fresh[2205], Fresh[2204], Fresh[2203], Fresh[2202], Fresh[2201], Fresh[2200], Fresh[2199], Fresh[2198], Fresh[2197], Fresh[2196], Fresh[2195], Fresh[2194], Fresh[2193], Fresh[2192], Fresh[2191], Fresh[2190], Fresh[2189], Fresh[2188], Fresh[2187], Fresh[2186], Fresh[2185], Fresh[2184], Fresh[2183], Fresh[2182], Fresh[2181], Fresh[2180], Fresh[2179], Fresh[2178], Fresh[2177], Fresh[2176], Fresh[2175], Fresh[2174], Fresh[2173], Fresh[2172], Fresh[2171], Fresh[2170], Fresh[2169], Fresh[2168], Fresh[2167], Fresh[2166], Fresh[2165], Fresh[2164], Fresh[2163], Fresh[2162], Fresh[2161], Fresh[2160], Fresh[2159], Fresh[2158], Fresh[2157], Fresh[2156], Fresh[2155], Fresh[2154], Fresh[2153], Fresh[2152], Fresh[2151], Fresh[2150], Fresh[2149], Fresh[2148], Fresh[2147], Fresh[2146], Fresh[2145], Fresh[2144], Fresh[2143], Fresh[2142], Fresh[2141], Fresh[2140], Fresh[2139], Fresh[2138], Fresh[2137], Fresh[2136], Fresh[2135], Fresh[2134], Fresh[2133], Fresh[2132], Fresh[2131], Fresh[2130], Fresh[2129], Fresh[2128], Fresh[2127], Fresh[2126], Fresh[2125], Fresh[2124], Fresh[2123], Fresh[2122], Fresh[2121], Fresh[2120], Fresh[2119], Fresh[2118], Fresh[2117], Fresh[2116], Fresh[2115], Fresh[2114], Fresh[2113], Fresh[2112], Fresh[2111], Fresh[2110], Fresh[2109], Fresh[2108], Fresh[2107], Fresh[2106], Fresh[2105], Fresh[2104], Fresh[2103], Fresh[2102], Fresh[2101], Fresh[2100], Fresh[2099], Fresh[2098], Fresh[2097], Fresh[2096], Fresh[2095], Fresh[2094], Fresh[2093], Fresh[2092], Fresh[2091], Fresh[2090], Fresh[2089], Fresh[2088], Fresh[2087], Fresh[2086], Fresh[2085], Fresh[2084], Fresh[2083], Fresh[2082], Fresh[2081], Fresh[2080], Fresh[2079], Fresh[2078], Fresh[2077], Fresh[2076], Fresh[2075], Fresh[2074], Fresh[2073], Fresh[2072], Fresh[2071], Fresh[2070], Fresh[2069], Fresh[2068], Fresh[2067], Fresh[2066], Fresh[2065], Fresh[2064], Fresh[2063], Fresh[2062], Fresh[2061], Fresh[2060], Fresh[2059], Fresh[2058], Fresh[2057], Fresh[2056], Fresh[2055], Fresh[2054], Fresh[2053], Fresh[2052], Fresh[2051], Fresh[2050], Fresh[2049], Fresh[2048], Fresh[2047], Fresh[2046], Fresh[2045], Fresh[2044], Fresh[2043], Fresh[2042], Fresh[2041], Fresh[2040], Fresh[2039], Fresh[2038], Fresh[2037], Fresh[2036], Fresh[2035], Fresh[2034], Fresh[2033], Fresh[2032], Fresh[2031], Fresh[2030], Fresh[2029], Fresh[2028], Fresh[2027], Fresh[2026], Fresh[2025], Fresh[2024], Fresh[2023], Fresh[2022], Fresh[2021], Fresh[2020], Fresh[2019], Fresh[2018], Fresh[2017], Fresh[2016], Fresh[2015], Fresh[2014], Fresh[2013], Fresh[2012], Fresh[2011], Fresh[2010], Fresh[2009], Fresh[2008], Fresh[2007], Fresh[2006], Fresh[2005], Fresh[2004], Fresh[2003], Fresh[2002], Fresh[2001], Fresh[2000], Fresh[1999], Fresh[1998], Fresh[1997], Fresh[1996], Fresh[1995], Fresh[1994], Fresh[1993], Fresh[1992], Fresh[1991], Fresh[1990], Fresh[1989], Fresh[1988], Fresh[1987], Fresh[1986], Fresh[1985], Fresh[1984], Fresh[1983], Fresh[1982], Fresh[1981], Fresh[1980], Fresh[1979], Fresh[1978], Fresh[1977], Fresh[1976], Fresh[1975], Fresh[1974], Fresh[1973], Fresh[1972], Fresh[1971], Fresh[1970], Fresh[1969], Fresh[1968], Fresh[1967], Fresh[1966], Fresh[1965], Fresh[1964], Fresh[1963], Fresh[1962], Fresh[1961], Fresh[1960], Fresh[1959], Fresh[1958], Fresh[1957], Fresh[1956], Fresh[1955], Fresh[1954], Fresh[1953], Fresh[1952], Fresh[1951], Fresh[1950], Fresh[1949], Fresh[1948], Fresh[1947], Fresh[1946], Fresh[1945], Fresh[1944], Fresh[1943], Fresh[1942], Fresh[1941], Fresh[1940], Fresh[1939], Fresh[1938], Fresh[1937], Fresh[1936], Fresh[1935], Fresh[1934], Fresh[1933], Fresh[1932], Fresh[1931], Fresh[1930], Fresh[1929], Fresh[1928], Fresh[1927], Fresh[1926], Fresh[1925], Fresh[1924], Fresh[1923], Fresh[1922], Fresh[1921], Fresh[1920], Fresh[1919], Fresh[1918], Fresh[1917], Fresh[1916], Fresh[1915], Fresh[1914], Fresh[1913], Fresh[1912], Fresh[1911], Fresh[1910], Fresh[1909], Fresh[1908], Fresh[1907], Fresh[1906], Fresh[1905], Fresh[1904], Fresh[1903], Fresh[1902], Fresh[1901], Fresh[1900], Fresh[1899], Fresh[1898], Fresh[1897], Fresh[1896], Fresh[1895], Fresh[1894], Fresh[1893], Fresh[1892], Fresh[1891], Fresh[1890], Fresh[1889], Fresh[1888], Fresh[1887], Fresh[1886], Fresh[1885], Fresh[1884], Fresh[1883], Fresh[1882], Fresh[1881], Fresh[1880], Fresh[1879], Fresh[1878], Fresh[1877], Fresh[1876], Fresh[1875], Fresh[1874], Fresh[1873], Fresh[1872], Fresh[1871], Fresh[1870], Fresh[1869], Fresh[1868], Fresh[1867], Fresh[1866], Fresh[1865], Fresh[1864], Fresh[1863], Fresh[1862], Fresh[1861], Fresh[1860], Fresh[1859], Fresh[1858], Fresh[1857], Fresh[1856], Fresh[1855], Fresh[1854], Fresh[1853], Fresh[1852], Fresh[1851], Fresh[1850], Fresh[1849], Fresh[1848], Fresh[1847], Fresh[1846], Fresh[1845], Fresh[1844], Fresh[1843], Fresh[1842], Fresh[1841], Fresh[1840], Fresh[1839], Fresh[1838], Fresh[1837], Fresh[1836], Fresh[1835], Fresh[1834], Fresh[1833], Fresh[1832], Fresh[1831], Fresh[1830], Fresh[1829], Fresh[1828], Fresh[1827], Fresh[1826], Fresh[1825], Fresh[1824], Fresh[1823], Fresh[1822], Fresh[1821], Fresh[1820], Fresh[1819], Fresh[1818], Fresh[1817], Fresh[1816], Fresh[1815], Fresh[1814], Fresh[1813], Fresh[1812], Fresh[1811], Fresh[1810], Fresh[1809], Fresh[1808], Fresh[1807], Fresh[1806], Fresh[1805], Fresh[1804], Fresh[1803], Fresh[1802], Fresh[1801], Fresh[1800], Fresh[1799], Fresh[1798], Fresh[1797], Fresh[1796], Fresh[1795], Fresh[1794], Fresh[1793], Fresh[1792], Fresh[1791], Fresh[1790], Fresh[1789], Fresh[1788], Fresh[1787], Fresh[1786], Fresh[1785], Fresh[1784], Fresh[1783], Fresh[1782], Fresh[1781], Fresh[1780], Fresh[1779], Fresh[1778], Fresh[1777], Fresh[1776], Fresh[1775], Fresh[1774], Fresh[1773], Fresh[1772], Fresh[1771], Fresh[1770], Fresh[1769], Fresh[1768], Fresh[1767], Fresh[1766], Fresh[1765], Fresh[1764], Fresh[1763], Fresh[1762], Fresh[1761], Fresh[1760], Fresh[1759], Fresh[1758], Fresh[1757], Fresh[1756], Fresh[1755], Fresh[1754], Fresh[1753], Fresh[1752], Fresh[1751], Fresh[1750], Fresh[1749], Fresh[1748], Fresh[1747], Fresh[1746], Fresh[1745], Fresh[1744], Fresh[1743], Fresh[1742], Fresh[1741], Fresh[1740], Fresh[1739], Fresh[1738], Fresh[1737], Fresh[1736], Fresh[1735], Fresh[1734], Fresh[1733], Fresh[1732], Fresh[1731], Fresh[1730], Fresh[1729], Fresh[1728], Fresh[1727], Fresh[1726], Fresh[1725], Fresh[1724], Fresh[1723], Fresh[1722], Fresh[1721], Fresh[1720], Fresh[1719], Fresh[1718], Fresh[1717], Fresh[1716], Fresh[1715], Fresh[1714], Fresh[1713], Fresh[1712], Fresh[1711], Fresh[1710], Fresh[1709], Fresh[1708], Fresh[1707], Fresh[1706], Fresh[1705], Fresh[1704], Fresh[1703], Fresh[1702], Fresh[1701], Fresh[1700], Fresh[1699], Fresh[1698], Fresh[1697], Fresh[1696], Fresh[1695], Fresh[1694], Fresh[1693], Fresh[1692], Fresh[1691], Fresh[1690], Fresh[1689], Fresh[1688], Fresh[1687], Fresh[1686], Fresh[1685], Fresh[1684], Fresh[1683], Fresh[1682], Fresh[1681], Fresh[1680], Fresh[1679], Fresh[1678], Fresh[1677], Fresh[1676], Fresh[1675], Fresh[1674], Fresh[1673], Fresh[1672], Fresh[1671], Fresh[1670], Fresh[1669], Fresh[1668], Fresh[1667], Fresh[1666], Fresh[1665], Fresh[1664], Fresh[1663], Fresh[1662], Fresh[1661], Fresh[1660], Fresh[1659], Fresh[1658], Fresh[1657], Fresh[1656], Fresh[1655], Fresh[1654], Fresh[1653], Fresh[1652], Fresh[1651], Fresh[1650], Fresh[1649], Fresh[1648], Fresh[1647], Fresh[1646], Fresh[1645], Fresh[1644], Fresh[1643], Fresh[1642], Fresh[1641], Fresh[1640], Fresh[1639], Fresh[1638], Fresh[1637], Fresh[1636], Fresh[1635], Fresh[1634], Fresh[1633], Fresh[1632], Fresh[1631], Fresh[1630], Fresh[1629], Fresh[1628], Fresh[1627], Fresh[1626], Fresh[1625], Fresh[1624], Fresh[1623], Fresh[1622], Fresh[1621], Fresh[1620], Fresh[1619], Fresh[1618], Fresh[1617], Fresh[1616], Fresh[1615], Fresh[1614], Fresh[1613], Fresh[1612], Fresh[1611], Fresh[1610], Fresh[1609], Fresh[1608], Fresh[1607], Fresh[1606], Fresh[1605], Fresh[1604], Fresh[1603], Fresh[1602], Fresh[1601], Fresh[1600], Fresh[1599], Fresh[1598], Fresh[1597], Fresh[1596], Fresh[1595], Fresh[1594], Fresh[1593], Fresh[1592], Fresh[1591], Fresh[1590], Fresh[1589], Fresh[1588], Fresh[1587], Fresh[1586], Fresh[1585], Fresh[1584], Fresh[1583], Fresh[1582], Fresh[1581], Fresh[1580], Fresh[1579], Fresh[1578], Fresh[1577], Fresh[1576], Fresh[1575], Fresh[1574], Fresh[1573], Fresh[1572], Fresh[1571], Fresh[1570], Fresh[1569], Fresh[1568], Fresh[1567], Fresh[1566], Fresh[1565], Fresh[1564], Fresh[1563], Fresh[1562], Fresh[1561], Fresh[1560], Fresh[1559], Fresh[1558], Fresh[1557], Fresh[1556], Fresh[1555], Fresh[1554], Fresh[1553], Fresh[1552], Fresh[1551], Fresh[1550], Fresh[1549], Fresh[1548], Fresh[1547], Fresh[1546], Fresh[1545], Fresh[1544], Fresh[1543], Fresh[1542], Fresh[1541], Fresh[1540], Fresh[1539], Fresh[1538], Fresh[1537], Fresh[1536], Fresh[1535], Fresh[1534], Fresh[1533], Fresh[1532], Fresh[1531], Fresh[1530], Fresh[1529], Fresh[1528], Fresh[1527], Fresh[1526], Fresh[1525], Fresh[1524], Fresh[1523], Fresh[1522], Fresh[1521], Fresh[1520], Fresh[1519], Fresh[1518], Fresh[1517], Fresh[1516], Fresh[1515], Fresh[1514], Fresh[1513], Fresh[1512], Fresh[1511], Fresh[1510], Fresh[1509], Fresh[1508], Fresh[1507], Fresh[1506], Fresh[1505], Fresh[1504], Fresh[1503], Fresh[1502], Fresh[1501], Fresh[1500], Fresh[1499], Fresh[1498], Fresh[1497], Fresh[1496], Fresh[1495], Fresh[1494], Fresh[1493], Fresh[1492], Fresh[1491], Fresh[1490], Fresh[1489], Fresh[1488], Fresh[1487], Fresh[1486], Fresh[1485], Fresh[1484], Fresh[1483], Fresh[1482], Fresh[1481], Fresh[1480], Fresh[1479], Fresh[1478], Fresh[1477], Fresh[1476], Fresh[1475], Fresh[1474], Fresh[1473], Fresh[1472], Fresh[1471], Fresh[1470], Fresh[1469], Fresh[1468], Fresh[1467], Fresh[1466], Fresh[1465], Fresh[1464], Fresh[1463], Fresh[1462], Fresh[1461], Fresh[1460], Fresh[1459], Fresh[1458], Fresh[1457], Fresh[1456], Fresh[1455], Fresh[1454], Fresh[1453], Fresh[1452], Fresh[1451], Fresh[1450], Fresh[1449], Fresh[1448], Fresh[1447], Fresh[1446], Fresh[1445], Fresh[1444], Fresh[1443], Fresh[1442], Fresh[1441], Fresh[1440], Fresh[1439], Fresh[1438], Fresh[1437], Fresh[1436], Fresh[1435], Fresh[1434], Fresh[1433], Fresh[1432], Fresh[1431], Fresh[1430], Fresh[1429], Fresh[1428], Fresh[1427], Fresh[1426], Fresh[1425], Fresh[1424], Fresh[1423], Fresh[1422], Fresh[1421], Fresh[1420], Fresh[1419], Fresh[1418], Fresh[1417], Fresh[1416], Fresh[1415], Fresh[1414], Fresh[1413], Fresh[1412], Fresh[1411], Fresh[1410], Fresh[1409], Fresh[1408], Fresh[1407], Fresh[1406], Fresh[1405], Fresh[1404], Fresh[1403], Fresh[1402], Fresh[1401], Fresh[1400], Fresh[1399], Fresh[1398], Fresh[1397], Fresh[1396], Fresh[1395], Fresh[1394], Fresh[1393], Fresh[1392], Fresh[1391], Fresh[1390], Fresh[1389], Fresh[1388], Fresh[1387], Fresh[1386], Fresh[1385], Fresh[1384], Fresh[1383], Fresh[1382], Fresh[1381], Fresh[1380], Fresh[1379], Fresh[1378], Fresh[1377], Fresh[1376], Fresh[1375], Fresh[1374], Fresh[1373], Fresh[1372], Fresh[1371], Fresh[1370], Fresh[1369], Fresh[1368], Fresh[1367], Fresh[1366], Fresh[1365], Fresh[1364], Fresh[1363], Fresh[1362], Fresh[1361], Fresh[1360], Fresh[1359], Fresh[1358], Fresh[1357], Fresh[1356], Fresh[1355], Fresh[1354], Fresh[1353], Fresh[1352], Fresh[1351], Fresh[1350], Fresh[1349], Fresh[1348], Fresh[1347], Fresh[1346], Fresh[1345], Fresh[1344], Fresh[1343], Fresh[1342], Fresh[1341], Fresh[1340], Fresh[1339], Fresh[1338], Fresh[1337], Fresh[1336], Fresh[1335], Fresh[1334], Fresh[1333], Fresh[1332], Fresh[1331], Fresh[1330], Fresh[1329], Fresh[1328], Fresh[1327], Fresh[1326], Fresh[1325], Fresh[1324], Fresh[1323], Fresh[1322], Fresh[1321], Fresh[1320], Fresh[1319], Fresh[1318], Fresh[1317], Fresh[1316], Fresh[1315], Fresh[1314], Fresh[1313], Fresh[1312], Fresh[1311], Fresh[1310], Fresh[1309], Fresh[1308], Fresh[1307], Fresh[1306], Fresh[1305], Fresh[1304], Fresh[1303], Fresh[1302], Fresh[1301], Fresh[1300], Fresh[1299], Fresh[1298], Fresh[1297], Fresh[1296], Fresh[1295], Fresh[1294], Fresh[1293], Fresh[1292], Fresh[1291], Fresh[1290], Fresh[1289], Fresh[1288], Fresh[1287], Fresh[1286], Fresh[1285], Fresh[1284], Fresh[1283], Fresh[1282], Fresh[1281], Fresh[1280], Fresh[1279], Fresh[1278], Fresh[1277], Fresh[1276], Fresh[1275], Fresh[1274], Fresh[1273], Fresh[1272], Fresh[1271], Fresh[1270], Fresh[1269], Fresh[1268], Fresh[1267], Fresh[1266], Fresh[1265], Fresh[1264], Fresh[1263], Fresh[1262], Fresh[1261], Fresh[1260], Fresh[1259], Fresh[1258], Fresh[1257], Fresh[1256], Fresh[1255], Fresh[1254], Fresh[1253], Fresh[1252], Fresh[1251], Fresh[1250], Fresh[1249], Fresh[1248], Fresh[1247], Fresh[1246], Fresh[1245], Fresh[1244], Fresh[1243], Fresh[1242], Fresh[1241], Fresh[1240], Fresh[1239], Fresh[1238], Fresh[1237], Fresh[1236], Fresh[1235], Fresh[1234], Fresh[1233], Fresh[1232], Fresh[1231], Fresh[1230], Fresh[1229], Fresh[1228], Fresh[1227], Fresh[1226], Fresh[1225], Fresh[1224], Fresh[1223], Fresh[1222], Fresh[1221], Fresh[1220], Fresh[1219], Fresh[1218], Fresh[1217], Fresh[1216], Fresh[1215], Fresh[1214], Fresh[1213], Fresh[1212], Fresh[1211], Fresh[1210], Fresh[1209], Fresh[1208], Fresh[1207], Fresh[1206], Fresh[1205], Fresh[1204], Fresh[1203], Fresh[1202], Fresh[1201], Fresh[1200], Fresh[1199], Fresh[1198], Fresh[1197], Fresh[1196], Fresh[1195], Fresh[1194], Fresh[1193], Fresh[1192], Fresh[1191], Fresh[1190], Fresh[1189], Fresh[1188], Fresh[1187], Fresh[1186], Fresh[1185], Fresh[1184], Fresh[1183], Fresh[1182], Fresh[1181], Fresh[1180], Fresh[1179], Fresh[1178], Fresh[1177], Fresh[1176], Fresh[1175], Fresh[1174], Fresh[1173], Fresh[1172], Fresh[1171], Fresh[1170], Fresh[1169], Fresh[1168], Fresh[1167], Fresh[1166], Fresh[1165], Fresh[1164], Fresh[1163], Fresh[1162], Fresh[1161], Fresh[1160], Fresh[1159], Fresh[1158], Fresh[1157], Fresh[1156], Fresh[1155], Fresh[1154], Fresh[1153], Fresh[1152], Fresh[1151], Fresh[1150], Fresh[1149], Fresh[1148], Fresh[1147], Fresh[1146], Fresh[1145], Fresh[1144], Fresh[1143], Fresh[1142], Fresh[1141], Fresh[1140], Fresh[1139], Fresh[1138], Fresh[1137], Fresh[1136], Fresh[1135], Fresh[1134], Fresh[1133], Fresh[1132], Fresh[1131], Fresh[1130], Fresh[1129], Fresh[1128], Fresh[1127], Fresh[1126], Fresh[1125], Fresh[1124], Fresh[1123], Fresh[1122], Fresh[1121], Fresh[1120], Fresh[1119], Fresh[1118], Fresh[1117], Fresh[1116], Fresh[1115], Fresh[1114], Fresh[1113], Fresh[1112], Fresh[1111], Fresh[1110], Fresh[1109], Fresh[1108], Fresh[1107], Fresh[1106], Fresh[1105], Fresh[1104], Fresh[1103], Fresh[1102], Fresh[1101], Fresh[1100], Fresh[1099], Fresh[1098], Fresh[1097], Fresh[1096], Fresh[1095], Fresh[1094], Fresh[1093], Fresh[1092], Fresh[1091], Fresh[1090], Fresh[1089], Fresh[1088], Fresh[1087], Fresh[1086], Fresh[1085], Fresh[1084], Fresh[1083], Fresh[1082], Fresh[1081], Fresh[1080], Fresh[1079], Fresh[1078], Fresh[1077], Fresh[1076], Fresh[1075], Fresh[1074], Fresh[1073], Fresh[1072], Fresh[1071], Fresh[1070], Fresh[1069], Fresh[1068], Fresh[1067], Fresh[1066], Fresh[1065], Fresh[1064], Fresh[1063], Fresh[1062], Fresh[1061], Fresh[1060], Fresh[1059], Fresh[1058], Fresh[1057], Fresh[1056], Fresh[1055], Fresh[1054], Fresh[1053], Fresh[1052], Fresh[1051], Fresh[1050], Fresh[1049], Fresh[1048], Fresh[1047], Fresh[1046], Fresh[1045], Fresh[1044], Fresh[1043], Fresh[1042], Fresh[1041], Fresh[1040], Fresh[1039], Fresh[1038], Fresh[1037], Fresh[1036], Fresh[1035], Fresh[1034], Fresh[1033], Fresh[1032], Fresh[1031], Fresh[1030], Fresh[1029], Fresh[1028], Fresh[1027], Fresh[1026], Fresh[1025], Fresh[1024], Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008], Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992], Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976], Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960], Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944], Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928], Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912], Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896], Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880], Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864], Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848], Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832], Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816], Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800], Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784], Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768], Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752], Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736], Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720], Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704], Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688], Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672], Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656], Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640], Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624], Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608], Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592], Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576], Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560], Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544], Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528], Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512], Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496], Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480], Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464], Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448], Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432], Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416], Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400], Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384], Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368], Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352], Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336], Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320], Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304], Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288], Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272], Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256], Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240], Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224], Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208], Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192], Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176], Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160], Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144], Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128], Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112], Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96], Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80], Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64], Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48], Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32], Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16], Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .out0 ({signal_2337, signal_2336, signal_2335, signal_2334, signal_2333, signal_2332, signal_2331, signal_2330, signal_2329, signal_2328, signal_2327, signal_2326, signal_2325, signal_2324, signal_2323, signal_2322, signal_2321, signal_2320, signal_2319, signal_2318, signal_2317, signal_2316, signal_2315, signal_2314, signal_2305, signal_2303, signal_2300, signal_2299, signal_2298, signal_1876, signal_1875, signal_1874, signal_1873, signal_1872, signal_1871, signal_1870, signal_1869, signal_1867, signal_1866, signal_1865, signal_1864, signal_1863, signal_1862, signal_1861, signal_1860, signal_1859, signal_1858, signal_1857, signal_1856, signal_1855, signal_1854, signal_1853, signal_1852, signal_1851, signal_1850, signal_1849, signal_1848, signal_1847, signal_1846, signal_1845, signal_1843, signal_1842, signal_1216, signal_1153}), .out1 ({signal_3109, signal_3108, signal_3107, signal_3106, signal_3105, signal_3104, signal_3103, signal_3102, signal_3101, signal_3100, signal_3099, signal_3098, signal_3097, signal_3096, signal_3095, signal_3094, signal_3093, signal_3092, signal_3091, signal_3090, signal_3089, signal_3088, signal_3087, signal_3086, signal_3085, signal_3084, signal_3083, signal_3082, signal_3081, signal_3080, signal_3079, signal_3078, signal_3077, signal_3076, signal_3075, signal_3074, signal_3073, signal_3072, signal_3071, signal_3070, signal_3069, signal_3068, signal_3067, signal_3066, signal_3065, signal_3064, signal_3063, signal_3062, signal_3061, signal_3060, signal_3059, signal_3058, signal_3057, signal_3056, signal_3055, signal_3054, signal_3053, signal_3052, signal_3051, signal_3050, signal_3049, signal_3048, signal_3047, signal_3046}) ) ;
    buf_clk cell_2062 ( .C (clk), .D (reset), .Q (signal_11952) ) ;
    buf_sca_clk cell_2063 ( .C (clk), .D (plaintext_s0[0]), .Q (signal_11953) ) ;
    buf_sca_clk cell_2064 ( .C (clk), .D (plaintext_s1[0]), .Q (signal_11954) ) ;
    buf_sca_clk cell_2065 ( .C (clk), .D (plaintext_s0[1]), .Q (signal_11955) ) ;
    buf_sca_clk cell_2066 ( .C (clk), .D (plaintext_s1[1]), .Q (signal_11956) ) ;
    buf_sca_clk cell_2067 ( .C (clk), .D (plaintext_s0[2]), .Q (signal_11957) ) ;
    buf_sca_clk cell_2068 ( .C (clk), .D (plaintext_s1[2]), .Q (signal_11958) ) ;
    buf_sca_clk cell_2069 ( .C (clk), .D (plaintext_s0[3]), .Q (signal_11959) ) ;
    buf_sca_clk cell_2070 ( .C (clk), .D (plaintext_s1[3]), .Q (signal_11960) ) ;
    buf_sca_clk cell_2071 ( .C (clk), .D (plaintext_s0[4]), .Q (signal_11961) ) ;
    buf_sca_clk cell_2072 ( .C (clk), .D (plaintext_s1[4]), .Q (signal_11962) ) ;
    buf_sca_clk cell_2073 ( .C (clk), .D (plaintext_s0[5]), .Q (signal_11963) ) ;
    buf_sca_clk cell_2074 ( .C (clk), .D (plaintext_s1[5]), .Q (signal_11964) ) ;
    buf_sca_clk cell_2075 ( .C (clk), .D (plaintext_s0[6]), .Q (signal_11965) ) ;
    buf_sca_clk cell_2076 ( .C (clk), .D (plaintext_s1[6]), .Q (signal_11966) ) ;
    buf_sca_clk cell_2077 ( .C (clk), .D (plaintext_s0[7]), .Q (signal_11967) ) ;
    buf_sca_clk cell_2078 ( .C (clk), .D (plaintext_s1[7]), .Q (signal_11968) ) ;
    buf_sca_clk cell_2079 ( .C (clk), .D (plaintext_s0[8]), .Q (signal_11969) ) ;
    buf_sca_clk cell_2080 ( .C (clk), .D (plaintext_s1[8]), .Q (signal_11970) ) ;
    buf_sca_clk cell_2081 ( .C (clk), .D (plaintext_s0[9]), .Q (signal_11971) ) ;
    buf_sca_clk cell_2082 ( .C (clk), .D (plaintext_s1[9]), .Q (signal_11972) ) ;
    buf_sca_clk cell_2083 ( .C (clk), .D (plaintext_s0[10]), .Q (signal_11973) ) ;
    buf_sca_clk cell_2084 ( .C (clk), .D (plaintext_s1[10]), .Q (signal_11974) ) ;
    buf_sca_clk cell_2085 ( .C (clk), .D (plaintext_s0[11]), .Q (signal_11975) ) ;
    buf_sca_clk cell_2086 ( .C (clk), .D (plaintext_s1[11]), .Q (signal_11976) ) ;
    buf_sca_clk cell_2087 ( .C (clk), .D (plaintext_s0[12]), .Q (signal_11977) ) ;
    buf_sca_clk cell_2088 ( .C (clk), .D (plaintext_s1[12]), .Q (signal_11978) ) ;
    buf_sca_clk cell_2089 ( .C (clk), .D (plaintext_s0[13]), .Q (signal_11979) ) ;
    buf_sca_clk cell_2090 ( .C (clk), .D (plaintext_s1[13]), .Q (signal_11980) ) ;
    buf_sca_clk cell_2091 ( .C (clk), .D (plaintext_s0[14]), .Q (signal_11981) ) ;
    buf_sca_clk cell_2092 ( .C (clk), .D (plaintext_s1[14]), .Q (signal_11982) ) ;
    buf_sca_clk cell_2093 ( .C (clk), .D (plaintext_s0[15]), .Q (signal_11983) ) ;
    buf_sca_clk cell_2094 ( .C (clk), .D (plaintext_s1[15]), .Q (signal_11984) ) ;
    buf_sca_clk cell_2095 ( .C (clk), .D (plaintext_s0[16]), .Q (signal_11985) ) ;
    buf_sca_clk cell_2096 ( .C (clk), .D (plaintext_s1[16]), .Q (signal_11986) ) ;
    buf_sca_clk cell_2097 ( .C (clk), .D (plaintext_s0[17]), .Q (signal_11987) ) ;
    buf_sca_clk cell_2098 ( .C (clk), .D (plaintext_s1[17]), .Q (signal_11988) ) ;
    buf_sca_clk cell_2099 ( .C (clk), .D (plaintext_s0[18]), .Q (signal_11989) ) ;
    buf_sca_clk cell_2100 ( .C (clk), .D (plaintext_s1[18]), .Q (signal_11990) ) ;
    buf_sca_clk cell_2101 ( .C (clk), .D (plaintext_s0[19]), .Q (signal_11991) ) ;
    buf_sca_clk cell_2102 ( .C (clk), .D (plaintext_s1[19]), .Q (signal_11992) ) ;
    buf_sca_clk cell_2103 ( .C (clk), .D (plaintext_s0[20]), .Q (signal_11993) ) ;
    buf_sca_clk cell_2104 ( .C (clk), .D (plaintext_s1[20]), .Q (signal_11994) ) ;
    buf_sca_clk cell_2105 ( .C (clk), .D (plaintext_s0[21]), .Q (signal_11995) ) ;
    buf_sca_clk cell_2106 ( .C (clk), .D (plaintext_s1[21]), .Q (signal_11996) ) ;
    buf_sca_clk cell_2107 ( .C (clk), .D (plaintext_s0[22]), .Q (signal_11997) ) ;
    buf_sca_clk cell_2108 ( .C (clk), .D (plaintext_s1[22]), .Q (signal_11998) ) ;
    buf_sca_clk cell_2109 ( .C (clk), .D (plaintext_s0[23]), .Q (signal_11999) ) ;
    buf_sca_clk cell_2110 ( .C (clk), .D (plaintext_s1[23]), .Q (signal_12000) ) ;
    buf_sca_clk cell_2111 ( .C (clk), .D (plaintext_s0[24]), .Q (signal_12001) ) ;
    buf_sca_clk cell_2112 ( .C (clk), .D (plaintext_s1[24]), .Q (signal_12002) ) ;
    buf_sca_clk cell_2113 ( .C (clk), .D (plaintext_s0[25]), .Q (signal_12003) ) ;
    buf_sca_clk cell_2114 ( .C (clk), .D (plaintext_s1[25]), .Q (signal_12004) ) ;
    buf_sca_clk cell_2115 ( .C (clk), .D (plaintext_s0[26]), .Q (signal_12005) ) ;
    buf_sca_clk cell_2116 ( .C (clk), .D (plaintext_s1[26]), .Q (signal_12006) ) ;
    buf_sca_clk cell_2117 ( .C (clk), .D (plaintext_s0[27]), .Q (signal_12007) ) ;
    buf_sca_clk cell_2118 ( .C (clk), .D (plaintext_s1[27]), .Q (signal_12008) ) ;
    buf_sca_clk cell_2119 ( .C (clk), .D (plaintext_s0[28]), .Q (signal_12009) ) ;
    buf_sca_clk cell_2120 ( .C (clk), .D (plaintext_s1[28]), .Q (signal_12010) ) ;
    buf_sca_clk cell_2121 ( .C (clk), .D (plaintext_s0[29]), .Q (signal_12011) ) ;
    buf_sca_clk cell_2122 ( .C (clk), .D (plaintext_s1[29]), .Q (signal_12012) ) ;
    buf_sca_clk cell_2123 ( .C (clk), .D (plaintext_s0[30]), .Q (signal_12013) ) ;
    buf_sca_clk cell_2124 ( .C (clk), .D (plaintext_s1[30]), .Q (signal_12014) ) ;
    buf_sca_clk cell_2125 ( .C (clk), .D (plaintext_s0[31]), .Q (signal_12015) ) ;
    buf_sca_clk cell_2126 ( .C (clk), .D (plaintext_s1[31]), .Q (signal_12016) ) ;
    buf_clk cell_2127 ( .C (clk), .D (signal_1218), .Q (signal_12017) ) ;
    buf_clk cell_2128 ( .C (clk), .D (signal_394), .Q (signal_12018) ) ;
    buf_clk cell_2129 ( .C (clk), .D (signal_1219), .Q (signal_12019) ) ;
    buf_clk cell_2130 ( .C (clk), .D (signal_393), .Q (signal_12020) ) ;
    buf_sca_clk cell_2131 ( .C (clk), .D (signal_1777), .Q (signal_12021) ) ;
    buf_sca_clk cell_2132 ( .C (clk), .D (signal_2499), .Q (signal_12022) ) ;
    buf_clk cell_2133 ( .C (clk), .D (signal_1226), .Q (signal_12023) ) ;
    buf_sca_clk cell_2134 ( .C (clk), .D (signal_1776), .Q (signal_12024) ) ;
    buf_sca_clk cell_2135 ( .C (clk), .D (signal_2502), .Q (signal_12025) ) ;
    buf_clk cell_2136 ( .C (clk), .D (signal_1225), .Q (signal_12026) ) ;
    buf_sca_clk cell_2137 ( .C (clk), .D (signal_1775), .Q (signal_12027) ) ;
    buf_sca_clk cell_2138 ( .C (clk), .D (signal_2505), .Q (signal_12028) ) ;
    buf_clk cell_2139 ( .C (clk), .D (signal_1224), .Q (signal_12029) ) ;
    buf_sca_clk cell_2140 ( .C (clk), .D (signal_1774), .Q (signal_12030) ) ;
    buf_sca_clk cell_2141 ( .C (clk), .D (signal_2508), .Q (signal_12031) ) ;
    buf_clk cell_2142 ( .C (clk), .D (signal_1223), .Q (signal_12032) ) ;
    buf_sca_clk cell_2143 ( .C (clk), .D (signal_1773), .Q (signal_12033) ) ;
    buf_sca_clk cell_2144 ( .C (clk), .D (signal_2511), .Q (signal_12034) ) ;
    buf_clk cell_2145 ( .C (clk), .D (signal_1222), .Q (signal_12035) ) ;
    buf_sca_clk cell_2146 ( .C (clk), .D (signal_1772), .Q (signal_12036) ) ;
    buf_sca_clk cell_2147 ( .C (clk), .D (signal_2514), .Q (signal_12037) ) ;
    buf_clk cell_2148 ( .C (clk), .D (signal_1221), .Q (signal_12038) ) ;
    buf_sca_clk cell_2149 ( .C (clk), .D (signal_1771), .Q (signal_12039) ) ;
    buf_sca_clk cell_2150 ( .C (clk), .D (signal_2517), .Q (signal_12040) ) ;
    buf_sca_clk cell_2151 ( .C (clk), .D (signal_1770), .Q (signal_12041) ) ;
    buf_sca_clk cell_2152 ( .C (clk), .D (signal_2520), .Q (signal_12042) ) ;
    buf_sca_clk cell_2153 ( .C (clk), .D (signal_1769), .Q (signal_12043) ) ;
    buf_sca_clk cell_2154 ( .C (clk), .D (signal_2631), .Q (signal_12044) ) ;
    buf_sca_clk cell_2155 ( .C (clk), .D (signal_1768), .Q (signal_12045) ) ;
    buf_sca_clk cell_2156 ( .C (clk), .D (signal_2634), .Q (signal_12046) ) ;
    buf_sca_clk cell_2157 ( .C (clk), .D (signal_1767), .Q (signal_12047) ) ;
    buf_sca_clk cell_2158 ( .C (clk), .D (signal_2637), .Q (signal_12048) ) ;
    buf_sca_clk cell_2159 ( .C (clk), .D (signal_1766), .Q (signal_12049) ) ;
    buf_sca_clk cell_2160 ( .C (clk), .D (signal_2640), .Q (signal_12050) ) ;
    buf_sca_clk cell_2161 ( .C (clk), .D (signal_1765), .Q (signal_12051) ) ;
    buf_sca_clk cell_2162 ( .C (clk), .D (signal_2643), .Q (signal_12052) ) ;
    buf_sca_clk cell_2163 ( .C (clk), .D (signal_1764), .Q (signal_12053) ) ;
    buf_sca_clk cell_2164 ( .C (clk), .D (signal_2646), .Q (signal_12054) ) ;
    buf_sca_clk cell_2165 ( .C (clk), .D (signal_1763), .Q (signal_12055) ) ;
    buf_sca_clk cell_2166 ( .C (clk), .D (signal_2649), .Q (signal_12056) ) ;
    buf_sca_clk cell_2167 ( .C (clk), .D (signal_1762), .Q (signal_12057) ) ;
    buf_sca_clk cell_2168 ( .C (clk), .D (signal_2652), .Q (signal_12058) ) ;
    buf_sca_clk cell_2169 ( .C (clk), .D (signal_1761), .Q (signal_12059) ) ;
    buf_sca_clk cell_2170 ( .C (clk), .D (signal_2382), .Q (signal_12060) ) ;
    buf_sca_clk cell_2171 ( .C (clk), .D (signal_1760), .Q (signal_12061) ) ;
    buf_sca_clk cell_2172 ( .C (clk), .D (signal_2385), .Q (signal_12062) ) ;
    buf_sca_clk cell_2173 ( .C (clk), .D (signal_1759), .Q (signal_12063) ) ;
    buf_sca_clk cell_2174 ( .C (clk), .D (signal_2388), .Q (signal_12064) ) ;
    buf_sca_clk cell_2175 ( .C (clk), .D (signal_1758), .Q (signal_12065) ) ;
    buf_sca_clk cell_2176 ( .C (clk), .D (signal_2391), .Q (signal_12066) ) ;
    buf_sca_clk cell_2177 ( .C (clk), .D (signal_1757), .Q (signal_12067) ) ;
    buf_sca_clk cell_2178 ( .C (clk), .D (signal_2394), .Q (signal_12068) ) ;
    buf_sca_clk cell_2179 ( .C (clk), .D (signal_1756), .Q (signal_12069) ) ;
    buf_sca_clk cell_2180 ( .C (clk), .D (signal_2397), .Q (signal_12070) ) ;
    buf_sca_clk cell_2181 ( .C (clk), .D (signal_1755), .Q (signal_12071) ) ;
    buf_sca_clk cell_2182 ( .C (clk), .D (signal_2400), .Q (signal_12072) ) ;
    buf_sca_clk cell_2183 ( .C (clk), .D (signal_1754), .Q (signal_12073) ) ;
    buf_sca_clk cell_2184 ( .C (clk), .D (signal_2403), .Q (signal_12074) ) ;
    buf_sca_clk cell_2185 ( .C (clk), .D (signal_1753), .Q (signal_12075) ) ;
    buf_sca_clk cell_2186 ( .C (clk), .D (signal_2472), .Q (signal_12076) ) ;
    buf_sca_clk cell_2187 ( .C (clk), .D (signal_1752), .Q (signal_12077) ) ;
    buf_sca_clk cell_2188 ( .C (clk), .D (signal_2475), .Q (signal_12078) ) ;
    buf_sca_clk cell_2189 ( .C (clk), .D (signal_1751), .Q (signal_12079) ) ;
    buf_sca_clk cell_2190 ( .C (clk), .D (signal_2478), .Q (signal_12080) ) ;
    buf_sca_clk cell_2191 ( .C (clk), .D (signal_1750), .Q (signal_12081) ) ;
    buf_sca_clk cell_2192 ( .C (clk), .D (signal_2481), .Q (signal_12082) ) ;
    buf_sca_clk cell_2193 ( .C (clk), .D (signal_1749), .Q (signal_12083) ) ;
    buf_sca_clk cell_2194 ( .C (clk), .D (signal_2484), .Q (signal_12084) ) ;
    buf_sca_clk cell_2195 ( .C (clk), .D (signal_1748), .Q (signal_12085) ) ;
    buf_sca_clk cell_2196 ( .C (clk), .D (signal_2487), .Q (signal_12086) ) ;
    buf_sca_clk cell_2197 ( .C (clk), .D (signal_1747), .Q (signal_12087) ) ;
    buf_sca_clk cell_2198 ( .C (clk), .D (signal_2493), .Q (signal_12088) ) ;
    buf_sca_clk cell_2199 ( .C (clk), .D (signal_1746), .Q (signal_12089) ) ;
    buf_sca_clk cell_2200 ( .C (clk), .D (signal_2496), .Q (signal_12090) ) ;
    buf_sca_clk cell_2201 ( .C (clk), .D (key_s0[0]), .Q (signal_12091) ) ;
    buf_sca_clk cell_2202 ( .C (clk), .D (key_s1[0]), .Q (signal_12092) ) ;
    buf_sca_clk cell_2203 ( .C (clk), .D (key_s0[1]), .Q (signal_12093) ) ;
    buf_sca_clk cell_2204 ( .C (clk), .D (key_s1[1]), .Q (signal_12094) ) ;
    buf_sca_clk cell_2205 ( .C (clk), .D (key_s0[2]), .Q (signal_12095) ) ;
    buf_sca_clk cell_2206 ( .C (clk), .D (key_s1[2]), .Q (signal_12096) ) ;
    buf_sca_clk cell_2207 ( .C (clk), .D (key_s0[3]), .Q (signal_12097) ) ;
    buf_sca_clk cell_2208 ( .C (clk), .D (key_s1[3]), .Q (signal_12098) ) ;
    buf_sca_clk cell_2209 ( .C (clk), .D (key_s0[4]), .Q (signal_12099) ) ;
    buf_sca_clk cell_2210 ( .C (clk), .D (key_s1[4]), .Q (signal_12100) ) ;
    buf_sca_clk cell_2211 ( .C (clk), .D (key_s0[5]), .Q (signal_12101) ) ;
    buf_sca_clk cell_2212 ( .C (clk), .D (key_s1[5]), .Q (signal_12102) ) ;
    buf_sca_clk cell_2213 ( .C (clk), .D (key_s0[6]), .Q (signal_12103) ) ;
    buf_sca_clk cell_2214 ( .C (clk), .D (key_s1[6]), .Q (signal_12104) ) ;
    buf_sca_clk cell_2215 ( .C (clk), .D (key_s0[7]), .Q (signal_12105) ) ;
    buf_sca_clk cell_2216 ( .C (clk), .D (key_s1[7]), .Q (signal_12106) ) ;
    buf_sca_clk cell_2217 ( .C (clk), .D (key_s0[8]), .Q (signal_12107) ) ;
    buf_sca_clk cell_2218 ( .C (clk), .D (key_s1[8]), .Q (signal_12108) ) ;
    buf_sca_clk cell_2219 ( .C (clk), .D (key_s0[9]), .Q (signal_12109) ) ;
    buf_sca_clk cell_2220 ( .C (clk), .D (key_s1[9]), .Q (signal_12110) ) ;
    buf_sca_clk cell_2221 ( .C (clk), .D (key_s0[10]), .Q (signal_12111) ) ;
    buf_sca_clk cell_2222 ( .C (clk), .D (key_s1[10]), .Q (signal_12112) ) ;
    buf_sca_clk cell_2223 ( .C (clk), .D (key_s0[11]), .Q (signal_12113) ) ;
    buf_sca_clk cell_2224 ( .C (clk), .D (key_s1[11]), .Q (signal_12114) ) ;
    buf_sca_clk cell_2225 ( .C (clk), .D (key_s0[12]), .Q (signal_12115) ) ;
    buf_sca_clk cell_2226 ( .C (clk), .D (key_s1[12]), .Q (signal_12116) ) ;
    buf_sca_clk cell_2227 ( .C (clk), .D (key_s0[13]), .Q (signal_12117) ) ;
    buf_sca_clk cell_2228 ( .C (clk), .D (key_s1[13]), .Q (signal_12118) ) ;
    buf_sca_clk cell_2229 ( .C (clk), .D (key_s0[14]), .Q (signal_12119) ) ;
    buf_sca_clk cell_2230 ( .C (clk), .D (key_s1[14]), .Q (signal_12120) ) ;
    buf_sca_clk cell_2231 ( .C (clk), .D (key_s0[15]), .Q (signal_12121) ) ;
    buf_sca_clk cell_2232 ( .C (clk), .D (key_s1[15]), .Q (signal_12122) ) ;
    buf_sca_clk cell_2233 ( .C (clk), .D (key_s0[16]), .Q (signal_12123) ) ;
    buf_sca_clk cell_2234 ( .C (clk), .D (key_s1[16]), .Q (signal_12124) ) ;
    buf_sca_clk cell_2235 ( .C (clk), .D (key_s0[17]), .Q (signal_12125) ) ;
    buf_sca_clk cell_2236 ( .C (clk), .D (key_s1[17]), .Q (signal_12126) ) ;
    buf_sca_clk cell_2237 ( .C (clk), .D (key_s0[18]), .Q (signal_12127) ) ;
    buf_sca_clk cell_2238 ( .C (clk), .D (key_s1[18]), .Q (signal_12128) ) ;
    buf_sca_clk cell_2239 ( .C (clk), .D (key_s0[19]), .Q (signal_12129) ) ;
    buf_sca_clk cell_2240 ( .C (clk), .D (key_s1[19]), .Q (signal_12130) ) ;
    buf_sca_clk cell_2241 ( .C (clk), .D (key_s0[20]), .Q (signal_12131) ) ;
    buf_sca_clk cell_2242 ( .C (clk), .D (key_s1[20]), .Q (signal_12132) ) ;
    buf_sca_clk cell_2243 ( .C (clk), .D (key_s0[21]), .Q (signal_12133) ) ;
    buf_sca_clk cell_2244 ( .C (clk), .D (key_s1[21]), .Q (signal_12134) ) ;
    buf_sca_clk cell_2245 ( .C (clk), .D (key_s0[22]), .Q (signal_12135) ) ;
    buf_sca_clk cell_2246 ( .C (clk), .D (key_s1[22]), .Q (signal_12136) ) ;
    buf_sca_clk cell_2247 ( .C (clk), .D (key_s0[23]), .Q (signal_12137) ) ;
    buf_sca_clk cell_2248 ( .C (clk), .D (key_s1[23]), .Q (signal_12138) ) ;
    buf_sca_clk cell_2249 ( .C (clk), .D (key_s0[24]), .Q (signal_12139) ) ;
    buf_sca_clk cell_2250 ( .C (clk), .D (key_s1[24]), .Q (signal_12140) ) ;
    buf_sca_clk cell_2251 ( .C (clk), .D (key_s0[25]), .Q (signal_12141) ) ;
    buf_sca_clk cell_2252 ( .C (clk), .D (key_s1[25]), .Q (signal_12142) ) ;
    buf_sca_clk cell_2253 ( .C (clk), .D (key_s0[26]), .Q (signal_12143) ) ;
    buf_sca_clk cell_2254 ( .C (clk), .D (key_s1[26]), .Q (signal_12144) ) ;
    buf_sca_clk cell_2255 ( .C (clk), .D (key_s0[27]), .Q (signal_12145) ) ;
    buf_sca_clk cell_2256 ( .C (clk), .D (key_s1[27]), .Q (signal_12146) ) ;
    buf_sca_clk cell_2257 ( .C (clk), .D (key_s0[28]), .Q (signal_12147) ) ;
    buf_sca_clk cell_2258 ( .C (clk), .D (key_s1[28]), .Q (signal_12148) ) ;
    buf_sca_clk cell_2259 ( .C (clk), .D (key_s0[29]), .Q (signal_12149) ) ;
    buf_sca_clk cell_2260 ( .C (clk), .D (key_s1[29]), .Q (signal_12150) ) ;
    buf_sca_clk cell_2261 ( .C (clk), .D (key_s0[30]), .Q (signal_12151) ) ;
    buf_sca_clk cell_2262 ( .C (clk), .D (key_s1[30]), .Q (signal_12152) ) ;
    buf_sca_clk cell_2263 ( .C (clk), .D (key_s0[31]), .Q (signal_12153) ) ;
    buf_sca_clk cell_2264 ( .C (clk), .D (key_s1[31]), .Q (signal_12154) ) ;
    buf_sca_clk cell_2265 ( .C (clk), .D (key_s0[32]), .Q (signal_12155) ) ;
    buf_sca_clk cell_2266 ( .C (clk), .D (key_s1[32]), .Q (signal_12156) ) ;
    buf_sca_clk cell_2267 ( .C (clk), .D (key_s0[33]), .Q (signal_12157) ) ;
    buf_sca_clk cell_2268 ( .C (clk), .D (key_s1[33]), .Q (signal_12158) ) ;
    buf_sca_clk cell_2269 ( .C (clk), .D (key_s0[34]), .Q (signal_12159) ) ;
    buf_sca_clk cell_2270 ( .C (clk), .D (key_s1[34]), .Q (signal_12160) ) ;
    buf_sca_clk cell_2271 ( .C (clk), .D (key_s0[35]), .Q (signal_12161) ) ;
    buf_sca_clk cell_2272 ( .C (clk), .D (key_s1[35]), .Q (signal_12162) ) ;
    buf_sca_clk cell_2273 ( .C (clk), .D (key_s0[36]), .Q (signal_12163) ) ;
    buf_sca_clk cell_2274 ( .C (clk), .D (key_s1[36]), .Q (signal_12164) ) ;
    buf_sca_clk cell_2275 ( .C (clk), .D (key_s0[37]), .Q (signal_12165) ) ;
    buf_sca_clk cell_2276 ( .C (clk), .D (key_s1[37]), .Q (signal_12166) ) ;
    buf_sca_clk cell_2277 ( .C (clk), .D (key_s0[38]), .Q (signal_12167) ) ;
    buf_sca_clk cell_2278 ( .C (clk), .D (key_s1[38]), .Q (signal_12168) ) ;
    buf_sca_clk cell_2279 ( .C (clk), .D (key_s0[39]), .Q (signal_12169) ) ;
    buf_sca_clk cell_2280 ( .C (clk), .D (key_s1[39]), .Q (signal_12170) ) ;
    buf_sca_clk cell_2281 ( .C (clk), .D (key_s0[40]), .Q (signal_12171) ) ;
    buf_sca_clk cell_2282 ( .C (clk), .D (key_s1[40]), .Q (signal_12172) ) ;
    buf_sca_clk cell_2283 ( .C (clk), .D (key_s0[41]), .Q (signal_12173) ) ;
    buf_sca_clk cell_2284 ( .C (clk), .D (key_s1[41]), .Q (signal_12174) ) ;
    buf_sca_clk cell_2285 ( .C (clk), .D (key_s0[42]), .Q (signal_12175) ) ;
    buf_sca_clk cell_2286 ( .C (clk), .D (key_s1[42]), .Q (signal_12176) ) ;
    buf_sca_clk cell_2287 ( .C (clk), .D (key_s0[43]), .Q (signal_12177) ) ;
    buf_sca_clk cell_2288 ( .C (clk), .D (key_s1[43]), .Q (signal_12178) ) ;
    buf_sca_clk cell_2289 ( .C (clk), .D (key_s0[44]), .Q (signal_12179) ) ;
    buf_sca_clk cell_2290 ( .C (clk), .D (key_s1[44]), .Q (signal_12180) ) ;
    buf_sca_clk cell_2291 ( .C (clk), .D (key_s0[45]), .Q (signal_12181) ) ;
    buf_sca_clk cell_2292 ( .C (clk), .D (key_s1[45]), .Q (signal_12182) ) ;
    buf_sca_clk cell_2293 ( .C (clk), .D (key_s0[46]), .Q (signal_12183) ) ;
    buf_sca_clk cell_2294 ( .C (clk), .D (key_s1[46]), .Q (signal_12184) ) ;
    buf_sca_clk cell_2295 ( .C (clk), .D (key_s0[47]), .Q (signal_12185) ) ;
    buf_sca_clk cell_2296 ( .C (clk), .D (key_s1[47]), .Q (signal_12186) ) ;
    buf_sca_clk cell_2297 ( .C (clk), .D (key_s0[48]), .Q (signal_12187) ) ;
    buf_sca_clk cell_2298 ( .C (clk), .D (key_s1[48]), .Q (signal_12188) ) ;
    buf_sca_clk cell_2299 ( .C (clk), .D (key_s0[49]), .Q (signal_12189) ) ;
    buf_sca_clk cell_2300 ( .C (clk), .D (key_s1[49]), .Q (signal_12190) ) ;
    buf_sca_clk cell_2301 ( .C (clk), .D (key_s0[50]), .Q (signal_12191) ) ;
    buf_sca_clk cell_2302 ( .C (clk), .D (key_s1[50]), .Q (signal_12192) ) ;
    buf_sca_clk cell_2303 ( .C (clk), .D (key_s0[51]), .Q (signal_12193) ) ;
    buf_sca_clk cell_2304 ( .C (clk), .D (key_s1[51]), .Q (signal_12194) ) ;
    buf_sca_clk cell_2305 ( .C (clk), .D (key_s0[52]), .Q (signal_12195) ) ;
    buf_sca_clk cell_2306 ( .C (clk), .D (key_s1[52]), .Q (signal_12196) ) ;
    buf_sca_clk cell_2307 ( .C (clk), .D (key_s0[53]), .Q (signal_12197) ) ;
    buf_sca_clk cell_2308 ( .C (clk), .D (key_s1[53]), .Q (signal_12198) ) ;
    buf_sca_clk cell_2309 ( .C (clk), .D (key_s0[54]), .Q (signal_12199) ) ;
    buf_sca_clk cell_2310 ( .C (clk), .D (key_s1[54]), .Q (signal_12200) ) ;
    buf_sca_clk cell_2311 ( .C (clk), .D (key_s0[55]), .Q (signal_12201) ) ;
    buf_sca_clk cell_2312 ( .C (clk), .D (key_s1[55]), .Q (signal_12202) ) ;
    buf_sca_clk cell_2313 ( .C (clk), .D (key_s0[56]), .Q (signal_12203) ) ;
    buf_sca_clk cell_2314 ( .C (clk), .D (key_s1[56]), .Q (signal_12204) ) ;
    buf_sca_clk cell_2315 ( .C (clk), .D (key_s0[57]), .Q (signal_12205) ) ;
    buf_sca_clk cell_2316 ( .C (clk), .D (key_s1[57]), .Q (signal_12206) ) ;
    buf_sca_clk cell_2317 ( .C (clk), .D (key_s0[58]), .Q (signal_12207) ) ;
    buf_sca_clk cell_2318 ( .C (clk), .D (key_s1[58]), .Q (signal_12208) ) ;
    buf_sca_clk cell_2319 ( .C (clk), .D (key_s0[59]), .Q (signal_12209) ) ;
    buf_sca_clk cell_2320 ( .C (clk), .D (key_s1[59]), .Q (signal_12210) ) ;
    buf_sca_clk cell_2321 ( .C (clk), .D (key_s0[60]), .Q (signal_12211) ) ;
    buf_sca_clk cell_2322 ( .C (clk), .D (key_s1[60]), .Q (signal_12212) ) ;
    buf_sca_clk cell_2323 ( .C (clk), .D (key_s0[61]), .Q (signal_12213) ) ;
    buf_sca_clk cell_2324 ( .C (clk), .D (key_s1[61]), .Q (signal_12214) ) ;
    buf_sca_clk cell_2325 ( .C (clk), .D (key_s0[62]), .Q (signal_12215) ) ;
    buf_sca_clk cell_2326 ( .C (clk), .D (key_s1[62]), .Q (signal_12216) ) ;
    buf_sca_clk cell_2327 ( .C (clk), .D (key_s0[63]), .Q (signal_12217) ) ;
    buf_sca_clk cell_2328 ( .C (clk), .D (key_s1[63]), .Q (signal_12218) ) ;
    buf_sca_clk cell_2329 ( .C (clk), .D (key_s0[64]), .Q (signal_12219) ) ;
    buf_sca_clk cell_2330 ( .C (clk), .D (key_s1[64]), .Q (signal_12220) ) ;
    buf_sca_clk cell_2331 ( .C (clk), .D (key_s0[65]), .Q (signal_12221) ) ;
    buf_sca_clk cell_2332 ( .C (clk), .D (key_s1[65]), .Q (signal_12222) ) ;
    buf_sca_clk cell_2333 ( .C (clk), .D (key_s0[66]), .Q (signal_12223) ) ;
    buf_sca_clk cell_2334 ( .C (clk), .D (key_s1[66]), .Q (signal_12224) ) ;
    buf_sca_clk cell_2335 ( .C (clk), .D (key_s0[67]), .Q (signal_12225) ) ;
    buf_sca_clk cell_2336 ( .C (clk), .D (key_s1[67]), .Q (signal_12226) ) ;
    buf_sca_clk cell_2337 ( .C (clk), .D (key_s0[68]), .Q (signal_12227) ) ;
    buf_sca_clk cell_2338 ( .C (clk), .D (key_s1[68]), .Q (signal_12228) ) ;
    buf_sca_clk cell_2339 ( .C (clk), .D (key_s0[69]), .Q (signal_12229) ) ;
    buf_sca_clk cell_2340 ( .C (clk), .D (key_s1[69]), .Q (signal_12230) ) ;
    buf_sca_clk cell_2341 ( .C (clk), .D (key_s0[70]), .Q (signal_12231) ) ;
    buf_sca_clk cell_2342 ( .C (clk), .D (key_s1[70]), .Q (signal_12232) ) ;
    buf_sca_clk cell_2343 ( .C (clk), .D (key_s0[71]), .Q (signal_12233) ) ;
    buf_sca_clk cell_2344 ( .C (clk), .D (key_s1[71]), .Q (signal_12234) ) ;
    buf_sca_clk cell_2345 ( .C (clk), .D (key_s0[72]), .Q (signal_12235) ) ;
    buf_sca_clk cell_2346 ( .C (clk), .D (key_s1[72]), .Q (signal_12236) ) ;
    buf_sca_clk cell_2347 ( .C (clk), .D (key_s0[73]), .Q (signal_12237) ) ;
    buf_sca_clk cell_2348 ( .C (clk), .D (key_s1[73]), .Q (signal_12238) ) ;
    buf_sca_clk cell_2349 ( .C (clk), .D (key_s0[74]), .Q (signal_12239) ) ;
    buf_sca_clk cell_2350 ( .C (clk), .D (key_s1[74]), .Q (signal_12240) ) ;
    buf_sca_clk cell_2351 ( .C (clk), .D (key_s0[75]), .Q (signal_12241) ) ;
    buf_sca_clk cell_2352 ( .C (clk), .D (key_s1[75]), .Q (signal_12242) ) ;
    buf_sca_clk cell_2353 ( .C (clk), .D (key_s0[76]), .Q (signal_12243) ) ;
    buf_sca_clk cell_2354 ( .C (clk), .D (key_s1[76]), .Q (signal_12244) ) ;
    buf_sca_clk cell_2355 ( .C (clk), .D (key_s0[77]), .Q (signal_12245) ) ;
    buf_sca_clk cell_2356 ( .C (clk), .D (key_s1[77]), .Q (signal_12246) ) ;
    buf_sca_clk cell_2357 ( .C (clk), .D (key_s0[78]), .Q (signal_12247) ) ;
    buf_sca_clk cell_2358 ( .C (clk), .D (key_s1[78]), .Q (signal_12248) ) ;
    buf_sca_clk cell_2359 ( .C (clk), .D (key_s0[79]), .Q (signal_12249) ) ;
    buf_sca_clk cell_2360 ( .C (clk), .D (key_s1[79]), .Q (signal_12250) ) ;
    buf_sca_clk cell_2361 ( .C (clk), .D (key_s0[80]), .Q (signal_12251) ) ;
    buf_sca_clk cell_2362 ( .C (clk), .D (key_s1[80]), .Q (signal_12252) ) ;
    buf_sca_clk cell_2363 ( .C (clk), .D (key_s0[81]), .Q (signal_12253) ) ;
    buf_sca_clk cell_2364 ( .C (clk), .D (key_s1[81]), .Q (signal_12254) ) ;
    buf_sca_clk cell_2365 ( .C (clk), .D (key_s0[82]), .Q (signal_12255) ) ;
    buf_sca_clk cell_2366 ( .C (clk), .D (key_s1[82]), .Q (signal_12256) ) ;
    buf_sca_clk cell_2367 ( .C (clk), .D (key_s0[83]), .Q (signal_12257) ) ;
    buf_sca_clk cell_2368 ( .C (clk), .D (key_s1[83]), .Q (signal_12258) ) ;
    buf_sca_clk cell_2369 ( .C (clk), .D (key_s0[84]), .Q (signal_12259) ) ;
    buf_sca_clk cell_2370 ( .C (clk), .D (key_s1[84]), .Q (signal_12260) ) ;
    buf_sca_clk cell_2371 ( .C (clk), .D (key_s0[85]), .Q (signal_12261) ) ;
    buf_sca_clk cell_2372 ( .C (clk), .D (key_s1[85]), .Q (signal_12262) ) ;
    buf_sca_clk cell_2373 ( .C (clk), .D (key_s0[86]), .Q (signal_12263) ) ;
    buf_sca_clk cell_2374 ( .C (clk), .D (key_s1[86]), .Q (signal_12264) ) ;
    buf_sca_clk cell_2375 ( .C (clk), .D (key_s0[87]), .Q (signal_12265) ) ;
    buf_sca_clk cell_2376 ( .C (clk), .D (key_s1[87]), .Q (signal_12266) ) ;
    buf_sca_clk cell_2377 ( .C (clk), .D (key_s0[88]), .Q (signal_12267) ) ;
    buf_sca_clk cell_2378 ( .C (clk), .D (key_s1[88]), .Q (signal_12268) ) ;
    buf_sca_clk cell_2379 ( .C (clk), .D (key_s0[89]), .Q (signal_12269) ) ;
    buf_sca_clk cell_2380 ( .C (clk), .D (key_s1[89]), .Q (signal_12270) ) ;
    buf_sca_clk cell_2381 ( .C (clk), .D (key_s0[90]), .Q (signal_12271) ) ;
    buf_sca_clk cell_2382 ( .C (clk), .D (key_s1[90]), .Q (signal_12272) ) ;
    buf_sca_clk cell_2383 ( .C (clk), .D (key_s0[91]), .Q (signal_12273) ) ;
    buf_sca_clk cell_2384 ( .C (clk), .D (key_s1[91]), .Q (signal_12274) ) ;
    buf_sca_clk cell_2385 ( .C (clk), .D (key_s0[92]), .Q (signal_12275) ) ;
    buf_sca_clk cell_2386 ( .C (clk), .D (key_s1[92]), .Q (signal_12276) ) ;
    buf_sca_clk cell_2387 ( .C (clk), .D (key_s0[93]), .Q (signal_12277) ) ;
    buf_sca_clk cell_2388 ( .C (clk), .D (key_s1[93]), .Q (signal_12278) ) ;
    buf_sca_clk cell_2389 ( .C (clk), .D (key_s0[94]), .Q (signal_12279) ) ;
    buf_sca_clk cell_2390 ( .C (clk), .D (key_s1[94]), .Q (signal_12280) ) ;
    buf_sca_clk cell_2391 ( .C (clk), .D (key_s0[95]), .Q (signal_12281) ) ;
    buf_sca_clk cell_2392 ( .C (clk), .D (key_s1[95]), .Q (signal_12282) ) ;
    buf_sca_clk cell_2393 ( .C (clk), .D (key_s0[96]), .Q (signal_12283) ) ;
    buf_sca_clk cell_2394 ( .C (clk), .D (key_s1[96]), .Q (signal_12284) ) ;
    buf_sca_clk cell_2395 ( .C (clk), .D (key_s0[97]), .Q (signal_12285) ) ;
    buf_sca_clk cell_2396 ( .C (clk), .D (key_s1[97]), .Q (signal_12286) ) ;
    buf_sca_clk cell_2397 ( .C (clk), .D (key_s0[98]), .Q (signal_12287) ) ;
    buf_sca_clk cell_2398 ( .C (clk), .D (key_s1[98]), .Q (signal_12288) ) ;
    buf_sca_clk cell_2399 ( .C (clk), .D (key_s0[99]), .Q (signal_12289) ) ;
    buf_sca_clk cell_2400 ( .C (clk), .D (key_s1[99]), .Q (signal_12290) ) ;
    buf_sca_clk cell_2401 ( .C (clk), .D (key_s0[100]), .Q (signal_12291) ) ;
    buf_sca_clk cell_2402 ( .C (clk), .D (key_s1[100]), .Q (signal_12292) ) ;
    buf_sca_clk cell_2403 ( .C (clk), .D (key_s0[101]), .Q (signal_12293) ) ;
    buf_sca_clk cell_2404 ( .C (clk), .D (key_s1[101]), .Q (signal_12294) ) ;
    buf_sca_clk cell_2405 ( .C (clk), .D (key_s0[102]), .Q (signal_12295) ) ;
    buf_sca_clk cell_2406 ( .C (clk), .D (key_s1[102]), .Q (signal_12296) ) ;
    buf_sca_clk cell_2407 ( .C (clk), .D (key_s0[103]), .Q (signal_12297) ) ;
    buf_sca_clk cell_2408 ( .C (clk), .D (key_s1[103]), .Q (signal_12298) ) ;
    buf_sca_clk cell_2409 ( .C (clk), .D (key_s0[104]), .Q (signal_12299) ) ;
    buf_sca_clk cell_2410 ( .C (clk), .D (key_s1[104]), .Q (signal_12300) ) ;
    buf_sca_clk cell_2411 ( .C (clk), .D (key_s0[105]), .Q (signal_12301) ) ;
    buf_sca_clk cell_2412 ( .C (clk), .D (key_s1[105]), .Q (signal_12302) ) ;
    buf_sca_clk cell_2413 ( .C (clk), .D (key_s0[106]), .Q (signal_12303) ) ;
    buf_sca_clk cell_2414 ( .C (clk), .D (key_s1[106]), .Q (signal_12304) ) ;
    buf_sca_clk cell_2415 ( .C (clk), .D (key_s0[107]), .Q (signal_12305) ) ;
    buf_sca_clk cell_2416 ( .C (clk), .D (key_s1[107]), .Q (signal_12306) ) ;
    buf_sca_clk cell_2417 ( .C (clk), .D (key_s0[108]), .Q (signal_12307) ) ;
    buf_sca_clk cell_2418 ( .C (clk), .D (key_s1[108]), .Q (signal_12308) ) ;
    buf_sca_clk cell_2419 ( .C (clk), .D (key_s0[109]), .Q (signal_12309) ) ;
    buf_sca_clk cell_2420 ( .C (clk), .D (key_s1[109]), .Q (signal_12310) ) ;
    buf_sca_clk cell_2421 ( .C (clk), .D (key_s0[110]), .Q (signal_12311) ) ;
    buf_sca_clk cell_2422 ( .C (clk), .D (key_s1[110]), .Q (signal_12312) ) ;
    buf_sca_clk cell_2423 ( .C (clk), .D (key_s0[111]), .Q (signal_12313) ) ;
    buf_sca_clk cell_2424 ( .C (clk), .D (key_s1[111]), .Q (signal_12314) ) ;
    buf_sca_clk cell_2425 ( .C (clk), .D (key_s0[112]), .Q (signal_12315) ) ;
    buf_sca_clk cell_2426 ( .C (clk), .D (key_s1[112]), .Q (signal_12316) ) ;
    buf_sca_clk cell_2427 ( .C (clk), .D (key_s0[113]), .Q (signal_12317) ) ;
    buf_sca_clk cell_2428 ( .C (clk), .D (key_s1[113]), .Q (signal_12318) ) ;
    buf_sca_clk cell_2429 ( .C (clk), .D (key_s0[114]), .Q (signal_12319) ) ;
    buf_sca_clk cell_2430 ( .C (clk), .D (key_s1[114]), .Q (signal_12320) ) ;
    buf_sca_clk cell_2431 ( .C (clk), .D (key_s0[115]), .Q (signal_12321) ) ;
    buf_sca_clk cell_2432 ( .C (clk), .D (key_s1[115]), .Q (signal_12322) ) ;
    buf_sca_clk cell_2433 ( .C (clk), .D (key_s0[116]), .Q (signal_12323) ) ;
    buf_sca_clk cell_2434 ( .C (clk), .D (key_s1[116]), .Q (signal_12324) ) ;
    buf_sca_clk cell_2435 ( .C (clk), .D (key_s0[117]), .Q (signal_12325) ) ;
    buf_sca_clk cell_2436 ( .C (clk), .D (key_s1[117]), .Q (signal_12326) ) ;
    buf_sca_clk cell_2437 ( .C (clk), .D (key_s0[118]), .Q (signal_12327) ) ;
    buf_sca_clk cell_2438 ( .C (clk), .D (key_s1[118]), .Q (signal_12328) ) ;
    buf_sca_clk cell_2439 ( .C (clk), .D (key_s0[119]), .Q (signal_12329) ) ;
    buf_sca_clk cell_2440 ( .C (clk), .D (key_s1[119]), .Q (signal_12330) ) ;
    buf_sca_clk cell_2441 ( .C (clk), .D (key_s0[120]), .Q (signal_12331) ) ;
    buf_sca_clk cell_2442 ( .C (clk), .D (key_s1[120]), .Q (signal_12332) ) ;
    buf_sca_clk cell_2443 ( .C (clk), .D (key_s0[121]), .Q (signal_12333) ) ;
    buf_sca_clk cell_2444 ( .C (clk), .D (key_s1[121]), .Q (signal_12334) ) ;
    buf_sca_clk cell_2445 ( .C (clk), .D (key_s0[122]), .Q (signal_12335) ) ;
    buf_sca_clk cell_2446 ( .C (clk), .D (key_s1[122]), .Q (signal_12336) ) ;
    buf_sca_clk cell_2447 ( .C (clk), .D (key_s0[123]), .Q (signal_12337) ) ;
    buf_sca_clk cell_2448 ( .C (clk), .D (key_s1[123]), .Q (signal_12338) ) ;
    buf_sca_clk cell_2449 ( .C (clk), .D (key_s0[124]), .Q (signal_12339) ) ;
    buf_sca_clk cell_2450 ( .C (clk), .D (key_s1[124]), .Q (signal_12340) ) ;
    buf_sca_clk cell_2451 ( .C (clk), .D (key_s0[125]), .Q (signal_12341) ) ;
    buf_sca_clk cell_2452 ( .C (clk), .D (key_s1[125]), .Q (signal_12342) ) ;
    buf_sca_clk cell_2453 ( .C (clk), .D (key_s0[126]), .Q (signal_12343) ) ;
    buf_sca_clk cell_2454 ( .C (clk), .D (key_s1[126]), .Q (signal_12344) ) ;
    buf_sca_clk cell_2455 ( .C (clk), .D (key_s0[127]), .Q (signal_12345) ) ;
    buf_sca_clk cell_2456 ( .C (clk), .D (key_s1[127]), .Q (signal_12346) ) ;
    buf_sca_clk cell_2457 ( .C (clk), .D (signal_1800), .Q (signal_12347) ) ;
    buf_sca_clk cell_2458 ( .C (clk), .D (signal_2720), .Q (signal_12348) ) ;
    buf_sca_clk cell_2459 ( .C (clk), .D (signal_1801), .Q (signal_12349) ) ;
    buf_sca_clk cell_2460 ( .C (clk), .D (signal_2687), .Q (signal_12350) ) ;
    buf_sca_clk cell_2461 ( .C (clk), .D (signal_1786), .Q (signal_12351) ) ;
    buf_sca_clk cell_2462 ( .C (clk), .D (signal_2654), .Q (signal_12352) ) ;
    buf_sca_clk cell_2463 ( .C (clk), .D (signal_1787), .Q (signal_12353) ) ;
    buf_sca_clk cell_2464 ( .C (clk), .D (signal_2621), .Q (signal_12354) ) ;
    buf_sca_clk cell_2465 ( .C (clk), .D (signal_1788), .Q (signal_12355) ) ;
    buf_sca_clk cell_2466 ( .C (clk), .D (signal_2588), .Q (signal_12356) ) ;
    buf_sca_clk cell_2467 ( .C (clk), .D (signal_1789), .Q (signal_12357) ) ;
    buf_sca_clk cell_2468 ( .C (clk), .D (signal_2555), .Q (signal_12358) ) ;
    buf_sca_clk cell_2469 ( .C (clk), .D (signal_2124), .Q (signal_12359) ) ;
    buf_sca_clk cell_2470 ( .C (clk), .D (signal_2528), .Q (signal_12360) ) ;
    buf_sca_clk cell_2471 ( .C (clk), .D (signal_2092), .Q (signal_12361) ) ;
    buf_sca_clk cell_2472 ( .C (clk), .D (signal_2633), .Q (signal_12362) ) ;
    buf_sca_clk cell_2473 ( .C (clk), .D (signal_2125), .Q (signal_12363) ) ;
    buf_sca_clk cell_2474 ( .C (clk), .D (signal_2525), .Q (signal_12364) ) ;
    buf_sca_clk cell_2475 ( .C (clk), .D (signal_2093), .Q (signal_12365) ) ;
    buf_sca_clk cell_2476 ( .C (clk), .D (signal_2630), .Q (signal_12366) ) ;
    buf_sca_clk cell_2477 ( .C (clk), .D (signal_1790), .Q (signal_12367) ) ;
    buf_sca_clk cell_2478 ( .C (clk), .D (signal_2522), .Q (signal_12368) ) ;
    buf_sca_clk cell_2479 ( .C (clk), .D (signal_2126), .Q (signal_12369) ) ;
    buf_sca_clk cell_2480 ( .C (clk), .D (signal_2519), .Q (signal_12370) ) ;
    buf_sca_clk cell_2481 ( .C (clk), .D (signal_2094), .Q (signal_12371) ) ;
    buf_sca_clk cell_2482 ( .C (clk), .D (signal_2627), .Q (signal_12372) ) ;
    buf_sca_clk cell_2483 ( .C (clk), .D (signal_2127), .Q (signal_12373) ) ;
    buf_sca_clk cell_2484 ( .C (clk), .D (signal_2516), .Q (signal_12374) ) ;
    buf_sca_clk cell_2485 ( .C (clk), .D (signal_2095), .Q (signal_12375) ) ;
    buf_sca_clk cell_2486 ( .C (clk), .D (signal_2624), .Q (signal_12376) ) ;
    buf_sca_clk cell_2487 ( .C (clk), .D (signal_2128), .Q (signal_12377) ) ;
    buf_sca_clk cell_2488 ( .C (clk), .D (signal_2513), .Q (signal_12378) ) ;
    buf_sca_clk cell_2489 ( .C (clk), .D (signal_2096), .Q (signal_12379) ) ;
    buf_sca_clk cell_2490 ( .C (clk), .D (signal_2618), .Q (signal_12380) ) ;
    buf_sca_clk cell_2491 ( .C (clk), .D (signal_2129), .Q (signal_12381) ) ;
    buf_sca_clk cell_2492 ( .C (clk), .D (signal_2510), .Q (signal_12382) ) ;
    buf_sca_clk cell_2493 ( .C (clk), .D (signal_2097), .Q (signal_12383) ) ;
    buf_sca_clk cell_2494 ( .C (clk), .D (signal_2615), .Q (signal_12384) ) ;
    buf_sca_clk cell_2495 ( .C (clk), .D (signal_2130), .Q (signal_12385) ) ;
    buf_sca_clk cell_2496 ( .C (clk), .D (signal_2507), .Q (signal_12386) ) ;
    buf_sca_clk cell_2497 ( .C (clk), .D (signal_2098), .Q (signal_12387) ) ;
    buf_sca_clk cell_2498 ( .C (clk), .D (signal_2612), .Q (signal_12388) ) ;
    buf_sca_clk cell_2499 ( .C (clk), .D (signal_2066), .Q (signal_12389) ) ;
    buf_sca_clk cell_2500 ( .C (clk), .D (signal_2717), .Q (signal_12390) ) ;
    buf_sca_clk cell_2501 ( .C (clk), .D (signal_1778), .Q (signal_12391) ) ;
    buf_sca_clk cell_2502 ( .C (clk), .D (signal_2495), .Q (signal_12392) ) ;
    buf_sca_clk cell_2503 ( .C (clk), .D (signal_2102), .Q (signal_12393) ) ;
    buf_sca_clk cell_2504 ( .C (clk), .D (signal_2600), .Q (signal_12394) ) ;
    buf_sca_clk cell_2505 ( .C (clk), .D (signal_2070), .Q (signal_12395) ) ;
    buf_sca_clk cell_2506 ( .C (clk), .D (signal_2705), .Q (signal_12396) ) ;
    buf_sca_clk cell_2507 ( .C (clk), .D (signal_1779), .Q (signal_12397) ) ;
    buf_sca_clk cell_2508 ( .C (clk), .D (signal_2492), .Q (signal_12398) ) ;
    buf_sca_clk cell_2509 ( .C (clk), .D (signal_2103), .Q (signal_12399) ) ;
    buf_sca_clk cell_2510 ( .C (clk), .D (signal_2597), .Q (signal_12400) ) ;
    buf_sca_clk cell_2511 ( .C (clk), .D (signal_2071), .Q (signal_12401) ) ;
    buf_sca_clk cell_2512 ( .C (clk), .D (signal_2702), .Q (signal_12402) ) ;
    buf_sca_clk cell_2513 ( .C (clk), .D (signal_1791), .Q (signal_12403) ) ;
    buf_sca_clk cell_2514 ( .C (clk), .D (signal_2489), .Q (signal_12404) ) ;
    buf_sca_clk cell_2515 ( .C (clk), .D (signal_2131), .Q (signal_12405) ) ;
    buf_sca_clk cell_2516 ( .C (clk), .D (signal_2504), .Q (signal_12406) ) ;
    buf_sca_clk cell_2517 ( .C (clk), .D (signal_2099), .Q (signal_12407) ) ;
    buf_sca_clk cell_2518 ( .C (clk), .D (signal_2609), .Q (signal_12408) ) ;
    buf_sca_clk cell_2519 ( .C (clk), .D (signal_2067), .Q (signal_12409) ) ;
    buf_sca_clk cell_2520 ( .C (clk), .D (signal_2714), .Q (signal_12410) ) ;
    buf_sca_clk cell_2521 ( .C (clk), .D (signal_1780), .Q (signal_12411) ) ;
    buf_sca_clk cell_2522 ( .C (clk), .D (signal_2486), .Q (signal_12412) ) ;
    buf_sca_clk cell_2523 ( .C (clk), .D (signal_2104), .Q (signal_12413) ) ;
    buf_sca_clk cell_2524 ( .C (clk), .D (signal_2594), .Q (signal_12414) ) ;
    buf_sca_clk cell_2525 ( .C (clk), .D (signal_2072), .Q (signal_12415) ) ;
    buf_sca_clk cell_2526 ( .C (clk), .D (signal_2699), .Q (signal_12416) ) ;
    buf_sca_clk cell_2527 ( .C (clk), .D (signal_1781), .Q (signal_12417) ) ;
    buf_sca_clk cell_2528 ( .C (clk), .D (signal_2483), .Q (signal_12418) ) ;
    buf_sca_clk cell_2529 ( .C (clk), .D (signal_2105), .Q (signal_12419) ) ;
    buf_sca_clk cell_2530 ( .C (clk), .D (signal_2591), .Q (signal_12420) ) ;
    buf_sca_clk cell_2531 ( .C (clk), .D (signal_2073), .Q (signal_12421) ) ;
    buf_sca_clk cell_2532 ( .C (clk), .D (signal_2696), .Q (signal_12422) ) ;
    buf_sca_clk cell_2533 ( .C (clk), .D (signal_1782), .Q (signal_12423) ) ;
    buf_sca_clk cell_2534 ( .C (clk), .D (signal_2480), .Q (signal_12424) ) ;
    buf_sca_clk cell_2535 ( .C (clk), .D (signal_2106), .Q (signal_12425) ) ;
    buf_sca_clk cell_2536 ( .C (clk), .D (signal_2585), .Q (signal_12426) ) ;
    buf_sca_clk cell_2537 ( .C (clk), .D (signal_2074), .Q (signal_12427) ) ;
    buf_sca_clk cell_2538 ( .C (clk), .D (signal_2693), .Q (signal_12428) ) ;
    buf_sca_clk cell_2539 ( .C (clk), .D (signal_1783), .Q (signal_12429) ) ;
    buf_sca_clk cell_2540 ( .C (clk), .D (signal_2477), .Q (signal_12430) ) ;
    buf_sca_clk cell_2541 ( .C (clk), .D (signal_2107), .Q (signal_12431) ) ;
    buf_sca_clk cell_2542 ( .C (clk), .D (signal_2582), .Q (signal_12432) ) ;
    buf_sca_clk cell_2543 ( .C (clk), .D (signal_2075), .Q (signal_12433) ) ;
    buf_sca_clk cell_2544 ( .C (clk), .D (signal_2690), .Q (signal_12434) ) ;
    buf_sca_clk cell_2545 ( .C (clk), .D (signal_1784), .Q (signal_12435) ) ;
    buf_sca_clk cell_2546 ( .C (clk), .D (signal_2474), .Q (signal_12436) ) ;
    buf_sca_clk cell_2547 ( .C (clk), .D (signal_2108), .Q (signal_12437) ) ;
    buf_sca_clk cell_2548 ( .C (clk), .D (signal_2579), .Q (signal_12438) ) ;
    buf_sca_clk cell_2549 ( .C (clk), .D (signal_2076), .Q (signal_12439) ) ;
    buf_sca_clk cell_2550 ( .C (clk), .D (signal_2684), .Q (signal_12440) ) ;
    buf_sca_clk cell_2551 ( .C (clk), .D (signal_1785), .Q (signal_12441) ) ;
    buf_sca_clk cell_2552 ( .C (clk), .D (signal_2471), .Q (signal_12442) ) ;
    buf_sca_clk cell_2553 ( .C (clk), .D (signal_2109), .Q (signal_12443) ) ;
    buf_sca_clk cell_2554 ( .C (clk), .D (signal_2576), .Q (signal_12444) ) ;
    buf_sca_clk cell_2555 ( .C (clk), .D (signal_2077), .Q (signal_12445) ) ;
    buf_sca_clk cell_2556 ( .C (clk), .D (signal_2681), .Q (signal_12446) ) ;
    buf_sca_clk cell_2557 ( .C (clk), .D (signal_1802), .Q (signal_12447) ) ;
    buf_sca_clk cell_2558 ( .C (clk), .D (signal_2468), .Q (signal_12448) ) ;
    buf_sca_clk cell_2559 ( .C (clk), .D (signal_2110), .Q (signal_12449) ) ;
    buf_sca_clk cell_2560 ( .C (clk), .D (signal_2573), .Q (signal_12450) ) ;
    buf_sca_clk cell_2561 ( .C (clk), .D (signal_2078), .Q (signal_12451) ) ;
    buf_sca_clk cell_2562 ( .C (clk), .D (signal_2678), .Q (signal_12452) ) ;
    buf_sca_clk cell_2563 ( .C (clk), .D (signal_1803), .Q (signal_12453) ) ;
    buf_sca_clk cell_2564 ( .C (clk), .D (signal_2465), .Q (signal_12454) ) ;
    buf_sca_clk cell_2565 ( .C (clk), .D (signal_2111), .Q (signal_12455) ) ;
    buf_sca_clk cell_2566 ( .C (clk), .D (signal_2570), .Q (signal_12456) ) ;
    buf_sca_clk cell_2567 ( .C (clk), .D (signal_2079), .Q (signal_12457) ) ;
    buf_sca_clk cell_2568 ( .C (clk), .D (signal_2675), .Q (signal_12458) ) ;
    buf_sca_clk cell_2569 ( .C (clk), .D (signal_1804), .Q (signal_12459) ) ;
    buf_sca_clk cell_2570 ( .C (clk), .D (signal_2462), .Q (signal_12460) ) ;
    buf_sca_clk cell_2571 ( .C (clk), .D (signal_2112), .Q (signal_12461) ) ;
    buf_sca_clk cell_2572 ( .C (clk), .D (signal_2567), .Q (signal_12462) ) ;
    buf_sca_clk cell_2573 ( .C (clk), .D (signal_2080), .Q (signal_12463) ) ;
    buf_sca_clk cell_2574 ( .C (clk), .D (signal_2672), .Q (signal_12464) ) ;
    buf_sca_clk cell_2575 ( .C (clk), .D (signal_1805), .Q (signal_12465) ) ;
    buf_sca_clk cell_2576 ( .C (clk), .D (signal_2459), .Q (signal_12466) ) ;
    buf_sca_clk cell_2577 ( .C (clk), .D (signal_2113), .Q (signal_12467) ) ;
    buf_sca_clk cell_2578 ( .C (clk), .D (signal_2564), .Q (signal_12468) ) ;
    buf_sca_clk cell_2579 ( .C (clk), .D (signal_2081), .Q (signal_12469) ) ;
    buf_sca_clk cell_2580 ( .C (clk), .D (signal_2669), .Q (signal_12470) ) ;
    buf_sca_clk cell_2581 ( .C (clk), .D (signal_1792), .Q (signal_12471) ) ;
    buf_sca_clk cell_2582 ( .C (clk), .D (signal_2456), .Q (signal_12472) ) ;
    buf_sca_clk cell_2583 ( .C (clk), .D (signal_2132), .Q (signal_12473) ) ;
    buf_sca_clk cell_2584 ( .C (clk), .D (signal_2501), .Q (signal_12474) ) ;
    buf_sca_clk cell_2585 ( .C (clk), .D (signal_2100), .Q (signal_12475) ) ;
    buf_sca_clk cell_2586 ( .C (clk), .D (signal_2606), .Q (signal_12476) ) ;
    buf_sca_clk cell_2587 ( .C (clk), .D (signal_2068), .Q (signal_12477) ) ;
    buf_sca_clk cell_2588 ( .C (clk), .D (signal_2711), .Q (signal_12478) ) ;
    buf_sca_clk cell_2589 ( .C (clk), .D (signal_1806), .Q (signal_12479) ) ;
    buf_sca_clk cell_2590 ( .C (clk), .D (signal_2453), .Q (signal_12480) ) ;
    buf_sca_clk cell_2591 ( .C (clk), .D (signal_2114), .Q (signal_12481) ) ;
    buf_sca_clk cell_2592 ( .C (clk), .D (signal_2561), .Q (signal_12482) ) ;
    buf_sca_clk cell_2593 ( .C (clk), .D (signal_2082), .Q (signal_12483) ) ;
    buf_sca_clk cell_2594 ( .C (clk), .D (signal_2666), .Q (signal_12484) ) ;
    buf_sca_clk cell_2595 ( .C (clk), .D (signal_1807), .Q (signal_12485) ) ;
    buf_sca_clk cell_2596 ( .C (clk), .D (signal_2450), .Q (signal_12486) ) ;
    buf_sca_clk cell_2597 ( .C (clk), .D (signal_2115), .Q (signal_12487) ) ;
    buf_sca_clk cell_2598 ( .C (clk), .D (signal_2558), .Q (signal_12488) ) ;
    buf_sca_clk cell_2599 ( .C (clk), .D (signal_2083), .Q (signal_12489) ) ;
    buf_sca_clk cell_2600 ( .C (clk), .D (signal_2663), .Q (signal_12490) ) ;
    buf_sca_clk cell_2601 ( .C (clk), .D (signal_1808), .Q (signal_12491) ) ;
    buf_sca_clk cell_2602 ( .C (clk), .D (signal_2447), .Q (signal_12492) ) ;
    buf_sca_clk cell_2603 ( .C (clk), .D (signal_2116), .Q (signal_12493) ) ;
    buf_sca_clk cell_2604 ( .C (clk), .D (signal_2552), .Q (signal_12494) ) ;
    buf_sca_clk cell_2605 ( .C (clk), .D (signal_2084), .Q (signal_12495) ) ;
    buf_sca_clk cell_2606 ( .C (clk), .D (signal_2660), .Q (signal_12496) ) ;
    buf_sca_clk cell_2607 ( .C (clk), .D (signal_1809), .Q (signal_12497) ) ;
    buf_sca_clk cell_2608 ( .C (clk), .D (signal_2444), .Q (signal_12498) ) ;
    buf_sca_clk cell_2609 ( .C (clk), .D (signal_2117), .Q (signal_12499) ) ;
    buf_sca_clk cell_2610 ( .C (clk), .D (signal_2549), .Q (signal_12500) ) ;
    buf_sca_clk cell_2611 ( .C (clk), .D (signal_2085), .Q (signal_12501) ) ;
    buf_sca_clk cell_2612 ( .C (clk), .D (signal_2657), .Q (signal_12502) ) ;
    buf_sca_clk cell_2613 ( .C (clk), .D (signal_1794), .Q (signal_12503) ) ;
    buf_sca_clk cell_2614 ( .C (clk), .D (signal_2441), .Q (signal_12504) ) ;
    buf_sca_clk cell_2615 ( .C (clk), .D (signal_2118), .Q (signal_12505) ) ;
    buf_sca_clk cell_2616 ( .C (clk), .D (signal_2546), .Q (signal_12506) ) ;
    buf_sca_clk cell_2617 ( .C (clk), .D (signal_2086), .Q (signal_12507) ) ;
    buf_sca_clk cell_2618 ( .C (clk), .D (signal_2651), .Q (signal_12508) ) ;
    buf_sca_clk cell_2619 ( .C (clk), .D (signal_1795), .Q (signal_12509) ) ;
    buf_sca_clk cell_2620 ( .C (clk), .D (signal_2438), .Q (signal_12510) ) ;
    buf_sca_clk cell_2621 ( .C (clk), .D (signal_2119), .Q (signal_12511) ) ;
    buf_sca_clk cell_2622 ( .C (clk), .D (signal_2543), .Q (signal_12512) ) ;
    buf_sca_clk cell_2623 ( .C (clk), .D (signal_2087), .Q (signal_12513) ) ;
    buf_sca_clk cell_2624 ( .C (clk), .D (signal_2648), .Q (signal_12514) ) ;
    buf_sca_clk cell_2625 ( .C (clk), .D (signal_1796), .Q (signal_12515) ) ;
    buf_sca_clk cell_2626 ( .C (clk), .D (signal_2435), .Q (signal_12516) ) ;
    buf_sca_clk cell_2627 ( .C (clk), .D (signal_2120), .Q (signal_12517) ) ;
    buf_sca_clk cell_2628 ( .C (clk), .D (signal_2540), .Q (signal_12518) ) ;
    buf_sca_clk cell_2629 ( .C (clk), .D (signal_2088), .Q (signal_12519) ) ;
    buf_sca_clk cell_2630 ( .C (clk), .D (signal_2645), .Q (signal_12520) ) ;
    buf_sca_clk cell_2631 ( .C (clk), .D (signal_1797), .Q (signal_12521) ) ;
    buf_sca_clk cell_2632 ( .C (clk), .D (signal_2432), .Q (signal_12522) ) ;
    buf_sca_clk cell_2633 ( .C (clk), .D (signal_2121), .Q (signal_12523) ) ;
    buf_sca_clk cell_2634 ( .C (clk), .D (signal_2537), .Q (signal_12524) ) ;
    buf_sca_clk cell_2635 ( .C (clk), .D (signal_2089), .Q (signal_12525) ) ;
    buf_sca_clk cell_2636 ( .C (clk), .D (signal_2642), .Q (signal_12526) ) ;
    buf_sca_clk cell_2637 ( .C (clk), .D (signal_2038), .Q (signal_12527) ) ;
    buf_sca_clk cell_2638 ( .C (clk), .D (signal_2429), .Q (signal_12528) ) ;
    buf_sca_clk cell_2639 ( .C (clk), .D (signal_2039), .Q (signal_12529) ) ;
    buf_sca_clk cell_2640 ( .C (clk), .D (signal_2426), .Q (signal_12530) ) ;
    buf_sca_clk cell_2641 ( .C (clk), .D (signal_2040), .Q (signal_12531) ) ;
    buf_sca_clk cell_2642 ( .C (clk), .D (signal_2423), .Q (signal_12532) ) ;
    buf_sca_clk cell_2643 ( .C (clk), .D (signal_2041), .Q (signal_12533) ) ;
    buf_sca_clk cell_2644 ( .C (clk), .D (signal_2420), .Q (signal_12534) ) ;
    buf_sca_clk cell_2645 ( .C (clk), .D (signal_2042), .Q (signal_12535) ) ;
    buf_sca_clk cell_2646 ( .C (clk), .D (signal_2417), .Q (signal_12536) ) ;
    buf_sca_clk cell_2647 ( .C (clk), .D (signal_2043), .Q (signal_12537) ) ;
    buf_sca_clk cell_2648 ( .C (clk), .D (signal_2414), .Q (signal_12538) ) ;
    buf_sca_clk cell_2649 ( .C (clk), .D (signal_2044), .Q (signal_12539) ) ;
    buf_sca_clk cell_2650 ( .C (clk), .D (signal_2411), .Q (signal_12540) ) ;
    buf_sca_clk cell_2651 ( .C (clk), .D (signal_2045), .Q (signal_12541) ) ;
    buf_sca_clk cell_2652 ( .C (clk), .D (signal_2408), .Q (signal_12542) ) ;
    buf_sca_clk cell_2653 ( .C (clk), .D (signal_1798), .Q (signal_12543) ) ;
    buf_sca_clk cell_2654 ( .C (clk), .D (signal_2405), .Q (signal_12544) ) ;
    buf_sca_clk cell_2655 ( .C (clk), .D (signal_2122), .Q (signal_12545) ) ;
    buf_sca_clk cell_2656 ( .C (clk), .D (signal_2534), .Q (signal_12546) ) ;
    buf_sca_clk cell_2657 ( .C (clk), .D (signal_2090), .Q (signal_12547) ) ;
    buf_sca_clk cell_2658 ( .C (clk), .D (signal_2639), .Q (signal_12548) ) ;
    buf_sca_clk cell_2659 ( .C (clk), .D (signal_2046), .Q (signal_12549) ) ;
    buf_sca_clk cell_2660 ( .C (clk), .D (signal_2402), .Q (signal_12550) ) ;
    buf_sca_clk cell_2661 ( .C (clk), .D (signal_2047), .Q (signal_12551) ) ;
    buf_sca_clk cell_2662 ( .C (clk), .D (signal_2399), .Q (signal_12552) ) ;
    buf_sca_clk cell_2663 ( .C (clk), .D (signal_2048), .Q (signal_12553) ) ;
    buf_sca_clk cell_2664 ( .C (clk), .D (signal_2396), .Q (signal_12554) ) ;
    buf_sca_clk cell_2665 ( .C (clk), .D (signal_2049), .Q (signal_12555) ) ;
    buf_sca_clk cell_2666 ( .C (clk), .D (signal_2393), .Q (signal_12556) ) ;
    buf_sca_clk cell_2667 ( .C (clk), .D (signal_2050), .Q (signal_12557) ) ;
    buf_sca_clk cell_2668 ( .C (clk), .D (signal_2390), .Q (signal_12558) ) ;
    buf_sca_clk cell_2669 ( .C (clk), .D (signal_2051), .Q (signal_12559) ) ;
    buf_sca_clk cell_2670 ( .C (clk), .D (signal_2387), .Q (signal_12560) ) ;
    buf_sca_clk cell_2671 ( .C (clk), .D (signal_2052), .Q (signal_12561) ) ;
    buf_sca_clk cell_2672 ( .C (clk), .D (signal_2384), .Q (signal_12562) ) ;
    buf_sca_clk cell_2673 ( .C (clk), .D (signal_2053), .Q (signal_12563) ) ;
    buf_sca_clk cell_2674 ( .C (clk), .D (signal_2381), .Q (signal_12564) ) ;
    buf_sca_clk cell_2675 ( .C (clk), .D (signal_2054), .Q (signal_12565) ) ;
    buf_sca_clk cell_2676 ( .C (clk), .D (signal_2378), .Q (signal_12566) ) ;
    buf_sca_clk cell_2677 ( .C (clk), .D (signal_2055), .Q (signal_12567) ) ;
    buf_sca_clk cell_2678 ( .C (clk), .D (signal_2375), .Q (signal_12568) ) ;
    buf_sca_clk cell_2679 ( .C (clk), .D (signal_1799), .Q (signal_12569) ) ;
    buf_sca_clk cell_2680 ( .C (clk), .D (signal_2372), .Q (signal_12570) ) ;
    buf_sca_clk cell_2681 ( .C (clk), .D (signal_2123), .Q (signal_12571) ) ;
    buf_sca_clk cell_2682 ( .C (clk), .D (signal_2531), .Q (signal_12572) ) ;
    buf_sca_clk cell_2683 ( .C (clk), .D (signal_2091), .Q (signal_12573) ) ;
    buf_sca_clk cell_2684 ( .C (clk), .D (signal_2636), .Q (signal_12574) ) ;
    buf_sca_clk cell_2685 ( .C (clk), .D (signal_2056), .Q (signal_12575) ) ;
    buf_sca_clk cell_2686 ( .C (clk), .D (signal_2369), .Q (signal_12576) ) ;
    buf_sca_clk cell_2687 ( .C (clk), .D (signal_2057), .Q (signal_12577) ) ;
    buf_sca_clk cell_2688 ( .C (clk), .D (signal_2366), .Q (signal_12578) ) ;
    buf_sca_clk cell_2689 ( .C (clk), .D (signal_2058), .Q (signal_12579) ) ;
    buf_sca_clk cell_2690 ( .C (clk), .D (signal_2363), .Q (signal_12580) ) ;
    buf_sca_clk cell_2691 ( .C (clk), .D (signal_2059), .Q (signal_12581) ) ;
    buf_sca_clk cell_2692 ( .C (clk), .D (signal_2360), .Q (signal_12582) ) ;
    buf_sca_clk cell_2693 ( .C (clk), .D (signal_2060), .Q (signal_12583) ) ;
    buf_sca_clk cell_2694 ( .C (clk), .D (signal_2357), .Q (signal_12584) ) ;
    buf_sca_clk cell_2695 ( .C (clk), .D (signal_2061), .Q (signal_12585) ) ;
    buf_sca_clk cell_2696 ( .C (clk), .D (signal_2354), .Q (signal_12586) ) ;
    buf_sca_clk cell_2697 ( .C (clk), .D (signal_2062), .Q (signal_12587) ) ;
    buf_sca_clk cell_2698 ( .C (clk), .D (signal_2351), .Q (signal_12588) ) ;
    buf_sca_clk cell_2699 ( .C (clk), .D (signal_2063), .Q (signal_12589) ) ;
    buf_sca_clk cell_2700 ( .C (clk), .D (signal_2348), .Q (signal_12590) ) ;
    buf_sca_clk cell_2701 ( .C (clk), .D (signal_2064), .Q (signal_12591) ) ;
    buf_sca_clk cell_2702 ( .C (clk), .D (signal_2345), .Q (signal_12592) ) ;
    buf_sca_clk cell_2703 ( .C (clk), .D (signal_2065), .Q (signal_12593) ) ;
    buf_sca_clk cell_2704 ( .C (clk), .D (signal_2342), .Q (signal_12594) ) ;
    buf_sca_clk cell_2705 ( .C (clk), .D (signal_1793), .Q (signal_12595) ) ;
    buf_sca_clk cell_2706 ( .C (clk), .D (signal_2339), .Q (signal_12596) ) ;
    buf_sca_clk cell_2707 ( .C (clk), .D (signal_2133), .Q (signal_12597) ) ;
    buf_sca_clk cell_2708 ( .C (clk), .D (signal_2498), .Q (signal_12598) ) ;
    buf_sca_clk cell_2709 ( .C (clk), .D (signal_2101), .Q (signal_12599) ) ;
    buf_sca_clk cell_2710 ( .C (clk), .D (signal_2603), .Q (signal_12600) ) ;
    buf_sca_clk cell_2711 ( .C (clk), .D (signal_2069), .Q (signal_12601) ) ;
    buf_sca_clk cell_2712 ( .C (clk), .D (signal_2708), .Q (signal_12602) ) ;
    buf_clk cell_2713 ( .C (clk), .D (signal_2134), .Q (signal_12603) ) ;
    buf_clk cell_2714 ( .C (clk), .D (signal_2135), .Q (signal_12604) ) ;
    buf_clk cell_2715 ( .C (clk), .D (signal_2136), .Q (signal_12605) ) ;
    buf_clk cell_2716 ( .C (clk), .D (signal_2137), .Q (signal_12606) ) ;
    buf_clk cell_2717 ( .C (clk), .D (signal_2138), .Q (signal_12607) ) ;
    buf_clk cell_2718 ( .C (clk), .D (signal_2139), .Q (signal_12608) ) ;
    buf_clk cell_2719 ( .C (clk), .D (signal_2140), .Q (signal_12609) ) ;
    buf_clk cell_2720 ( .C (clk), .D (signal_2141), .Q (signal_12610) ) ;
    buf_clk cell_2721 ( .C (clk), .D (signal_1489), .Q (signal_12611) ) ;
    buf_clk cell_2722 ( .C (clk), .D (signal_1488), .Q (signal_12612) ) ;
    buf_clk cell_2723 ( .C (clk), .D (signal_1487), .Q (signal_12613) ) ;
    buf_clk cell_2724 ( .C (clk), .D (signal_1486), .Q (signal_12614) ) ;
    buf_clk cell_2725 ( .C (clk), .D (signal_1485), .Q (signal_12615) ) ;
    buf_clk cell_2726 ( .C (clk), .D (signal_1484), .Q (signal_12616) ) ;
    buf_clk cell_2727 ( .C (clk), .D (signal_1490), .Q (signal_12617) ) ;
    buf_sca_clk cell_2728 ( .C (clk), .D (signal_478), .Q (signal_12618) ) ;
    buf_sca_clk cell_2729 ( .C (clk), .D (signal_2851), .Q (signal_12619) ) ;
    buf_sca_clk cell_2730 ( .C (clk), .D (signal_480), .Q (signal_12620) ) ;
    buf_sca_clk cell_2731 ( .C (clk), .D (signal_2853), .Q (signal_12621) ) ;
    buf_sca_clk cell_2732 ( .C (clk), .D (signal_482), .Q (signal_12622) ) ;
    buf_sca_clk cell_2733 ( .C (clk), .D (signal_2855), .Q (signal_12623) ) ;
    buf_sca_clk cell_2734 ( .C (clk), .D (signal_484), .Q (signal_12624) ) ;
    buf_sca_clk cell_2735 ( .C (clk), .D (signal_2857), .Q (signal_12625) ) ;
    buf_sca_clk cell_2736 ( .C (clk), .D (signal_486), .Q (signal_12626) ) ;
    buf_sca_clk cell_2737 ( .C (clk), .D (signal_2859), .Q (signal_12627) ) ;
    buf_sca_clk cell_2738 ( .C (clk), .D (signal_488), .Q (signal_12628) ) ;
    buf_sca_clk cell_2739 ( .C (clk), .D (signal_2861), .Q (signal_12629) ) ;
    buf_sca_clk cell_2740 ( .C (clk), .D (signal_490), .Q (signal_12630) ) ;
    buf_sca_clk cell_2741 ( .C (clk), .D (signal_2863), .Q (signal_12631) ) ;
    buf_sca_clk cell_2742 ( .C (clk), .D (signal_492), .Q (signal_12632) ) ;
    buf_sca_clk cell_2743 ( .C (clk), .D (signal_2865), .Q (signal_12633) ) ;
    buf_sca_clk cell_2744 ( .C (clk), .D (signal_494), .Q (signal_12634) ) ;
    buf_sca_clk cell_2745 ( .C (clk), .D (signal_2867), .Q (signal_12635) ) ;
    buf_sca_clk cell_2746 ( .C (clk), .D (signal_496), .Q (signal_12636) ) ;
    buf_sca_clk cell_2747 ( .C (clk), .D (signal_2869), .Q (signal_12637) ) ;
    buf_sca_clk cell_2748 ( .C (clk), .D (signal_498), .Q (signal_12638) ) ;
    buf_sca_clk cell_2749 ( .C (clk), .D (signal_2871), .Q (signal_12639) ) ;
    buf_sca_clk cell_2750 ( .C (clk), .D (signal_500), .Q (signal_12640) ) ;
    buf_sca_clk cell_2751 ( .C (clk), .D (signal_2873), .Q (signal_12641) ) ;
    buf_sca_clk cell_2752 ( .C (clk), .D (signal_502), .Q (signal_12642) ) ;
    buf_sca_clk cell_2753 ( .C (clk), .D (signal_2875), .Q (signal_12643) ) ;
    buf_sca_clk cell_2754 ( .C (clk), .D (signal_504), .Q (signal_12644) ) ;
    buf_sca_clk cell_2755 ( .C (clk), .D (signal_2877), .Q (signal_12645) ) ;
    buf_sca_clk cell_2756 ( .C (clk), .D (signal_506), .Q (signal_12646) ) ;
    buf_sca_clk cell_2757 ( .C (clk), .D (signal_2879), .Q (signal_12647) ) ;
    buf_sca_clk cell_2758 ( .C (clk), .D (signal_508), .Q (signal_12648) ) ;
    buf_sca_clk cell_2759 ( .C (clk), .D (signal_2881), .Q (signal_12649) ) ;
    buf_sca_clk cell_2760 ( .C (clk), .D (signal_510), .Q (signal_12650) ) ;
    buf_sca_clk cell_2761 ( .C (clk), .D (signal_2883), .Q (signal_12651) ) ;
    buf_sca_clk cell_2762 ( .C (clk), .D (signal_512), .Q (signal_12652) ) ;
    buf_sca_clk cell_2763 ( .C (clk), .D (signal_2885), .Q (signal_12653) ) ;
    buf_sca_clk cell_2764 ( .C (clk), .D (signal_514), .Q (signal_12654) ) ;
    buf_sca_clk cell_2765 ( .C (clk), .D (signal_2887), .Q (signal_12655) ) ;
    buf_sca_clk cell_2766 ( .C (clk), .D (signal_516), .Q (signal_12656) ) ;
    buf_sca_clk cell_2767 ( .C (clk), .D (signal_2889), .Q (signal_12657) ) ;
    buf_sca_clk cell_2768 ( .C (clk), .D (signal_518), .Q (signal_12658) ) ;
    buf_sca_clk cell_2769 ( .C (clk), .D (signal_2891), .Q (signal_12659) ) ;
    buf_sca_clk cell_2770 ( .C (clk), .D (signal_520), .Q (signal_12660) ) ;
    buf_sca_clk cell_2771 ( .C (clk), .D (signal_2893), .Q (signal_12661) ) ;
    buf_sca_clk cell_2772 ( .C (clk), .D (signal_522), .Q (signal_12662) ) ;
    buf_sca_clk cell_2773 ( .C (clk), .D (signal_2895), .Q (signal_12663) ) ;
    buf_sca_clk cell_2774 ( .C (clk), .D (signal_524), .Q (signal_12664) ) ;
    buf_sca_clk cell_2775 ( .C (clk), .D (signal_2897), .Q (signal_12665) ) ;
    buf_sca_clk cell_2776 ( .C (clk), .D (signal_526), .Q (signal_12666) ) ;
    buf_sca_clk cell_2777 ( .C (clk), .D (signal_2899), .Q (signal_12667) ) ;
    buf_sca_clk cell_2778 ( .C (clk), .D (signal_528), .Q (signal_12668) ) ;
    buf_sca_clk cell_2779 ( .C (clk), .D (signal_2901), .Q (signal_12669) ) ;
    buf_sca_clk cell_2780 ( .C (clk), .D (signal_530), .Q (signal_12670) ) ;
    buf_sca_clk cell_2781 ( .C (clk), .D (signal_2903), .Q (signal_12671) ) ;
    buf_sca_clk cell_2782 ( .C (clk), .D (signal_532), .Q (signal_12672) ) ;
    buf_sca_clk cell_2783 ( .C (clk), .D (signal_2905), .Q (signal_12673) ) ;
    buf_sca_clk cell_2784 ( .C (clk), .D (signal_534), .Q (signal_12674) ) ;
    buf_sca_clk cell_2785 ( .C (clk), .D (signal_2907), .Q (signal_12675) ) ;
    buf_sca_clk cell_2786 ( .C (clk), .D (signal_536), .Q (signal_12676) ) ;
    buf_sca_clk cell_2787 ( .C (clk), .D (signal_2909), .Q (signal_12677) ) ;
    buf_sca_clk cell_2788 ( .C (clk), .D (signal_538), .Q (signal_12678) ) ;
    buf_sca_clk cell_2789 ( .C (clk), .D (signal_2911), .Q (signal_12679) ) ;
    buf_sca_clk cell_2790 ( .C (clk), .D (signal_540), .Q (signal_12680) ) ;
    buf_sca_clk cell_2791 ( .C (clk), .D (signal_2913), .Q (signal_12681) ) ;
    buf_sca_clk cell_2792 ( .C (clk), .D (signal_542), .Q (signal_12682) ) ;
    buf_sca_clk cell_2793 ( .C (clk), .D (signal_2915), .Q (signal_12683) ) ;
    buf_sca_clk cell_2794 ( .C (clk), .D (signal_544), .Q (signal_12684) ) ;
    buf_sca_clk cell_2795 ( .C (clk), .D (signal_2917), .Q (signal_12685) ) ;
    buf_sca_clk cell_2796 ( .C (clk), .D (signal_546), .Q (signal_12686) ) ;
    buf_sca_clk cell_2797 ( .C (clk), .D (signal_2919), .Q (signal_12687) ) ;
    buf_sca_clk cell_2798 ( .C (clk), .D (signal_548), .Q (signal_12688) ) ;
    buf_sca_clk cell_2799 ( .C (clk), .D (signal_2921), .Q (signal_12689) ) ;
    buf_sca_clk cell_2800 ( .C (clk), .D (signal_550), .Q (signal_12690) ) ;
    buf_sca_clk cell_2801 ( .C (clk), .D (signal_2923), .Q (signal_12691) ) ;
    buf_sca_clk cell_2802 ( .C (clk), .D (signal_552), .Q (signal_12692) ) ;
    buf_sca_clk cell_2803 ( .C (clk), .D (signal_2925), .Q (signal_12693) ) ;
    buf_sca_clk cell_2804 ( .C (clk), .D (signal_554), .Q (signal_12694) ) ;
    buf_sca_clk cell_2805 ( .C (clk), .D (signal_2927), .Q (signal_12695) ) ;
    buf_sca_clk cell_2806 ( .C (clk), .D (signal_556), .Q (signal_12696) ) ;
    buf_sca_clk cell_2807 ( .C (clk), .D (signal_2929), .Q (signal_12697) ) ;
    buf_sca_clk cell_2808 ( .C (clk), .D (signal_558), .Q (signal_12698) ) ;
    buf_sca_clk cell_2809 ( .C (clk), .D (signal_2931), .Q (signal_12699) ) ;
    buf_sca_clk cell_2810 ( .C (clk), .D (signal_560), .Q (signal_12700) ) ;
    buf_sca_clk cell_2811 ( .C (clk), .D (signal_2933), .Q (signal_12701) ) ;
    buf_sca_clk cell_2812 ( .C (clk), .D (signal_562), .Q (signal_12702) ) ;
    buf_sca_clk cell_2813 ( .C (clk), .D (signal_2935), .Q (signal_12703) ) ;
    buf_sca_clk cell_2814 ( .C (clk), .D (signal_564), .Q (signal_12704) ) ;
    buf_sca_clk cell_2815 ( .C (clk), .D (signal_2937), .Q (signal_12705) ) ;
    buf_sca_clk cell_2816 ( .C (clk), .D (signal_566), .Q (signal_12706) ) ;
    buf_sca_clk cell_2817 ( .C (clk), .D (signal_2939), .Q (signal_12707) ) ;
    buf_sca_clk cell_2818 ( .C (clk), .D (signal_568), .Q (signal_12708) ) ;
    buf_sca_clk cell_2819 ( .C (clk), .D (signal_2941), .Q (signal_12709) ) ;
    buf_sca_clk cell_2820 ( .C (clk), .D (signal_570), .Q (signal_12710) ) ;
    buf_sca_clk cell_2821 ( .C (clk), .D (signal_2943), .Q (signal_12711) ) ;
    buf_sca_clk cell_2822 ( .C (clk), .D (signal_572), .Q (signal_12712) ) ;
    buf_sca_clk cell_2823 ( .C (clk), .D (signal_2945), .Q (signal_12713) ) ;
    buf_sca_clk cell_2824 ( .C (clk), .D (signal_574), .Q (signal_12714) ) ;
    buf_sca_clk cell_2825 ( .C (clk), .D (signal_2947), .Q (signal_12715) ) ;
    buf_sca_clk cell_2826 ( .C (clk), .D (signal_576), .Q (signal_12716) ) ;
    buf_sca_clk cell_2827 ( .C (clk), .D (signal_2949), .Q (signal_12717) ) ;
    buf_sca_clk cell_2828 ( .C (clk), .D (signal_578), .Q (signal_12718) ) ;
    buf_sca_clk cell_2829 ( .C (clk), .D (signal_2951), .Q (signal_12719) ) ;
    buf_sca_clk cell_2830 ( .C (clk), .D (signal_580), .Q (signal_12720) ) ;
    buf_sca_clk cell_2831 ( .C (clk), .D (signal_2953), .Q (signal_12721) ) ;
    buf_sca_clk cell_2832 ( .C (clk), .D (signal_582), .Q (signal_12722) ) ;
    buf_sca_clk cell_2833 ( .C (clk), .D (signal_2955), .Q (signal_12723) ) ;
    buf_sca_clk cell_2834 ( .C (clk), .D (signal_584), .Q (signal_12724) ) ;
    buf_sca_clk cell_2835 ( .C (clk), .D (signal_2957), .Q (signal_12725) ) ;
    buf_sca_clk cell_2836 ( .C (clk), .D (signal_586), .Q (signal_12726) ) ;
    buf_sca_clk cell_2837 ( .C (clk), .D (signal_2959), .Q (signal_12727) ) ;
    buf_sca_clk cell_2838 ( .C (clk), .D (signal_588), .Q (signal_12728) ) ;
    buf_sca_clk cell_2839 ( .C (clk), .D (signal_2961), .Q (signal_12729) ) ;
    buf_sca_clk cell_2840 ( .C (clk), .D (signal_590), .Q (signal_12730) ) ;
    buf_sca_clk cell_2841 ( .C (clk), .D (signal_2963), .Q (signal_12731) ) ;
    buf_sca_clk cell_2842 ( .C (clk), .D (signal_592), .Q (signal_12732) ) ;
    buf_sca_clk cell_2843 ( .C (clk), .D (signal_2965), .Q (signal_12733) ) ;
    buf_sca_clk cell_2844 ( .C (clk), .D (signal_594), .Q (signal_12734) ) ;
    buf_sca_clk cell_2845 ( .C (clk), .D (signal_2967), .Q (signal_12735) ) ;
    buf_sca_clk cell_2846 ( .C (clk), .D (signal_596), .Q (signal_12736) ) ;
    buf_sca_clk cell_2847 ( .C (clk), .D (signal_2969), .Q (signal_12737) ) ;
    buf_sca_clk cell_2848 ( .C (clk), .D (signal_598), .Q (signal_12738) ) ;
    buf_sca_clk cell_2849 ( .C (clk), .D (signal_2971), .Q (signal_12739) ) ;
    buf_sca_clk cell_2850 ( .C (clk), .D (signal_600), .Q (signal_12740) ) ;
    buf_sca_clk cell_2851 ( .C (clk), .D (signal_2973), .Q (signal_12741) ) ;
    buf_sca_clk cell_2852 ( .C (clk), .D (signal_602), .Q (signal_12742) ) ;
    buf_sca_clk cell_2853 ( .C (clk), .D (signal_2975), .Q (signal_12743) ) ;
    buf_sca_clk cell_2854 ( .C (clk), .D (signal_604), .Q (signal_12744) ) ;
    buf_sca_clk cell_2855 ( .C (clk), .D (signal_2977), .Q (signal_12745) ) ;
    buf_sca_clk cell_2856 ( .C (clk), .D (signal_606), .Q (signal_12746) ) ;
    buf_sca_clk cell_2857 ( .C (clk), .D (signal_2979), .Q (signal_12747) ) ;
    buf_sca_clk cell_2858 ( .C (clk), .D (signal_608), .Q (signal_12748) ) ;
    buf_sca_clk cell_2859 ( .C (clk), .D (signal_2981), .Q (signal_12749) ) ;
    buf_sca_clk cell_2860 ( .C (clk), .D (signal_610), .Q (signal_12750) ) ;
    buf_sca_clk cell_2861 ( .C (clk), .D (signal_2983), .Q (signal_12751) ) ;
    buf_sca_clk cell_2862 ( .C (clk), .D (signal_612), .Q (signal_12752) ) ;
    buf_sca_clk cell_2863 ( .C (clk), .D (signal_2985), .Q (signal_12753) ) ;
    buf_sca_clk cell_2864 ( .C (clk), .D (signal_614), .Q (signal_12754) ) ;
    buf_sca_clk cell_2865 ( .C (clk), .D (signal_2987), .Q (signal_12755) ) ;
    buf_sca_clk cell_2866 ( .C (clk), .D (signal_616), .Q (signal_12756) ) ;
    buf_sca_clk cell_2867 ( .C (clk), .D (signal_2989), .Q (signal_12757) ) ;
    buf_sca_clk cell_2868 ( .C (clk), .D (signal_618), .Q (signal_12758) ) ;
    buf_sca_clk cell_2869 ( .C (clk), .D (signal_2991), .Q (signal_12759) ) ;
    buf_sca_clk cell_2870 ( .C (clk), .D (signal_620), .Q (signal_12760) ) ;
    buf_sca_clk cell_2871 ( .C (clk), .D (signal_2993), .Q (signal_12761) ) ;
    buf_sca_clk cell_2872 ( .C (clk), .D (signal_622), .Q (signal_12762) ) ;
    buf_sca_clk cell_2873 ( .C (clk), .D (signal_2995), .Q (signal_12763) ) ;
    buf_sca_clk cell_2874 ( .C (clk), .D (signal_624), .Q (signal_12764) ) ;
    buf_sca_clk cell_2875 ( .C (clk), .D (signal_2997), .Q (signal_12765) ) ;
    buf_sca_clk cell_2876 ( .C (clk), .D (signal_626), .Q (signal_12766) ) ;
    buf_sca_clk cell_2877 ( .C (clk), .D (signal_2999), .Q (signal_12767) ) ;
    buf_sca_clk cell_2878 ( .C (clk), .D (signal_628), .Q (signal_12768) ) ;
    buf_sca_clk cell_2879 ( .C (clk), .D (signal_3001), .Q (signal_12769) ) ;
    buf_sca_clk cell_2880 ( .C (clk), .D (signal_630), .Q (signal_12770) ) ;
    buf_sca_clk cell_2881 ( .C (clk), .D (signal_3003), .Q (signal_12771) ) ;
    buf_sca_clk cell_2882 ( .C (clk), .D (signal_632), .Q (signal_12772) ) ;
    buf_sca_clk cell_2883 ( .C (clk), .D (signal_3005), .Q (signal_12773) ) ;
    buf_sca_clk cell_2884 ( .C (clk), .D (signal_634), .Q (signal_12774) ) ;
    buf_sca_clk cell_2885 ( .C (clk), .D (signal_3007), .Q (signal_12775) ) ;
    buf_sca_clk cell_2886 ( .C (clk), .D (signal_636), .Q (signal_12776) ) ;
    buf_sca_clk cell_2887 ( .C (clk), .D (signal_3009), .Q (signal_12777) ) ;
    buf_sca_clk cell_2888 ( .C (clk), .D (signal_638), .Q (signal_12778) ) ;
    buf_sca_clk cell_2889 ( .C (clk), .D (signal_3011), .Q (signal_12779) ) ;
    buf_sca_clk cell_2890 ( .C (clk), .D (signal_640), .Q (signal_12780) ) ;
    buf_sca_clk cell_2891 ( .C (clk), .D (signal_3013), .Q (signal_12781) ) ;
    buf_sca_clk cell_2892 ( .C (clk), .D (signal_642), .Q (signal_12782) ) ;
    buf_sca_clk cell_2893 ( .C (clk), .D (signal_3015), .Q (signal_12783) ) ;
    buf_sca_clk cell_2894 ( .C (clk), .D (signal_644), .Q (signal_12784) ) ;
    buf_sca_clk cell_2895 ( .C (clk), .D (signal_3017), .Q (signal_12785) ) ;
    buf_sca_clk cell_2896 ( .C (clk), .D (signal_646), .Q (signal_12786) ) ;
    buf_sca_clk cell_2897 ( .C (clk), .D (signal_3019), .Q (signal_12787) ) ;
    buf_sca_clk cell_2898 ( .C (clk), .D (signal_648), .Q (signal_12788) ) ;
    buf_sca_clk cell_2899 ( .C (clk), .D (signal_3021), .Q (signal_12789) ) ;
    buf_sca_clk cell_2900 ( .C (clk), .D (signal_650), .Q (signal_12790) ) ;
    buf_sca_clk cell_2901 ( .C (clk), .D (signal_3023), .Q (signal_12791) ) ;
    buf_sca_clk cell_2902 ( .C (clk), .D (signal_652), .Q (signal_12792) ) ;
    buf_sca_clk cell_2903 ( .C (clk), .D (signal_3025), .Q (signal_12793) ) ;
    buf_sca_clk cell_2904 ( .C (clk), .D (signal_654), .Q (signal_12794) ) ;
    buf_sca_clk cell_2905 ( .C (clk), .D (signal_3027), .Q (signal_12795) ) ;
    buf_sca_clk cell_2906 ( .C (clk), .D (signal_656), .Q (signal_12796) ) ;
    buf_sca_clk cell_2907 ( .C (clk), .D (signal_3029), .Q (signal_12797) ) ;
    buf_sca_clk cell_2908 ( .C (clk), .D (signal_658), .Q (signal_12798) ) ;
    buf_sca_clk cell_2909 ( .C (clk), .D (signal_3031), .Q (signal_12799) ) ;
    buf_sca_clk cell_2910 ( .C (clk), .D (signal_660), .Q (signal_12800) ) ;
    buf_sca_clk cell_2911 ( .C (clk), .D (signal_3033), .Q (signal_12801) ) ;
    buf_sca_clk cell_2912 ( .C (clk), .D (signal_662), .Q (signal_12802) ) ;
    buf_sca_clk cell_2913 ( .C (clk), .D (signal_3035), .Q (signal_12803) ) ;
    buf_sca_clk cell_2914 ( .C (clk), .D (signal_664), .Q (signal_12804) ) ;
    buf_sca_clk cell_2915 ( .C (clk), .D (signal_3037), .Q (signal_12805) ) ;
    buf_sca_clk cell_2916 ( .C (clk), .D (signal_666), .Q (signal_12806) ) ;
    buf_sca_clk cell_2917 ( .C (clk), .D (signal_3039), .Q (signal_12807) ) ;
    buf_sca_clk cell_2918 ( .C (clk), .D (signal_668), .Q (signal_12808) ) ;
    buf_sca_clk cell_2919 ( .C (clk), .D (signal_3041), .Q (signal_12809) ) ;
    buf_clk cell_2920 ( .C (clk), .D (signal_1502), .Q (signal_12810) ) ;
    buf_clk cell_2921 ( .C (clk), .D (signal_1501), .Q (signal_12811) ) ;
    buf_clk cell_2922 ( .C (clk), .D (signal_1499), .Q (signal_12812) ) ;
    buf_clk cell_2923 ( .C (clk), .D (signal_1498), .Q (signal_12813) ) ;
    buf_clk cell_2924 ( .C (clk), .D (signal_1520), .Q (signal_12814) ) ;
    buf_clk cell_2925 ( .C (clk), .D (signal_1519), .Q (signal_12815) ) ;
    buf_clk cell_2926 ( .C (clk), .D (signal_1518), .Q (signal_12816) ) ;

    /* register cells */
    reg_masked #(.low_latency(1), .pipeline(1)) cell_159 ( .D ({signal_3437, signal_414}), .clk (clk), .Q ({ciphertext_s1[32], ciphertext_s0[32]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_162 ( .D ({signal_3263, signal_416}), .clk (clk), .Q ({ciphertext_s1[33], ciphertext_s0[33]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_165 ( .D ({signal_3265, signal_418}), .clk (clk), .Q ({ciphertext_s1[34], ciphertext_s0[34]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_168 ( .D ({signal_3267, signal_420}), .clk (clk), .Q ({ciphertext_s1[35], ciphertext_s0[35]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_171 ( .D ({signal_3269, signal_422}), .clk (clk), .Q ({ciphertext_s1[36], ciphertext_s0[36]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_174 ( .D ({signal_3271, signal_424}), .clk (clk), .Q ({ciphertext_s1[37], ciphertext_s0[37]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_177 ( .D ({signal_3273, signal_426}), .clk (clk), .Q ({ciphertext_s1[38], ciphertext_s0[38]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_180 ( .D ({signal_3275, signal_428}), .clk (clk), .Q ({ciphertext_s1[39], ciphertext_s0[39]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_183 ( .D ({signal_3277, signal_430}), .clk (clk), .Q ({ciphertext_s1[72], ciphertext_s0[72]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_186 ( .D ({signal_3439, signal_432}), .clk (clk), .Q ({ciphertext_s1[73], ciphertext_s0[73]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_189 ( .D ({signal_3279, signal_434}), .clk (clk), .Q ({ciphertext_s1[74], ciphertext_s0[74]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_192 ( .D ({signal_3281, signal_436}), .clk (clk), .Q ({ciphertext_s1[75], ciphertext_s0[75]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_195 ( .D ({signal_3283, signal_438}), .clk (clk), .Q ({ciphertext_s1[76], ciphertext_s0[76]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_198 ( .D ({signal_3285, signal_440}), .clk (clk), .Q ({ciphertext_s1[77], ciphertext_s0[77]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_201 ( .D ({signal_3287, signal_442}), .clk (clk), .Q ({ciphertext_s1[78], ciphertext_s0[78]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_204 ( .D ({signal_3289, signal_444}), .clk (clk), .Q ({ciphertext_s1[79], ciphertext_s0[79]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_207 ( .D ({signal_3291, signal_446}), .clk (clk), .Q ({ciphertext_s1[112], ciphertext_s0[112]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_210 ( .D ({signal_3293, signal_448}), .clk (clk), .Q ({ciphertext_s1[113], ciphertext_s0[113]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_213 ( .D ({signal_3295, signal_450}), .clk (clk), .Q ({ciphertext_s1[114], ciphertext_s0[114]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_216 ( .D ({signal_3297, signal_452}), .clk (clk), .Q ({ciphertext_s1[115], ciphertext_s0[115]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_219 ( .D ({signal_3299, signal_454}), .clk (clk), .Q ({ciphertext_s1[116], ciphertext_s0[116]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_222 ( .D ({signal_3301, signal_456}), .clk (clk), .Q ({ciphertext_s1[117], ciphertext_s0[117]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_225 ( .D ({signal_3303, signal_458}), .clk (clk), .Q ({ciphertext_s1[118], ciphertext_s0[118]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_228 ( .D ({signal_3305, signal_460}), .clk (clk), .Q ({ciphertext_s1[119], ciphertext_s0[119]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_231 ( .D ({signal_3307, signal_462}), .clk (clk), .Q ({ciphertext_s1[24], ciphertext_s0[24]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_234 ( .D ({signal_3309, signal_464}), .clk (clk), .Q ({ciphertext_s1[25], ciphertext_s0[25]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_237 ( .D ({signal_3311, signal_466}), .clk (clk), .Q ({ciphertext_s1[26], ciphertext_s0[26]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_240 ( .D ({signal_3313, signal_468}), .clk (clk), .Q ({ciphertext_s1[27], ciphertext_s0[27]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_243 ( .D ({signal_3315, signal_470}), .clk (clk), .Q ({ciphertext_s1[28], ciphertext_s0[28]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_246 ( .D ({signal_3317, signal_472}), .clk (clk), .Q ({ciphertext_s1[29], ciphertext_s0[29]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_249 ( .D ({signal_3319, signal_474}), .clk (clk), .Q ({ciphertext_s1[30], ciphertext_s0[30]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_252 ( .D ({signal_3321, signal_476}), .clk (clk), .Q ({ciphertext_s1[31], ciphertext_s0[31]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_255 ( .D ({signal_12619, signal_12618}), .clk (clk), .Q ({ciphertext_s1[64], ciphertext_s0[64]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_258 ( .D ({signal_12621, signal_12620}), .clk (clk), .Q ({ciphertext_s1[65], ciphertext_s0[65]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_261 ( .D ({signal_12623, signal_12622}), .clk (clk), .Q ({ciphertext_s1[66], ciphertext_s0[66]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_264 ( .D ({signal_12625, signal_12624}), .clk (clk), .Q ({ciphertext_s1[67], ciphertext_s0[67]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_267 ( .D ({signal_12627, signal_12626}), .clk (clk), .Q ({ciphertext_s1[68], ciphertext_s0[68]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_270 ( .D ({signal_12629, signal_12628}), .clk (clk), .Q ({ciphertext_s1[69], ciphertext_s0[69]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_273 ( .D ({signal_12631, signal_12630}), .clk (clk), .Q ({ciphertext_s1[70], ciphertext_s0[70]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_276 ( .D ({signal_12633, signal_12632}), .clk (clk), .Q ({ciphertext_s1[71], ciphertext_s0[71]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_279 ( .D ({signal_12635, signal_12634}), .clk (clk), .Q ({ciphertext_s1[104], ciphertext_s0[104]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_282 ( .D ({signal_12637, signal_12636}), .clk (clk), .Q ({ciphertext_s1[105], ciphertext_s0[105]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_285 ( .D ({signal_12639, signal_12638}), .clk (clk), .Q ({ciphertext_s1[106], ciphertext_s0[106]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_288 ( .D ({signal_12641, signal_12640}), .clk (clk), .Q ({ciphertext_s1[107], ciphertext_s0[107]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_291 ( .D ({signal_12643, signal_12642}), .clk (clk), .Q ({ciphertext_s1[108], ciphertext_s0[108]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_294 ( .D ({signal_12645, signal_12644}), .clk (clk), .Q ({ciphertext_s1[109], ciphertext_s0[109]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_297 ( .D ({signal_12647, signal_12646}), .clk (clk), .Q ({ciphertext_s1[110], ciphertext_s0[110]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_300 ( .D ({signal_12649, signal_12648}), .clk (clk), .Q ({ciphertext_s1[111], ciphertext_s0[111]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_303 ( .D ({signal_12651, signal_12650}), .clk (clk), .Q ({ciphertext_s1[16], ciphertext_s0[16]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_306 ( .D ({signal_12653, signal_12652}), .clk (clk), .Q ({ciphertext_s1[17], ciphertext_s0[17]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_309 ( .D ({signal_12655, signal_12654}), .clk (clk), .Q ({ciphertext_s1[18], ciphertext_s0[18]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_312 ( .D ({signal_12657, signal_12656}), .clk (clk), .Q ({ciphertext_s1[19], ciphertext_s0[19]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_315 ( .D ({signal_12659, signal_12658}), .clk (clk), .Q ({ciphertext_s1[20], ciphertext_s0[20]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_318 ( .D ({signal_12661, signal_12660}), .clk (clk), .Q ({ciphertext_s1[21], ciphertext_s0[21]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_321 ( .D ({signal_12663, signal_12662}), .clk (clk), .Q ({ciphertext_s1[22], ciphertext_s0[22]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_324 ( .D ({signal_12665, signal_12664}), .clk (clk), .Q ({ciphertext_s1[23], ciphertext_s0[23]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_327 ( .D ({signal_12667, signal_12666}), .clk (clk), .Q ({ciphertext_s1[56], ciphertext_s0[56]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_330 ( .D ({signal_12669, signal_12668}), .clk (clk), .Q ({ciphertext_s1[57], ciphertext_s0[57]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_333 ( .D ({signal_12671, signal_12670}), .clk (clk), .Q ({ciphertext_s1[58], ciphertext_s0[58]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_336 ( .D ({signal_12673, signal_12672}), .clk (clk), .Q ({ciphertext_s1[59], ciphertext_s0[59]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_339 ( .D ({signal_12675, signal_12674}), .clk (clk), .Q ({ciphertext_s1[60], ciphertext_s0[60]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_342 ( .D ({signal_12677, signal_12676}), .clk (clk), .Q ({ciphertext_s1[61], ciphertext_s0[61]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_345 ( .D ({signal_12679, signal_12678}), .clk (clk), .Q ({ciphertext_s1[62], ciphertext_s0[62]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_348 ( .D ({signal_12681, signal_12680}), .clk (clk), .Q ({ciphertext_s1[63], ciphertext_s0[63]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_351 ( .D ({signal_12683, signal_12682}), .clk (clk), .Q ({ciphertext_s1[96], ciphertext_s0[96]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_354 ( .D ({signal_12685, signal_12684}), .clk (clk), .Q ({ciphertext_s1[97], ciphertext_s0[97]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_357 ( .D ({signal_12687, signal_12686}), .clk (clk), .Q ({ciphertext_s1[98], ciphertext_s0[98]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_360 ( .D ({signal_12689, signal_12688}), .clk (clk), .Q ({ciphertext_s1[99], ciphertext_s0[99]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_363 ( .D ({signal_12691, signal_12690}), .clk (clk), .Q ({ciphertext_s1[100], ciphertext_s0[100]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_366 ( .D ({signal_12693, signal_12692}), .clk (clk), .Q ({ciphertext_s1[101], ciphertext_s0[101]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_369 ( .D ({signal_12695, signal_12694}), .clk (clk), .Q ({ciphertext_s1[102], ciphertext_s0[102]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_372 ( .D ({signal_12697, signal_12696}), .clk (clk), .Q ({ciphertext_s1[103], ciphertext_s0[103]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_375 ( .D ({signal_12699, signal_12698}), .clk (clk), .Q ({ciphertext_s1[8], ciphertext_s0[8]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_378 ( .D ({signal_12701, signal_12700}), .clk (clk), .Q ({ciphertext_s1[9], ciphertext_s0[9]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_381 ( .D ({signal_12703, signal_12702}), .clk (clk), .Q ({ciphertext_s1[10], ciphertext_s0[10]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_384 ( .D ({signal_12705, signal_12704}), .clk (clk), .Q ({ciphertext_s1[11], ciphertext_s0[11]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_387 ( .D ({signal_12707, signal_12706}), .clk (clk), .Q ({ciphertext_s1[12], ciphertext_s0[12]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_390 ( .D ({signal_12709, signal_12708}), .clk (clk), .Q ({ciphertext_s1[13], ciphertext_s0[13]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_393 ( .D ({signal_12711, signal_12710}), .clk (clk), .Q ({ciphertext_s1[14], ciphertext_s0[14]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_396 ( .D ({signal_12713, signal_12712}), .clk (clk), .Q ({ciphertext_s1[15], ciphertext_s0[15]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_399 ( .D ({signal_12715, signal_12714}), .clk (clk), .Q ({ciphertext_s1[48], ciphertext_s0[48]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_402 ( .D ({signal_12717, signal_12716}), .clk (clk), .Q ({ciphertext_s1[49], ciphertext_s0[49]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_405 ( .D ({signal_12719, signal_12718}), .clk (clk), .Q ({ciphertext_s1[50], ciphertext_s0[50]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_408 ( .D ({signal_12721, signal_12720}), .clk (clk), .Q ({ciphertext_s1[51], ciphertext_s0[51]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_411 ( .D ({signal_12723, signal_12722}), .clk (clk), .Q ({ciphertext_s1[52], ciphertext_s0[52]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_414 ( .D ({signal_12725, signal_12724}), .clk (clk), .Q ({ciphertext_s1[53], ciphertext_s0[53]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_417 ( .D ({signal_12727, signal_12726}), .clk (clk), .Q ({ciphertext_s1[54], ciphertext_s0[54]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_420 ( .D ({signal_12729, signal_12728}), .clk (clk), .Q ({ciphertext_s1[55], ciphertext_s0[55]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_423 ( .D ({signal_12731, signal_12730}), .clk (clk), .Q ({ciphertext_s1[88], ciphertext_s0[88]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_426 ( .D ({signal_12733, signal_12732}), .clk (clk), .Q ({ciphertext_s1[89], ciphertext_s0[89]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_429 ( .D ({signal_12735, signal_12734}), .clk (clk), .Q ({ciphertext_s1[90], ciphertext_s0[90]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_432 ( .D ({signal_12737, signal_12736}), .clk (clk), .Q ({ciphertext_s1[91], ciphertext_s0[91]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_435 ( .D ({signal_12739, signal_12738}), .clk (clk), .Q ({ciphertext_s1[92], ciphertext_s0[92]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_438 ( .D ({signal_12741, signal_12740}), .clk (clk), .Q ({ciphertext_s1[93], ciphertext_s0[93]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_441 ( .D ({signal_12743, signal_12742}), .clk (clk), .Q ({ciphertext_s1[94], ciphertext_s0[94]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_444 ( .D ({signal_12745, signal_12744}), .clk (clk), .Q ({ciphertext_s1[95], ciphertext_s0[95]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_447 ( .D ({signal_12747, signal_12746}), .clk (clk), .Q ({ciphertext_s1[0], ciphertext_s0[0]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_450 ( .D ({signal_12749, signal_12748}), .clk (clk), .Q ({ciphertext_s1[1], ciphertext_s0[1]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_453 ( .D ({signal_12751, signal_12750}), .clk (clk), .Q ({ciphertext_s1[2], ciphertext_s0[2]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_456 ( .D ({signal_12753, signal_12752}), .clk (clk), .Q ({ciphertext_s1[3], ciphertext_s0[3]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_459 ( .D ({signal_12755, signal_12754}), .clk (clk), .Q ({ciphertext_s1[4], ciphertext_s0[4]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_462 ( .D ({signal_12757, signal_12756}), .clk (clk), .Q ({ciphertext_s1[5], ciphertext_s0[5]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_465 ( .D ({signal_12759, signal_12758}), .clk (clk), .Q ({ciphertext_s1[6], ciphertext_s0[6]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_468 ( .D ({signal_12761, signal_12760}), .clk (clk), .Q ({ciphertext_s1[7], ciphertext_s0[7]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_471 ( .D ({signal_12763, signal_12762}), .clk (clk), .Q ({ciphertext_s1[40], ciphertext_s0[40]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_474 ( .D ({signal_12765, signal_12764}), .clk (clk), .Q ({ciphertext_s1[41], ciphertext_s0[41]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_477 ( .D ({signal_12767, signal_12766}), .clk (clk), .Q ({ciphertext_s1[42], ciphertext_s0[42]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_480 ( .D ({signal_12769, signal_12768}), .clk (clk), .Q ({ciphertext_s1[43], ciphertext_s0[43]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_483 ( .D ({signal_12771, signal_12770}), .clk (clk), .Q ({ciphertext_s1[44], ciphertext_s0[44]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_486 ( .D ({signal_12773, signal_12772}), .clk (clk), .Q ({ciphertext_s1[45], ciphertext_s0[45]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_489 ( .D ({signal_12775, signal_12774}), .clk (clk), .Q ({ciphertext_s1[46], ciphertext_s0[46]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_492 ( .D ({signal_12777, signal_12776}), .clk (clk), .Q ({ciphertext_s1[47], ciphertext_s0[47]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_495 ( .D ({signal_12779, signal_12778}), .clk (clk), .Q ({ciphertext_s1[80], ciphertext_s0[80]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_498 ( .D ({signal_12781, signal_12780}), .clk (clk), .Q ({ciphertext_s1[81], ciphertext_s0[81]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_501 ( .D ({signal_12783, signal_12782}), .clk (clk), .Q ({ciphertext_s1[82], ciphertext_s0[82]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_504 ( .D ({signal_12785, signal_12784}), .clk (clk), .Q ({ciphertext_s1[83], ciphertext_s0[83]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_507 ( .D ({signal_12787, signal_12786}), .clk (clk), .Q ({ciphertext_s1[84], ciphertext_s0[84]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_510 ( .D ({signal_12789, signal_12788}), .clk (clk), .Q ({ciphertext_s1[85], ciphertext_s0[85]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_513 ( .D ({signal_12791, signal_12790}), .clk (clk), .Q ({ciphertext_s1[86], ciphertext_s0[86]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_516 ( .D ({signal_12793, signal_12792}), .clk (clk), .Q ({ciphertext_s1[87], ciphertext_s0[87]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_519 ( .D ({signal_12795, signal_12794}), .clk (clk), .Q ({ciphertext_s1[120], ciphertext_s0[120]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_522 ( .D ({signal_12797, signal_12796}), .clk (clk), .Q ({ciphertext_s1[121], ciphertext_s0[121]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_525 ( .D ({signal_12799, signal_12798}), .clk (clk), .Q ({ciphertext_s1[122], ciphertext_s0[122]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_528 ( .D ({signal_12801, signal_12800}), .clk (clk), .Q ({ciphertext_s1[123], ciphertext_s0[123]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_531 ( .D ({signal_12803, signal_12802}), .clk (clk), .Q ({ciphertext_s1[124], ciphertext_s0[124]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_534 ( .D ({signal_12805, signal_12804}), .clk (clk), .Q ({ciphertext_s1[125], ciphertext_s0[125]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_537 ( .D ({signal_12807, signal_12806}), .clk (clk), .Q ({ciphertext_s1[126], ciphertext_s0[126]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_540 ( .D ({signal_12809, signal_12808}), .clk (clk), .Q ({ciphertext_s1[127], ciphertext_s0[127]}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1368 ( .D ({signal_3673, signal_1227}), .clk (clk), .Q ({signal_2339, signal_1793}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1371 ( .D ({signal_3675, signal_1229}), .clk (clk), .Q ({signal_2456, signal_1792}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1374 ( .D ({signal_3677, signal_1231}), .clk (clk), .Q ({signal_2489, signal_1791}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1377 ( .D ({signal_3679, signal_1233}), .clk (clk), .Q ({signal_2522, signal_1790}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1380 ( .D ({signal_3681, signal_1235}), .clk (clk), .Q ({signal_2555, signal_1789}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1383 ( .D ({signal_3683, signal_1237}), .clk (clk), .Q ({signal_2588, signal_1788}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1386 ( .D ({signal_3685, signal_1239}), .clk (clk), .Q ({signal_2621, signal_1787}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1389 ( .D ({signal_3687, signal_1241}), .clk (clk), .Q ({signal_2654, signal_1786}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1392 ( .D ({signal_3689, signal_1243}), .clk (clk), .Q ({signal_2687, signal_1801}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1395 ( .D ({signal_3691, signal_1245}), .clk (clk), .Q ({signal_2720, signal_1800}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1398 ( .D ({signal_3693, signal_1247}), .clk (clk), .Q ({signal_2372, signal_1799}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1401 ( .D ({signal_3695, signal_1249}), .clk (clk), .Q ({signal_2405, signal_1798}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1404 ( .D ({signal_3697, signal_1251}), .clk (clk), .Q ({signal_2432, signal_1797}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1407 ( .D ({signal_3699, signal_1253}), .clk (clk), .Q ({signal_2435, signal_1796}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1410 ( .D ({signal_3701, signal_1255}), .clk (clk), .Q ({signal_2438, signal_1795}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1413 ( .D ({signal_3703, signal_1257}), .clk (clk), .Q ({signal_2441, signal_1794}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1416 ( .D ({signal_3705, signal_1259}), .clk (clk), .Q ({signal_2444, signal_1809}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1419 ( .D ({signal_3707, signal_1261}), .clk (clk), .Q ({signal_2447, signal_1808}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1422 ( .D ({signal_3709, signal_1263}), .clk (clk), .Q ({signal_2450, signal_1807}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1425 ( .D ({signal_3711, signal_1265}), .clk (clk), .Q ({signal_2453, signal_1806}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1428 ( .D ({signal_3713, signal_1267}), .clk (clk), .Q ({signal_2459, signal_1805}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1431 ( .D ({signal_3715, signal_1269}), .clk (clk), .Q ({signal_2462, signal_1804}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1434 ( .D ({signal_3717, signal_1271}), .clk (clk), .Q ({signal_2465, signal_1803}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1437 ( .D ({signal_3719, signal_1273}), .clk (clk), .Q ({signal_2468, signal_1802}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1440 ( .D ({signal_3745, signal_1275}), .clk (clk), .Q ({signal_2471, signal_1785}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1443 ( .D ({signal_3747, signal_1277}), .clk (clk), .Q ({signal_2474, signal_1784}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1446 ( .D ({signal_3749, signal_1279}), .clk (clk), .Q ({signal_2477, signal_1783}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1449 ( .D ({signal_3751, signal_1281}), .clk (clk), .Q ({signal_2480, signal_1782}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1452 ( .D ({signal_3753, signal_1283}), .clk (clk), .Q ({signal_2483, signal_1781}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1455 ( .D ({signal_3755, signal_1285}), .clk (clk), .Q ({signal_2486, signal_1780}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1458 ( .D ({signal_3757, signal_1287}), .clk (clk), .Q ({signal_2492, signal_1779}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1461 ( .D ({signal_3759, signal_1289}), .clk (clk), .Q ({signal_2495, signal_1778}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1464 ( .D ({signal_3569, signal_1291}), .clk (clk), .Q ({signal_2498, signal_2133}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1467 ( .D ({signal_3571, signal_1293}), .clk (clk), .Q ({signal_2501, signal_2132}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1470 ( .D ({signal_3573, signal_1295}), .clk (clk), .Q ({signal_2504, signal_2131}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1473 ( .D ({signal_3575, signal_1297}), .clk (clk), .Q ({signal_2507, signal_2130}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1476 ( .D ({signal_3577, signal_1299}), .clk (clk), .Q ({signal_2510, signal_2129}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1479 ( .D ({signal_3579, signal_1301}), .clk (clk), .Q ({signal_2513, signal_2128}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1482 ( .D ({signal_3581, signal_1303}), .clk (clk), .Q ({signal_2516, signal_2127}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1485 ( .D ({signal_3583, signal_1305}), .clk (clk), .Q ({signal_2519, signal_2126}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1488 ( .D ({signal_3585, signal_1307}), .clk (clk), .Q ({signal_2525, signal_2125}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1491 ( .D ({signal_3587, signal_1309}), .clk (clk), .Q ({signal_2528, signal_2124}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1494 ( .D ({signal_3589, signal_1311}), .clk (clk), .Q ({signal_2531, signal_2123}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1497 ( .D ({signal_3591, signal_1313}), .clk (clk), .Q ({signal_2534, signal_2122}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1500 ( .D ({signal_3593, signal_1315}), .clk (clk), .Q ({signal_2537, signal_2121}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1503 ( .D ({signal_3595, signal_1317}), .clk (clk), .Q ({signal_2540, signal_2120}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1506 ( .D ({signal_3597, signal_1319}), .clk (clk), .Q ({signal_2543, signal_2119}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1509 ( .D ({signal_3599, signal_1321}), .clk (clk), .Q ({signal_2546, signal_2118}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1512 ( .D ({signal_3601, signal_1323}), .clk (clk), .Q ({signal_2549, signal_2117}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1515 ( .D ({signal_3603, signal_1325}), .clk (clk), .Q ({signal_2552, signal_2116}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1518 ( .D ({signal_3605, signal_1327}), .clk (clk), .Q ({signal_2558, signal_2115}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1521 ( .D ({signal_3607, signal_1329}), .clk (clk), .Q ({signal_2561, signal_2114}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1524 ( .D ({signal_3609, signal_1331}), .clk (clk), .Q ({signal_2564, signal_2113}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1527 ( .D ({signal_3611, signal_1333}), .clk (clk), .Q ({signal_2567, signal_2112}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1530 ( .D ({signal_3613, signal_1335}), .clk (clk), .Q ({signal_2570, signal_2111}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1533 ( .D ({signal_3615, signal_1337}), .clk (clk), .Q ({signal_2573, signal_2110}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1536 ( .D ({signal_3721, signal_1339}), .clk (clk), .Q ({signal_2576, signal_2109}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1539 ( .D ({signal_3723, signal_1341}), .clk (clk), .Q ({signal_2579, signal_2108}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1542 ( .D ({signal_3725, signal_1343}), .clk (clk), .Q ({signal_2582, signal_2107}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1545 ( .D ({signal_3727, signal_1345}), .clk (clk), .Q ({signal_2585, signal_2106}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1548 ( .D ({signal_3729, signal_1347}), .clk (clk), .Q ({signal_2591, signal_2105}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1551 ( .D ({signal_3731, signal_1349}), .clk (clk), .Q ({signal_2594, signal_2104}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1554 ( .D ({signal_3733, signal_1351}), .clk (clk), .Q ({signal_2597, signal_2103}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1557 ( .D ({signal_3735, signal_1353}), .clk (clk), .Q ({signal_2600, signal_2102}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1560 ( .D ({signal_3441, signal_1355}), .clk (clk), .Q ({signal_2603, signal_2101}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1563 ( .D ({signal_3443, signal_1357}), .clk (clk), .Q ({signal_2606, signal_2100}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1566 ( .D ({signal_3445, signal_1359}), .clk (clk), .Q ({signal_2609, signal_2099}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1569 ( .D ({signal_3447, signal_1361}), .clk (clk), .Q ({signal_2612, signal_2098}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1572 ( .D ({signal_3449, signal_1363}), .clk (clk), .Q ({signal_2615, signal_2097}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1575 ( .D ({signal_3451, signal_1365}), .clk (clk), .Q ({signal_2618, signal_2096}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1578 ( .D ({signal_3453, signal_1367}), .clk (clk), .Q ({signal_2624, signal_2095}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1581 ( .D ({signal_3455, signal_1369}), .clk (clk), .Q ({signal_2627, signal_2094}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1584 ( .D ({signal_3457, signal_1371}), .clk (clk), .Q ({signal_2630, signal_2093}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1587 ( .D ({signal_3459, signal_1373}), .clk (clk), .Q ({signal_2633, signal_2092}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1590 ( .D ({signal_3461, signal_1375}), .clk (clk), .Q ({signal_2636, signal_2091}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1593 ( .D ({signal_3463, signal_1377}), .clk (clk), .Q ({signal_2639, signal_2090}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1596 ( .D ({signal_3465, signal_1379}), .clk (clk), .Q ({signal_2642, signal_2089}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1599 ( .D ({signal_3467, signal_1381}), .clk (clk), .Q ({signal_2645, signal_2088}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1602 ( .D ({signal_3469, signal_1383}), .clk (clk), .Q ({signal_2648, signal_2087}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1605 ( .D ({signal_3471, signal_1385}), .clk (clk), .Q ({signal_2651, signal_2086}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1608 ( .D ({signal_3473, signal_1387}), .clk (clk), .Q ({signal_2657, signal_2085}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1611 ( .D ({signal_3475, signal_1389}), .clk (clk), .Q ({signal_2660, signal_2084}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1614 ( .D ({signal_3477, signal_1391}), .clk (clk), .Q ({signal_2663, signal_2083}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1617 ( .D ({signal_3479, signal_1393}), .clk (clk), .Q ({signal_2666, signal_2082}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1620 ( .D ({signal_3481, signal_1395}), .clk (clk), .Q ({signal_2669, signal_2081}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1623 ( .D ({signal_3483, signal_1397}), .clk (clk), .Q ({signal_2672, signal_2080}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1626 ( .D ({signal_3485, signal_1399}), .clk (clk), .Q ({signal_2675, signal_2079}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1629 ( .D ({signal_3487, signal_1401}), .clk (clk), .Q ({signal_2678, signal_2078}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1632 ( .D ({signal_3617, signal_1403}), .clk (clk), .Q ({signal_2681, signal_2077}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1635 ( .D ({signal_3619, signal_1405}), .clk (clk), .Q ({signal_2684, signal_2076}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1638 ( .D ({signal_3621, signal_1407}), .clk (clk), .Q ({signal_2690, signal_2075}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1641 ( .D ({signal_3623, signal_1409}), .clk (clk), .Q ({signal_2693, signal_2074}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1644 ( .D ({signal_3625, signal_1411}), .clk (clk), .Q ({signal_2696, signal_2073}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1647 ( .D ({signal_3627, signal_1413}), .clk (clk), .Q ({signal_2699, signal_2072}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1650 ( .D ({signal_3629, signal_1415}), .clk (clk), .Q ({signal_2702, signal_2071}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1653 ( .D ({signal_3631, signal_1417}), .clk (clk), .Q ({signal_2705, signal_2070}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1656 ( .D ({signal_3325, signal_1419}), .clk (clk), .Q ({signal_2708, signal_2069}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1659 ( .D ({signal_3327, signal_1421}), .clk (clk), .Q ({signal_2711, signal_2068}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1662 ( .D ({signal_3329, signal_1423}), .clk (clk), .Q ({signal_2714, signal_2067}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1665 ( .D ({signal_3331, signal_1425}), .clk (clk), .Q ({signal_2717, signal_2066}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1668 ( .D ({signal_3333, signal_1427}), .clk (clk), .Q ({signal_2342, signal_2065}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1671 ( .D ({signal_3335, signal_1429}), .clk (clk), .Q ({signal_2345, signal_2064}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1674 ( .D ({signal_3337, signal_1431}), .clk (clk), .Q ({signal_2348, signal_2063}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1677 ( .D ({signal_3339, signal_1433}), .clk (clk), .Q ({signal_2351, signal_2062}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1680 ( .D ({signal_3341, signal_1435}), .clk (clk), .Q ({signal_2354, signal_2061}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1683 ( .D ({signal_3343, signal_1437}), .clk (clk), .Q ({signal_2357, signal_2060}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1686 ( .D ({signal_3345, signal_1439}), .clk (clk), .Q ({signal_2360, signal_2059}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1689 ( .D ({signal_3347, signal_1441}), .clk (clk), .Q ({signal_2363, signal_2058}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1692 ( .D ({signal_3349, signal_1443}), .clk (clk), .Q ({signal_2366, signal_2057}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1695 ( .D ({signal_3351, signal_1445}), .clk (clk), .Q ({signal_2369, signal_2056}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1698 ( .D ({signal_3353, signal_1447}), .clk (clk), .Q ({signal_2375, signal_2055}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1701 ( .D ({signal_3355, signal_1449}), .clk (clk), .Q ({signal_2378, signal_2054}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1704 ( .D ({signal_3357, signal_1451}), .clk (clk), .Q ({signal_2381, signal_2053}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1707 ( .D ({signal_3359, signal_1453}), .clk (clk), .Q ({signal_2384, signal_2052}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1710 ( .D ({signal_3361, signal_1455}), .clk (clk), .Q ({signal_2387, signal_2051}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1713 ( .D ({signal_3363, signal_1457}), .clk (clk), .Q ({signal_2390, signal_2050}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1716 ( .D ({signal_3365, signal_1459}), .clk (clk), .Q ({signal_2393, signal_2049}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1719 ( .D ({signal_3367, signal_1461}), .clk (clk), .Q ({signal_2396, signal_2048}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1722 ( .D ({signal_3369, signal_1463}), .clk (clk), .Q ({signal_2399, signal_2047}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1725 ( .D ({signal_3371, signal_1465}), .clk (clk), .Q ({signal_2402, signal_2046}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1728 ( .D ({signal_3489, signal_1467}), .clk (clk), .Q ({signal_2408, signal_2045}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1731 ( .D ({signal_3491, signal_1469}), .clk (clk), .Q ({signal_2411, signal_2044}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1734 ( .D ({signal_3493, signal_1471}), .clk (clk), .Q ({signal_2414, signal_2043}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1737 ( .D ({signal_3495, signal_1473}), .clk (clk), .Q ({signal_2417, signal_2042}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1740 ( .D ({signal_3497, signal_1475}), .clk (clk), .Q ({signal_2420, signal_2041}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1743 ( .D ({signal_3499, signal_1477}), .clk (clk), .Q ({signal_2423, signal_2040}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1746 ( .D ({signal_3501, signal_1479}), .clk (clk), .Q ({signal_2426, signal_2039}) ) ;
    reg_masked #(.low_latency(1), .pipeline(1)) cell_1749 ( .D ({signal_3503, signal_1481}), .clk (clk), .Q ({signal_2429, signal_2038}) ) ;
    DFF_X1 cell_2035 ( .D (signal_12810), .CK (clk), .Q (signal_2273), .QN () ) ;
    DFF_X1 cell_2037 ( .D (signal_12811), .CK (clk), .Q (signal_2272), .QN () ) ;
    DFF_X1 cell_2039 ( .D (signal_12812), .CK (clk), .Q (signal_2271), .QN () ) ;
    DFF_X1 cell_2041 ( .D (signal_12813), .CK (clk), .Q (signal_2270), .QN () ) ;
    DFF_X1 cell_2056 ( .D (signal_12814), .CK (clk), .Q (signal_2276), .QN () ) ;
    DFF_X1 cell_2058 ( .D (signal_12815), .CK (clk), .Q (signal_2275), .QN () ) ;
    DFF_X1 cell_2060 ( .D (signal_12816), .CK (clk), .Q (signal_2274), .QN () ) ;
endmodule
