/* modified netlist. Source: module LED in file ../CaseStudies/11_LED_round_based_encryption/FPGA_based/LED_synthesis.v */
/* clock gating is added to the circuit, the latency increased 1 time(s)  */

module LED_GHPCLL_ClockGating_d1 (CLK, IN_reset, IN_plaintext_s0, IN_key_s0, IN_key_s1, IN_plaintext_s1, Fresh, OUT_done, OUT_ciphertext_s0, OUT_ciphertext_s1, Synch);
    input CLK ;
    input IN_reset ;
    input [63:0] IN_plaintext_s0 ;
    input [127:0] IN_key_s0 ;
    input [127:0] IN_key_s1 ;
    input [63:0] IN_plaintext_s1 ;
    input [1023:0] Fresh ;
    output OUT_done ;
    output [63:0] OUT_ciphertext_s0 ;
    output [63:0] OUT_ciphertext_s1 ;
    output Synch ;
    wire \LED_128_Instance/addkey1_265 ;
    wire \LED_128_Instance/roundconstant[5]_roundconstant[4]_XOR_7_o ;
    wire \LED_128_Instance/addkey ;
    wire \LED_128_Instance/roundconstant_001001 ;
    wire \LED_128_Instance/ks[3]_INV_6_o ;
    wire [54:3] \LED_128_Instance/addconst_out ;
    wire N2 ;
    wire N4 ;
    wire N6 ;
    wire N8 ;
    wire N12 ;
    wire N14 ;
    wire N16 ;
    wire N18 ;
    wire N20 ;
    wire N22 ;
    wire N24 ;
    wire N26 ;
    wire N28 ;
    wire N32 ;
    wire N34 ;
    wire N36 ;
    wire N38 ;
    wire N40 ;
    wire N42 ;
    wire N44 ;
    wire N46 ;
    wire N48 ;
    wire N52 ;
    wire N54 ;
    wire N56 ;
    wire N58 ;
    wire N60 ;
    wire N62 ;
    wire N64 ;
    wire N66 ;
    wire N68 ;
    wire N72 ;
    wire N74 ;
    wire N76 ;
    wire N78 ;
    wire N80 ;
    wire internal_done_glue_set_843 ;
    wire N82 ;
    wire N84 ;
    wire N86 ;
    wire N88 ;
    wire N90 ;
    wire N92 ;
    wire N94 ;
    wire N96 ;
    wire N98 ;
    wire N100 ;
    wire N102 ;
    wire N104 ;
    wire [5:0] \LED_128_Instance/roundconstant ;
    wire [63:0] \LED_128_Instance/mixcolumns_out ;
    wire [63:0] \LED_128_Instance/subcells_out ;
    wire [63:0] \LED_128_Instance/addroundkey_out ;
    wire [3:0] \LED_128_Instance/ks ;
    wire [63:0] \LED_128_Instance/state ;
    wire new_AGEMA_signal_865 ;
    wire new_AGEMA_signal_869 ;
    wire new_AGEMA_signal_873 ;
    wire new_AGEMA_signal_877 ;
    wire new_AGEMA_signal_881 ;
    wire new_AGEMA_signal_885 ;
    wire new_AGEMA_signal_889 ;
    wire new_AGEMA_signal_893 ;
    wire new_AGEMA_signal_897 ;
    wire new_AGEMA_signal_901 ;
    wire new_AGEMA_signal_905 ;
    wire new_AGEMA_signal_909 ;
    wire new_AGEMA_signal_913 ;
    wire new_AGEMA_signal_917 ;
    wire new_AGEMA_signal_921 ;
    wire new_AGEMA_signal_925 ;
    wire new_AGEMA_signal_929 ;
    wire new_AGEMA_signal_933 ;
    wire new_AGEMA_signal_937 ;
    wire new_AGEMA_signal_941 ;
    wire new_AGEMA_signal_945 ;
    wire new_AGEMA_signal_949 ;
    wire new_AGEMA_signal_953 ;
    wire new_AGEMA_signal_957 ;
    wire new_AGEMA_signal_961 ;
    wire new_AGEMA_signal_965 ;
    wire new_AGEMA_signal_969 ;
    wire new_AGEMA_signal_973 ;
    wire new_AGEMA_signal_977 ;
    wire new_AGEMA_signal_981 ;
    wire new_AGEMA_signal_985 ;
    wire new_AGEMA_signal_989 ;
    wire new_AGEMA_signal_993 ;
    wire new_AGEMA_signal_997 ;
    wire new_AGEMA_signal_1001 ;
    wire new_AGEMA_signal_1005 ;
    wire new_AGEMA_signal_1009 ;
    wire new_AGEMA_signal_1013 ;
    wire new_AGEMA_signal_1017 ;
    wire new_AGEMA_signal_1021 ;
    wire new_AGEMA_signal_1025 ;
    wire new_AGEMA_signal_1029 ;
    wire new_AGEMA_signal_1033 ;
    wire new_AGEMA_signal_1037 ;
    wire new_AGEMA_signal_1041 ;
    wire new_AGEMA_signal_1045 ;
    wire new_AGEMA_signal_1049 ;
    wire new_AGEMA_signal_1053 ;
    wire new_AGEMA_signal_1057 ;
    wire new_AGEMA_signal_1061 ;
    wire new_AGEMA_signal_1065 ;
    wire new_AGEMA_signal_1069 ;
    wire new_AGEMA_signal_1073 ;
    wire new_AGEMA_signal_1077 ;
    wire new_AGEMA_signal_1081 ;
    wire new_AGEMA_signal_1085 ;
    wire new_AGEMA_signal_1089 ;
    wire new_AGEMA_signal_1093 ;
    wire new_AGEMA_signal_1097 ;
    wire new_AGEMA_signal_1101 ;
    wire new_AGEMA_signal_1105 ;
    wire new_AGEMA_signal_1109 ;
    wire new_AGEMA_signal_1113 ;
    wire new_AGEMA_signal_1117 ;
    wire new_AGEMA_signal_1118 ;
    wire new_AGEMA_signal_1119 ;
    wire new_AGEMA_signal_1120 ;
    wire new_AGEMA_signal_1121 ;
    wire new_AGEMA_signal_1122 ;
    wire new_AGEMA_signal_1123 ;
    wire new_AGEMA_signal_1124 ;
    wire new_AGEMA_signal_1125 ;
    wire new_AGEMA_signal_1126 ;
    wire new_AGEMA_signal_1127 ;
    wire new_AGEMA_signal_1128 ;
    wire new_AGEMA_signal_1129 ;
    wire new_AGEMA_signal_1130 ;
    wire new_AGEMA_signal_1131 ;
    wire new_AGEMA_signal_1132 ;
    wire new_AGEMA_signal_1133 ;
    wire new_AGEMA_signal_1134 ;
    wire new_AGEMA_signal_1135 ;
    wire new_AGEMA_signal_1136 ;
    wire new_AGEMA_signal_1137 ;
    wire new_AGEMA_signal_1138 ;
    wire new_AGEMA_signal_1139 ;
    wire new_AGEMA_signal_1140 ;
    wire new_AGEMA_signal_1141 ;
    wire new_AGEMA_signal_1142 ;
    wire new_AGEMA_signal_1143 ;
    wire new_AGEMA_signal_1144 ;
    wire new_AGEMA_signal_1145 ;
    wire new_AGEMA_signal_1146 ;
    wire new_AGEMA_signal_1147 ;
    wire new_AGEMA_signal_1148 ;
    wire new_AGEMA_signal_1149 ;
    wire new_AGEMA_signal_1150 ;
    wire new_AGEMA_signal_1151 ;
    wire new_AGEMA_signal_1152 ;
    wire new_AGEMA_signal_1153 ;
    wire new_AGEMA_signal_1154 ;
    wire new_AGEMA_signal_1155 ;
    wire new_AGEMA_signal_1156 ;
    wire new_AGEMA_signal_1157 ;
    wire new_AGEMA_signal_1158 ;
    wire new_AGEMA_signal_1159 ;
    wire new_AGEMA_signal_1160 ;
    wire new_AGEMA_signal_1161 ;
    wire new_AGEMA_signal_1162 ;
    wire new_AGEMA_signal_1163 ;
    wire new_AGEMA_signal_1164 ;
    wire new_AGEMA_signal_1165 ;
    wire new_AGEMA_signal_1166 ;
    wire new_AGEMA_signal_1167 ;
    wire new_AGEMA_signal_1168 ;
    wire new_AGEMA_signal_1169 ;
    wire new_AGEMA_signal_1170 ;
    wire new_AGEMA_signal_1171 ;
    wire new_AGEMA_signal_1172 ;
    wire new_AGEMA_signal_1173 ;
    wire new_AGEMA_signal_1174 ;
    wire new_AGEMA_signal_1175 ;
    wire new_AGEMA_signal_1176 ;
    wire new_AGEMA_signal_1177 ;
    wire new_AGEMA_signal_1178 ;
    wire new_AGEMA_signal_1179 ;
    wire new_AGEMA_signal_1180 ;
    wire new_AGEMA_signal_1181 ;
    wire new_AGEMA_signal_1182 ;
    wire new_AGEMA_signal_1183 ;
    wire new_AGEMA_signal_1184 ;
    wire new_AGEMA_signal_1185 ;
    wire new_AGEMA_signal_1186 ;
    wire new_AGEMA_signal_1187 ;
    wire new_AGEMA_signal_1188 ;
    wire new_AGEMA_signal_1189 ;
    wire new_AGEMA_signal_1190 ;
    wire new_AGEMA_signal_1191 ;
    wire new_AGEMA_signal_1192 ;
    wire new_AGEMA_signal_1193 ;
    wire new_AGEMA_signal_1194 ;
    wire new_AGEMA_signal_1195 ;
    wire new_AGEMA_signal_1196 ;
    wire new_AGEMA_signal_1197 ;
    wire new_AGEMA_signal_1198 ;
    wire new_AGEMA_signal_1199 ;
    wire new_AGEMA_signal_1200 ;
    wire new_AGEMA_signal_1201 ;
    wire new_AGEMA_signal_1202 ;
    wire new_AGEMA_signal_1203 ;
    wire new_AGEMA_signal_1204 ;
    wire new_AGEMA_signal_1205 ;
    wire new_AGEMA_signal_1206 ;
    wire new_AGEMA_signal_1207 ;
    wire new_AGEMA_signal_1208 ;
    wire new_AGEMA_signal_1209 ;
    wire new_AGEMA_signal_1210 ;
    wire new_AGEMA_signal_1211 ;
    wire new_AGEMA_signal_1212 ;
    wire new_AGEMA_signal_1213 ;
    wire new_AGEMA_signal_1214 ;
    wire new_AGEMA_signal_1215 ;
    wire new_AGEMA_signal_1216 ;
    wire new_AGEMA_signal_1217 ;
    wire new_AGEMA_signal_1218 ;
    wire new_AGEMA_signal_1219 ;
    wire new_AGEMA_signal_1220 ;
    wire new_AGEMA_signal_1221 ;
    wire new_AGEMA_signal_1222 ;
    wire new_AGEMA_signal_1223 ;
    wire new_AGEMA_signal_1224 ;
    wire new_AGEMA_signal_1225 ;
    wire new_AGEMA_signal_1226 ;
    wire new_AGEMA_signal_1227 ;
    wire new_AGEMA_signal_1228 ;
    wire new_AGEMA_signal_1229 ;
    wire new_AGEMA_signal_1230 ;
    wire new_AGEMA_signal_1231 ;
    wire new_AGEMA_signal_1232 ;
    wire new_AGEMA_signal_1233 ;
    wire new_AGEMA_signal_1234 ;
    wire new_AGEMA_signal_1235 ;
    wire new_AGEMA_signal_1236 ;
    wire new_AGEMA_signal_1237 ;
    wire new_AGEMA_signal_1238 ;
    wire new_AGEMA_signal_1239 ;
    wire new_AGEMA_signal_1240 ;
    wire new_AGEMA_signal_1241 ;
    wire new_AGEMA_signal_1242 ;
    wire new_AGEMA_signal_1243 ;
    wire new_AGEMA_signal_1244 ;
    wire new_AGEMA_signal_1245 ;
    wire new_AGEMA_signal_1246 ;
    wire new_AGEMA_signal_1247 ;
    wire new_AGEMA_signal_1248 ;
    wire new_AGEMA_signal_1249 ;
    wire new_AGEMA_signal_1250 ;
    wire new_AGEMA_signal_1251 ;
    wire new_AGEMA_signal_1252 ;
    wire new_AGEMA_signal_1253 ;
    wire new_AGEMA_signal_1254 ;
    wire new_AGEMA_signal_1255 ;
    wire new_AGEMA_signal_1256 ;
    wire new_AGEMA_signal_1257 ;
    wire new_AGEMA_signal_1258 ;
    wire new_AGEMA_signal_1259 ;
    wire new_AGEMA_signal_1260 ;
    wire new_AGEMA_signal_1261 ;
    wire new_AGEMA_signal_1262 ;
    wire new_AGEMA_signal_1263 ;
    wire new_AGEMA_signal_1265 ;
    wire new_AGEMA_signal_1267 ;
    wire new_AGEMA_signal_1269 ;
    wire new_AGEMA_signal_1271 ;
    wire new_AGEMA_signal_1273 ;
    wire new_AGEMA_signal_1275 ;
    wire new_AGEMA_signal_1277 ;
    wire new_AGEMA_signal_1279 ;
    wire new_AGEMA_signal_1281 ;
    wire new_AGEMA_signal_1283 ;
    wire new_AGEMA_signal_1285 ;
    wire new_AGEMA_signal_1287 ;
    wire new_AGEMA_signal_1289 ;
    wire new_AGEMA_signal_1291 ;
    wire new_AGEMA_signal_1293 ;
    wire new_AGEMA_signal_1295 ;
    wire new_AGEMA_signal_1296 ;
    wire new_AGEMA_signal_1297 ;
    wire new_AGEMA_signal_1298 ;
    wire new_AGEMA_signal_1299 ;
    wire new_AGEMA_signal_1300 ;
    wire new_AGEMA_signal_1301 ;
    wire new_AGEMA_signal_1302 ;
    wire new_AGEMA_signal_1303 ;
    wire new_AGEMA_signal_1304 ;
    wire new_AGEMA_signal_1305 ;
    wire new_AGEMA_signal_1306 ;
    wire new_AGEMA_signal_1307 ;
    wire new_AGEMA_signal_1308 ;
    wire new_AGEMA_signal_1309 ;
    wire new_AGEMA_signal_1310 ;
    wire new_AGEMA_signal_1311 ;
    wire new_AGEMA_signal_1312 ;
    wire new_AGEMA_signal_1313 ;
    wire new_AGEMA_signal_1314 ;
    wire new_AGEMA_signal_1315 ;
    wire new_AGEMA_signal_1316 ;
    wire new_AGEMA_signal_1317 ;
    wire new_AGEMA_signal_1318 ;
    wire new_AGEMA_signal_1319 ;
    wire new_AGEMA_signal_1320 ;
    wire new_AGEMA_signal_1321 ;
    wire new_AGEMA_signal_1322 ;
    wire new_AGEMA_signal_1323 ;
    wire new_AGEMA_signal_1324 ;
    wire new_AGEMA_signal_1325 ;
    wire new_AGEMA_signal_1326 ;
    wire new_AGEMA_signal_1327 ;
    wire new_AGEMA_signal_1328 ;
    wire new_AGEMA_signal_1329 ;
    wire new_AGEMA_signal_1330 ;
    wire new_AGEMA_signal_1331 ;
    wire new_AGEMA_signal_1332 ;
    wire new_AGEMA_signal_1333 ;
    wire new_AGEMA_signal_1334 ;
    wire new_AGEMA_signal_1335 ;
    wire new_AGEMA_signal_1336 ;
    wire new_AGEMA_signal_1337 ;
    wire new_AGEMA_signal_1338 ;
    wire new_AGEMA_signal_1339 ;
    wire new_AGEMA_signal_1340 ;
    wire new_AGEMA_signal_1341 ;
    wire new_AGEMA_signal_1342 ;
    wire new_AGEMA_signal_1343 ;
    wire new_AGEMA_signal_1345 ;
    wire new_AGEMA_signal_1347 ;
    wire new_AGEMA_signal_1349 ;
    wire new_AGEMA_signal_1351 ;
    wire new_AGEMA_signal_1353 ;
    wire new_AGEMA_signal_1355 ;
    wire new_AGEMA_signal_1357 ;
    wire new_AGEMA_signal_1359 ;
    wire new_AGEMA_signal_1361 ;
    wire new_AGEMA_signal_1363 ;
    wire new_AGEMA_signal_1365 ;
    wire new_AGEMA_signal_1367 ;
    wire new_AGEMA_signal_1369 ;
    wire new_AGEMA_signal_1371 ;
    wire new_AGEMA_signal_1373 ;
    wire new_AGEMA_signal_1375 ;
    wire new_AGEMA_signal_1377 ;
    wire new_AGEMA_signal_1379 ;
    wire new_AGEMA_signal_1381 ;
    wire new_AGEMA_signal_1383 ;
    wire new_AGEMA_signal_1385 ;
    wire new_AGEMA_signal_1387 ;
    wire new_AGEMA_signal_1389 ;
    wire new_AGEMA_signal_1391 ;
    wire new_AGEMA_signal_1393 ;
    wire new_AGEMA_signal_1395 ;
    wire new_AGEMA_signal_1397 ;
    wire new_AGEMA_signal_1399 ;
    wire new_AGEMA_signal_1401 ;
    wire new_AGEMA_signal_1403 ;
    wire new_AGEMA_signal_1405 ;
    wire new_AGEMA_signal_1407 ;
    wire new_AGEMA_signal_1409 ;
    wire new_AGEMA_signal_1411 ;
    wire new_AGEMA_signal_1413 ;
    wire new_AGEMA_signal_1415 ;
    wire new_AGEMA_signal_1417 ;
    wire new_AGEMA_signal_1419 ;
    wire new_AGEMA_signal_1421 ;
    wire new_AGEMA_signal_1423 ;
    wire new_AGEMA_signal_1425 ;
    wire new_AGEMA_signal_1427 ;
    wire new_AGEMA_signal_1429 ;
    wire new_AGEMA_signal_1431 ;
    wire new_AGEMA_signal_1433 ;
    wire new_AGEMA_signal_1435 ;
    wire new_AGEMA_signal_1437 ;
    wire new_AGEMA_signal_1439 ;
    wire clk_gated ;

    /* cells in depth 0 */
    LUT6 #( .INIT ( 64'h0000001000000000 ) ) \GND_3_o_roundconstant[5]_equal_1_o<5>1 ( .I0 (\LED_128_Instance/roundconstant [5]), .I1 (\LED_128_Instance/roundconstant [4]), .I2 (\LED_128_Instance/roundconstant [3]), .I3 (\LED_128_Instance/roundconstant [2]), .I4 (\LED_128_Instance/roundconstant [1]), .I5 (\LED_128_Instance/roundconstant [0]), .O (\LED_128_Instance/roundconstant_001001 ) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[9].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[73], IN_key_s0[73]}), .I1 ({IN_key_s1[9], IN_key_s0[9]}), .I2 ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[8].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[72], IN_key_s0[72]}), .I1 ({IN_key_s1[8], IN_key_s0[8]}), .I2 ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[7].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[71], IN_key_s0[71]}), .I1 ({IN_key_s1[7], IN_key_s0[7]}), .I2 ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[63].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[127], IN_key_s0[127]}), .I1 ({IN_key_s1[63], IN_key_s0[63]}), .I2 ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[62].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[126], IN_key_s0[126]}), .I1 ({IN_key_s1[62], IN_key_s0[62]}), .I2 ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[61].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[125], IN_key_s0[125]}), .I1 ({IN_key_s1[61], IN_key_s0[61]}), .I2 ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[60].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[124], IN_key_s0[124]}), .I1 ({IN_key_s1[60], IN_key_s0[60]}), .I2 ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[59].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[123], IN_key_s0[123]}), .I1 ({IN_key_s1[59], IN_key_s0[59]}), .I2 ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[58].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[122], IN_key_s0[122]}), .I1 ({IN_key_s1[58], IN_key_s0[58]}), .I2 ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[57].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[121], IN_key_s0[121]}), .I1 ({IN_key_s1[57], IN_key_s0[57]}), .I2 ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[56].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[120], IN_key_s0[120]}), .I1 ({IN_key_s1[56], IN_key_s0[56]}), .I2 ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[55].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[119], IN_key_s0[119]}), .I1 ({IN_key_s1[55], IN_key_s0[55]}), .I2 ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[51].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[115], IN_key_s0[115]}), .I1 ({IN_key_s1[51], IN_key_s0[51]}), .I2 ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[50].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[114], IN_key_s0[114]}), .I1 ({IN_key_s1[50], IN_key_s0[50]}), .I2 ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[47].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[111], IN_key_s0[111]}), .I1 ({IN_key_s1[47], IN_key_s0[47]}), .I2 ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[46].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[110], IN_key_s0[110]}), .I1 ({IN_key_s1[46], IN_key_s0[46]}), .I2 ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[45].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[109], IN_key_s0[109]}), .I1 ({IN_key_s1[45], IN_key_s0[45]}), .I2 ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[44].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[108], IN_key_s0[108]}), .I1 ({IN_key_s1[44], IN_key_s0[44]}), .I2 ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[43].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[107], IN_key_s0[107]}), .I1 ({IN_key_s1[43], IN_key_s0[43]}), .I2 ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[42].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[106], IN_key_s0[106]}), .I1 ({IN_key_s1[42], IN_key_s0[42]}), .I2 ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[41].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[105], IN_key_s0[105]}), .I1 ({IN_key_s1[41], IN_key_s0[41]}), .I2 ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[40].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[104], IN_key_s0[104]}), .I1 ({IN_key_s1[40], IN_key_s0[40]}), .I2 ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[39].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[103], IN_key_s0[103]}), .I1 ({IN_key_s1[39], IN_key_s0[39]}), .I2 ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[35].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[99], IN_key_s0[99]}), .I1 ({IN_key_s1[35], IN_key_s0[35]}), .I2 ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[34].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[98], IN_key_s0[98]}), .I1 ({IN_key_s1[34], IN_key_s0[34]}), .I2 ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[32].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[96], IN_key_s0[96]}), .I1 ({IN_key_s1[32], IN_key_s0[32]}), .I2 ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[31].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[95], IN_key_s0[95]}), .I1 ({IN_key_s1[31], IN_key_s0[31]}), .I2 ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[30].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[94], IN_key_s0[94]}), .I1 ({IN_key_s1[30], IN_key_s0[30]}), .I2 ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[2].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[66], IN_key_s0[66]}), .I1 ({IN_key_s1[2], IN_key_s0[2]}), .I2 ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[29].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[93], IN_key_s0[93]}), .I1 ({IN_key_s1[29], IN_key_s0[29]}), .I2 ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[28].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[92], IN_key_s0[92]}), .I1 ({IN_key_s1[28], IN_key_s0[28]}), .I2 ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[27].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[91], IN_key_s0[91]}), .I1 ({IN_key_s1[27], IN_key_s0[27]}), .I2 ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[26].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[90], IN_key_s0[90]}), .I1 ({IN_key_s1[26], IN_key_s0[26]}), .I2 ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[25].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[89], IN_key_s0[89]}), .I1 ({IN_key_s1[25], IN_key_s0[25]}), .I2 ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[24].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[88], IN_key_s0[88]}), .I1 ({IN_key_s1[24], IN_key_s0[24]}), .I2 ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[23].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[87], IN_key_s0[87]}), .I1 ({IN_key_s1[23], IN_key_s0[23]}), .I2 ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[1].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[65], IN_key_s0[65]}), .I1 ({IN_key_s1[1], IN_key_s0[1]}), .I2 ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[18].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[82], IN_key_s0[82]}), .I1 ({IN_key_s1[18], IN_key_s0[18]}), .I2 ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[17].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[81], IN_key_s0[81]}), .I1 ({IN_key_s1[17], IN_key_s0[17]}), .I2 ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[15].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[79], IN_key_s0[79]}), .I1 ({IN_key_s1[15], IN_key_s0[15]}), .I2 ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[14].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[78], IN_key_s0[78]}), .I1 ({IN_key_s1[14], IN_key_s0[14]}), .I2 ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[13].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[77], IN_key_s0[77]}), .I1 ({IN_key_s1[13], IN_key_s0[13]}), .I2 ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[12].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[76], IN_key_s0[76]}), .I1 ({IN_key_s1[12], IN_key_s0[12]}), .I2 ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[11].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[75], IN_key_s0[75]}), .I1 ({IN_key_s1[11], IN_key_s0[11]}), .I2 ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[10].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[74], IN_key_s0[74]}), .I1 ({IN_key_s1[10], IN_key_s0[10]}), .I2 ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h3CF05AF0 ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h3CF05AF0 ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[0].mux_inst/Mmux_Q11 ( .I0 ({IN_key_s1[64], IN_key_s0[64]}), .I1 ({IN_key_s1[0], IN_key_s0[0]}), .I2 ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[6].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[6], IN_key_s0[6]}), .I3 ({IN_key_s1[70], IN_key_s0[70]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1049, \LED_128_Instance/addroundkey_out [6]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[5].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[5], IN_key_s0[5]}), .I3 ({IN_key_s1[69], IN_key_s0[69]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1053, \LED_128_Instance/addroundkey_out [5]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[54].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[54], IN_key_s0[54]}), .I3 ({IN_key_s1[118], IN_key_s0[118]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1057, \LED_128_Instance/addroundkey_out [54]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[53].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[53], IN_key_s0[53]}), .I3 ({IN_key_s1[117], IN_key_s0[117]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1061, \LED_128_Instance/addroundkey_out [53]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[52].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[52], IN_key_s0[52]}), .I3 ({IN_key_s1[116], IN_key_s0[116]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1065, \LED_128_Instance/addroundkey_out [52]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[4].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[4], IN_key_s0[4]}), .I3 ({IN_key_s1[68], IN_key_s0[68]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1069, \LED_128_Instance/addroundkey_out [4]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[49].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[49], IN_key_s0[49]}), .I3 ({IN_key_s1[113], IN_key_s0[113]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1073, \LED_128_Instance/addroundkey_out [49]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[48].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[48], IN_key_s0[48]}), .I3 ({IN_key_s1[112], IN_key_s0[112]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1077, \LED_128_Instance/addroundkey_out [48]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[3].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[3], IN_key_s0[3]}), .I3 ({IN_key_s1[67], IN_key_s0[67]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1081, \LED_128_Instance/addroundkey_out [3]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[38].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[38], IN_key_s0[38]}), .I3 ({IN_key_s1[102], IN_key_s0[102]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1085, \LED_128_Instance/addroundkey_out [38]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[37].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[37], IN_key_s0[37]}), .I3 ({IN_key_s1[101], IN_key_s0[101]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1089, \LED_128_Instance/addroundkey_out [37]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[36].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[36], IN_key_s0[36]}), .I3 ({IN_key_s1[100], IN_key_s0[100]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1093, \LED_128_Instance/addroundkey_out [36]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[33].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[33], IN_key_s0[33]}), .I3 ({IN_key_s1[97], IN_key_s0[97]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1097, \LED_128_Instance/addroundkey_out [33]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[22].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[22], IN_key_s0[22]}), .I3 ({IN_key_s1[86], IN_key_s0[86]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1101, \LED_128_Instance/addroundkey_out [22]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[21].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[21], IN_key_s0[21]}), .I3 ({IN_key_s1[85], IN_key_s0[85]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1105, \LED_128_Instance/addroundkey_out [21]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[20].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[20], IN_key_s0[20]}), .I3 ({IN_key_s1[84], IN_key_s0[84]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1109, \LED_128_Instance/addroundkey_out [20]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[19].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[19], IN_key_s0[19]}), .I3 ({IN_key_s1[83], IN_key_s0[83]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1113, \LED_128_Instance/addroundkey_out [19]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h596AAAAA ) , .MASK ( 5'b10010 ), .INIT2 ( 32'h596AAAAA ) ) \LED_128_Instance/MUX_addroundkey_out/gen_mux[16].mux_inst/Mmux_Q11 ( .I0 ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .I1 ({1'b0, \LED_128_Instance/addkey1_265 }), .I2 ({IN_key_s1[16], IN_key_s0[16]}), .I3 ({IN_key_s1[80], IN_key_s0[80]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .O ({new_AGEMA_signal_1117, \LED_128_Instance/addroundkey_out [16]}) ) ;
    LUT4 #( .INIT ( 16'h8001 ) ) \LED_128_Instance/addkey1 ( .I0 (\LED_128_Instance/ks [0]), .I1 (\LED_128_Instance/ks [1]), .I2 (\LED_128_Instance/ks [2]), .I3 (\LED_128_Instance/ks [3]), .O (\LED_128_Instance/addkey ) ) ;
    LUT4 #( .INIT ( 16'h0001 ) ) \LED_128_Instance/addkey21 ( .I0 (\LED_128_Instance/ks [3]), .I1 (\LED_128_Instance/ks [2]), .I2 (\LED_128_Instance/ks [1]), .I3 (\LED_128_Instance/ks [0]), .O (\LED_128_Instance/addkey1_265 ) ) ;
    LUT2 #( .INIT ( 4'h9 ) ) \LED_128_Instance/Mxor_roundconstant[5]_roundconstant[4]_XOR_7_o_xo<0>1 ( .I0 (\LED_128_Instance/roundconstant [4]), .I1 (\LED_128_Instance/roundconstant [5]), .O (\LED_128_Instance/roundconstant[5]_roundconstant[4]_XOR_7_o ) ) ;
    LUT2 #( .INIT ( 4'hE ) ) internal_done_glue_set ( .I0 (OUT_done), .I1 (\LED_128_Instance/roundconstant_001001 ), .O (internal_done_glue_set_843) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<3:0>_3_xo<0>1 ( .I0 ({IN_key_s1[3], IN_key_s0[3]}), .I1 ({IN_key_s1[67], IN_key_s0[67]}), .I2 ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<35:32>_1_xo<0>1 ( .I0 ({IN_key_s1[33], IN_key_s0[33]}), .I1 ({IN_key_s1[97], IN_key_s0[97]}), .I2 ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<19:16>_3_xo<0>1 ( .I0 ({IN_key_s1[19], IN_key_s0[19]}), .I1 ({IN_key_s1[83], IN_key_s0[83]}), .I2 ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<19:16>_0_xo<0>1 ( .I0 ({IN_key_s1[16], IN_key_s0[16]}), .I1 ({IN_key_s1[80], IN_key_s0[80]}), .I2 ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<38:36>_2_xo<0>1 ( .I0 ({IN_key_s1[38], IN_key_s0[38]}), .I1 ({IN_key_s1[102], IN_key_s0[102]}), .I2 ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [5]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<38:36>_1_xo<0>1 ( .I0 ({IN_key_s1[37], IN_key_s0[37]}), .I1 ({IN_key_s1[101], IN_key_s0[101]}), .I2 ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [4]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<38:36>_0_xo<0>1 ( .I0 ({IN_key_s1[36], IN_key_s0[36]}), .I1 ({IN_key_s1[100], IN_key_s0[100]}), .I2 ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [3]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<6:4>_2_xo<0>1 ( .I0 ({IN_key_s1[6], IN_key_s0[6]}), .I1 ({IN_key_s1[70], IN_key_s0[70]}), .I2 ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [5]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<6:4>_1_xo<0>1 ( .I0 ({IN_key_s1[5], IN_key_s0[5]}), .I1 ({IN_key_s1[69], IN_key_s0[69]}), .I2 ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [4]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<6:4>_0_xo<0>1 ( .I0 ({IN_key_s1[4], IN_key_s0[4]}), .I1 ({IN_key_s1[68], IN_key_s0[68]}), .I2 ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [3]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<51:48>_1_xo<0>1 ( .I0 ({IN_key_s1[49], IN_key_s0[49]}), .I1 ({IN_key_s1[113], IN_key_s0[113]}), .I2 ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hA50FC30F ) , .MASK ( 5'b11000 ), .INIT2 ( 32'h5AF03CF0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<51:48>_0_xo<0>1 ( .I0 ({IN_key_s1[48], IN_key_s0[48]}), .I1 ({IN_key_s1[112], IN_key_s0[112]}), .I2 ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}), .I3 ({1'b0, \LED_128_Instance/addkey }), .I4 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<54:52>_2_xo<0>1 ( .I0 ({IN_key_s1[54], IN_key_s0[54]}), .I1 ({IN_key_s1[118], IN_key_s0[118]}), .I2 ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [2]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<54:52>_1_xo<0>1 ( .I0 ({IN_key_s1[53], IN_key_s0[53]}), .I1 ({IN_key_s1[117], IN_key_s0[117]}), .I2 ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [1]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<54:52>_0_xo<0>1 ( .I0 ({IN_key_s1[52], IN_key_s0[52]}), .I1 ({IN_key_s1[116], IN_key_s0[116]}), .I2 ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [0]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<22:20>_2_xo<0>1 ( .I0 ({IN_key_s1[22], IN_key_s0[22]}), .I1 ({IN_key_s1[86], IN_key_s0[86]}), .I2 ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [2]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<22:20>_1_xo<0>1 ( .I0 ({IN_key_s1[21], IN_key_s0[21]}), .I1 ({IN_key_s1[85], IN_key_s0[85]}), .I2 ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [1]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'hA55A0FF0C33C0FF0 ) , .MASK ( 6'b111000 ), .INIT2 ( 64'h5A5AF0F03C3CF0F0 ) ) \LED_128_Instance/AddConstants_instance/Mxor_OUT_cipherstate<22:20>_0_xo<0>1 ( .I0 ({IN_key_s1[20], IN_key_s0[20]}), .I1 ({IN_key_s1[84], IN_key_s0[84]}), .I2 ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}), .I3 ({1'b0, \LED_128_Instance/roundconstant [0]}), .I4 ({1'b0, \LED_128_Instance/addkey }), .I5 ({1'b0, \LED_128_Instance/addkey1_265 }), .O ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}) ) ;
    INV \LED_128_Instance/ks[3]_INV_6_o1_INV_0 ( .I (\LED_128_Instance/ks [3]), .O (\LED_128_Instance/ks[3]_INV_6_o ) ) ;
    ClockGatingController #(2) ClockGatingInst ( .clk (CLK), .rst (IN_reset), .GatedClk (clk_gated), .Synch (Synch) ) ;

    /* cells in depth 1 */
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[0].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I3 ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}), .clk (CLK), .r ({Fresh[15], Fresh[14], Fresh[13], Fresh[12], Fresh[11], Fresh[10], Fresh[9], Fresh[8], Fresh[7], Fresh[6], Fresh[5], Fresh[4], Fresh[3], Fresh[2], Fresh[1], Fresh[0]}), .O ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[0].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I3 ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}), .clk (CLK), .r ({Fresh[31], Fresh[30], Fresh[29], Fresh[28], Fresh[27], Fresh[26], Fresh[25], Fresh[24], Fresh[23], Fresh[22], Fresh[21], Fresh[20], Fresh[19], Fresh[18], Fresh[17], Fresh[16]}), .O ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[0].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I3 ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}), .clk (CLK), .r ({Fresh[47], Fresh[46], Fresh[45], Fresh[44], Fresh[43], Fresh[42], Fresh[41], Fresh[40], Fresh[39], Fresh[38], Fresh[37], Fresh[36], Fresh[35], Fresh[34], Fresh[33], Fresh[32]}), .O ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[0].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I3 ({new_AGEMA_signal_1118, \LED_128_Instance/addconst_out [3]}), .clk (CLK), .r ({Fresh[63], Fresh[62], Fresh[61], Fresh[60], Fresh[59], Fresh[58], Fresh[57], Fresh[56], Fresh[55], Fresh[54], Fresh[53], Fresh[52], Fresh[51], Fresh[50], Fresh[49], Fresh[48]}), .O ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[1].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}), .I1 ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}), .I2 ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}), .I3 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .clk (CLK), .r ({Fresh[79], Fresh[78], Fresh[77], Fresh[76], Fresh[75], Fresh[74], Fresh[73], Fresh[72], Fresh[71], Fresh[70], Fresh[69], Fresh[68], Fresh[67], Fresh[66], Fresh[65], Fresh[64]}), .O ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[1].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}), .I1 ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}), .I2 ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}), .I3 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .clk (CLK), .r ({Fresh[95], Fresh[94], Fresh[93], Fresh[92], Fresh[91], Fresh[90], Fresh[89], Fresh[88], Fresh[87], Fresh[86], Fresh[85], Fresh[84], Fresh[83], Fresh[82], Fresh[81], Fresh[80]}), .O ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[1].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}), .I1 ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}), .I2 ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}), .I3 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .clk (CLK), .r ({Fresh[111], Fresh[110], Fresh[109], Fresh[108], Fresh[107], Fresh[106], Fresh[105], Fresh[104], Fresh[103], Fresh[102], Fresh[101], Fresh[100], Fresh[99], Fresh[98], Fresh[97], Fresh[96]}), .O ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[1].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1127, \LED_128_Instance/addconst_out [4]}), .I1 ({new_AGEMA_signal_1126, \LED_128_Instance/addconst_out [5]}), .I2 ({new_AGEMA_signal_1125, \LED_128_Instance/addconst_out [6]}), .I3 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .clk (CLK), .r ({Fresh[127], Fresh[126], Fresh[125], Fresh[124], Fresh[123], Fresh[122], Fresh[121], Fresh[120], Fresh[119], Fresh[118], Fresh[117], Fresh[116], Fresh[115], Fresh[114], Fresh[113], Fresh[112]}), .O ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[2].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I3 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .clk (CLK), .r ({Fresh[143], Fresh[142], Fresh[141], Fresh[140], Fresh[139], Fresh[138], Fresh[137], Fresh[136], Fresh[135], Fresh[134], Fresh[133], Fresh[132], Fresh[131], Fresh[130], Fresh[129], Fresh[128]}), .O ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[2].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I3 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .clk (CLK), .r ({Fresh[159], Fresh[158], Fresh[157], Fresh[156], Fresh[155], Fresh[154], Fresh[153], Fresh[152], Fresh[151], Fresh[150], Fresh[149], Fresh[148], Fresh[147], Fresh[146], Fresh[145], Fresh[144]}), .O ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[2].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I3 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .clk (CLK), .r ({Fresh[175], Fresh[174], Fresh[173], Fresh[172], Fresh[171], Fresh[170], Fresh[169], Fresh[168], Fresh[167], Fresh[166], Fresh[165], Fresh[164], Fresh[163], Fresh[162], Fresh[161], Fresh[160]}), .O ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[2].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I3 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .clk (CLK), .r ({Fresh[191], Fresh[190], Fresh[189], Fresh[188], Fresh[187], Fresh[186], Fresh[185], Fresh[184], Fresh[183], Fresh[182], Fresh[181], Fresh[180], Fresh[179], Fresh[178], Fresh[177], Fresh[176]}), .O ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[3].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I3 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .clk (CLK), .r ({Fresh[207], Fresh[206], Fresh[205], Fresh[204], Fresh[203], Fresh[202], Fresh[201], Fresh[200], Fresh[199], Fresh[198], Fresh[197], Fresh[196], Fresh[195], Fresh[194], Fresh[193], Fresh[192]}), .O ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[3].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I3 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .clk (CLK), .r ({Fresh[223], Fresh[222], Fresh[221], Fresh[220], Fresh[219], Fresh[218], Fresh[217], Fresh[216], Fresh[215], Fresh[214], Fresh[213], Fresh[212], Fresh[211], Fresh[210], Fresh[209], Fresh[208]}), .O ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[3].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I3 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .clk (CLK), .r ({Fresh[239], Fresh[238], Fresh[237], Fresh[236], Fresh[235], Fresh[234], Fresh[233], Fresh[232], Fresh[231], Fresh[230], Fresh[229], Fresh[228], Fresh[227], Fresh[226], Fresh[225], Fresh[224]}), .O ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[3].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I3 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .clk (CLK), .r ({Fresh[255], Fresh[254], Fresh[253], Fresh[252], Fresh[251], Fresh[250], Fresh[249], Fresh[248], Fresh[247], Fresh[246], Fresh[245], Fresh[244], Fresh[243], Fresh[242], Fresh[241], Fresh[240]}), .O ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[4].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I3 ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}), .clk (CLK), .r ({Fresh[271], Fresh[270], Fresh[269], Fresh[268], Fresh[267], Fresh[266], Fresh[265], Fresh[264], Fresh[263], Fresh[262], Fresh[261], Fresh[260], Fresh[259], Fresh[258], Fresh[257], Fresh[256]}), .O ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[4].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I3 ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}), .clk (CLK), .r ({Fresh[287], Fresh[286], Fresh[285], Fresh[284], Fresh[283], Fresh[282], Fresh[281], Fresh[280], Fresh[279], Fresh[278], Fresh[277], Fresh[276], Fresh[275], Fresh[274], Fresh[273], Fresh[272]}), .O ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[4].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I3 ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}), .clk (CLK), .r ({Fresh[303], Fresh[302], Fresh[301], Fresh[300], Fresh[299], Fresh[298], Fresh[297], Fresh[296], Fresh[295], Fresh[294], Fresh[293], Fresh[292], Fresh[291], Fresh[290], Fresh[289], Fresh[288]}), .O ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[4].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1121, \LED_128_Instance/addconst_out [16]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I3 ({new_AGEMA_signal_1120, \LED_128_Instance/addconst_out [19]}), .clk (CLK), .r ({Fresh[319], Fresh[318], Fresh[317], Fresh[316], Fresh[315], Fresh[314], Fresh[313], Fresh[312], Fresh[311], Fresh[310], Fresh[309], Fresh[308], Fresh[307], Fresh[306], Fresh[305], Fresh[304]}), .O ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[5].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}), .I1 ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}), .I2 ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}), .I3 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .clk (CLK), .r ({Fresh[335], Fresh[334], Fresh[333], Fresh[332], Fresh[331], Fresh[330], Fresh[329], Fresh[328], Fresh[327], Fresh[326], Fresh[325], Fresh[324], Fresh[323], Fresh[322], Fresh[321], Fresh[320]}), .O ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[5].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}), .I1 ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}), .I2 ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}), .I3 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .clk (CLK), .r ({Fresh[351], Fresh[350], Fresh[349], Fresh[348], Fresh[347], Fresh[346], Fresh[345], Fresh[344], Fresh[343], Fresh[342], Fresh[341], Fresh[340], Fresh[339], Fresh[338], Fresh[337], Fresh[336]}), .O ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[5].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}), .I1 ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}), .I2 ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}), .I3 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .clk (CLK), .r ({Fresh[367], Fresh[366], Fresh[365], Fresh[364], Fresh[363], Fresh[362], Fresh[361], Fresh[360], Fresh[359], Fresh[358], Fresh[357], Fresh[356], Fresh[355], Fresh[354], Fresh[353], Fresh[352]}), .O ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[5].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1135, \LED_128_Instance/addconst_out [20]}), .I1 ({new_AGEMA_signal_1134, \LED_128_Instance/addconst_out [21]}), .I2 ({new_AGEMA_signal_1133, \LED_128_Instance/addconst_out [22]}), .I3 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .clk (CLK), .r ({Fresh[383], Fresh[382], Fresh[381], Fresh[380], Fresh[379], Fresh[378], Fresh[377], Fresh[376], Fresh[375], Fresh[374], Fresh[373], Fresh[372], Fresh[371], Fresh[370], Fresh[369], Fresh[368]}), .O ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[6].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I3 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .clk (CLK), .r ({Fresh[399], Fresh[398], Fresh[397], Fresh[396], Fresh[395], Fresh[394], Fresh[393], Fresh[392], Fresh[391], Fresh[390], Fresh[389], Fresh[388], Fresh[387], Fresh[386], Fresh[385], Fresh[384]}), .O ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[6].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I3 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .clk (CLK), .r ({Fresh[415], Fresh[414], Fresh[413], Fresh[412], Fresh[411], Fresh[410], Fresh[409], Fresh[408], Fresh[407], Fresh[406], Fresh[405], Fresh[404], Fresh[403], Fresh[402], Fresh[401], Fresh[400]}), .O ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[6].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I3 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .clk (CLK), .r ({Fresh[431], Fresh[430], Fresh[429], Fresh[428], Fresh[427], Fresh[426], Fresh[425], Fresh[424], Fresh[423], Fresh[422], Fresh[421], Fresh[420], Fresh[419], Fresh[418], Fresh[417], Fresh[416]}), .O ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[6].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I3 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .clk (CLK), .r ({Fresh[447], Fresh[446], Fresh[445], Fresh[444], Fresh[443], Fresh[442], Fresh[441], Fresh[440], Fresh[439], Fresh[438], Fresh[437], Fresh[436], Fresh[435], Fresh[434], Fresh[433], Fresh[432]}), .O ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[7].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I3 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .clk (CLK), .r ({Fresh[463], Fresh[462], Fresh[461], Fresh[460], Fresh[459], Fresh[458], Fresh[457], Fresh[456], Fresh[455], Fresh[454], Fresh[453], Fresh[452], Fresh[451], Fresh[450], Fresh[449], Fresh[448]}), .O ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[7].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I3 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .clk (CLK), .r ({Fresh[479], Fresh[478], Fresh[477], Fresh[476], Fresh[475], Fresh[474], Fresh[473], Fresh[472], Fresh[471], Fresh[470], Fresh[469], Fresh[468], Fresh[467], Fresh[466], Fresh[465], Fresh[464]}), .O ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[7].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I3 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .clk (CLK), .r ({Fresh[495], Fresh[494], Fresh[493], Fresh[492], Fresh[491], Fresh[490], Fresh[489], Fresh[488], Fresh[487], Fresh[486], Fresh[485], Fresh[484], Fresh[483], Fresh[482], Fresh[481], Fresh[480]}), .O ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[7].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I3 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .clk (CLK), .r ({Fresh[511], Fresh[510], Fresh[509], Fresh[508], Fresh[507], Fresh[506], Fresh[505], Fresh[504], Fresh[503], Fresh[502], Fresh[501], Fresh[500], Fresh[499], Fresh[498], Fresh[497], Fresh[496]}), .O ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[8].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I1 ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}), .I2 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I3 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .clk (CLK), .r ({Fresh[527], Fresh[526], Fresh[525], Fresh[524], Fresh[523], Fresh[522], Fresh[521], Fresh[520], Fresh[519], Fresh[518], Fresh[517], Fresh[516], Fresh[515], Fresh[514], Fresh[513], Fresh[512]}), .O ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[8].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I1 ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}), .I2 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I3 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .clk (CLK), .r ({Fresh[543], Fresh[542], Fresh[541], Fresh[540], Fresh[539], Fresh[538], Fresh[537], Fresh[536], Fresh[535], Fresh[534], Fresh[533], Fresh[532], Fresh[531], Fresh[530], Fresh[529], Fresh[528]}), .O ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[8].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I1 ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}), .I2 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I3 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .clk (CLK), .r ({Fresh[559], Fresh[558], Fresh[557], Fresh[556], Fresh[555], Fresh[554], Fresh[553], Fresh[552], Fresh[551], Fresh[550], Fresh[549], Fresh[548], Fresh[547], Fresh[546], Fresh[545], Fresh[544]}), .O ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[8].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I1 ({new_AGEMA_signal_1119, \LED_128_Instance/addconst_out [33]}), .I2 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I3 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .clk (CLK), .r ({Fresh[575], Fresh[574], Fresh[573], Fresh[572], Fresh[571], Fresh[570], Fresh[569], Fresh[568], Fresh[567], Fresh[566], Fresh[565], Fresh[564], Fresh[563], Fresh[562], Fresh[561], Fresh[560]}), .O ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[9].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}), .I1 ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}), .I2 ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}), .I3 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .clk (CLK), .r ({Fresh[591], Fresh[590], Fresh[589], Fresh[588], Fresh[587], Fresh[586], Fresh[585], Fresh[584], Fresh[583], Fresh[582], Fresh[581], Fresh[580], Fresh[579], Fresh[578], Fresh[577], Fresh[576]}), .O ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[9].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}), .I1 ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}), .I2 ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}), .I3 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .clk (CLK), .r ({Fresh[607], Fresh[606], Fresh[605], Fresh[604], Fresh[603], Fresh[602], Fresh[601], Fresh[600], Fresh[599], Fresh[598], Fresh[597], Fresh[596], Fresh[595], Fresh[594], Fresh[593], Fresh[592]}), .O ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[9].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}), .I1 ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}), .I2 ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}), .I3 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .clk (CLK), .r ({Fresh[623], Fresh[622], Fresh[621], Fresh[620], Fresh[619], Fresh[618], Fresh[617], Fresh[616], Fresh[615], Fresh[614], Fresh[613], Fresh[612], Fresh[611], Fresh[610], Fresh[609], Fresh[608]}), .O ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[9].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1124, \LED_128_Instance/addconst_out [36]}), .I1 ({new_AGEMA_signal_1123, \LED_128_Instance/addconst_out [37]}), .I2 ({new_AGEMA_signal_1122, \LED_128_Instance/addconst_out [38]}), .I3 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .clk (CLK), .r ({Fresh[639], Fresh[638], Fresh[637], Fresh[636], Fresh[635], Fresh[634], Fresh[633], Fresh[632], Fresh[631], Fresh[630], Fresh[629], Fresh[628], Fresh[627], Fresh[626], Fresh[625], Fresh[624]}), .O ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[10].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I3 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .clk (CLK), .r ({Fresh[655], Fresh[654], Fresh[653], Fresh[652], Fresh[651], Fresh[650], Fresh[649], Fresh[648], Fresh[647], Fresh[646], Fresh[645], Fresh[644], Fresh[643], Fresh[642], Fresh[641], Fresh[640]}), .O ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[10].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I3 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .clk (CLK), .r ({Fresh[671], Fresh[670], Fresh[669], Fresh[668], Fresh[667], Fresh[666], Fresh[665], Fresh[664], Fresh[663], Fresh[662], Fresh[661], Fresh[660], Fresh[659], Fresh[658], Fresh[657], Fresh[656]}), .O ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[10].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I3 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .clk (CLK), .r ({Fresh[687], Fresh[686], Fresh[685], Fresh[684], Fresh[683], Fresh[682], Fresh[681], Fresh[680], Fresh[679], Fresh[678], Fresh[677], Fresh[676], Fresh[675], Fresh[674], Fresh[673], Fresh[672]}), .O ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[10].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I3 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .clk (CLK), .r ({Fresh[703], Fresh[702], Fresh[701], Fresh[700], Fresh[699], Fresh[698], Fresh[697], Fresh[696], Fresh[695], Fresh[694], Fresh[693], Fresh[692], Fresh[691], Fresh[690], Fresh[689], Fresh[688]}), .O ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[11].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I3 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .clk (CLK), .r ({Fresh[719], Fresh[718], Fresh[717], Fresh[716], Fresh[715], Fresh[714], Fresh[713], Fresh[712], Fresh[711], Fresh[710], Fresh[709], Fresh[708], Fresh[707], Fresh[706], Fresh[705], Fresh[704]}), .O ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[11].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I3 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .clk (CLK), .r ({Fresh[735], Fresh[734], Fresh[733], Fresh[732], Fresh[731], Fresh[730], Fresh[729], Fresh[728], Fresh[727], Fresh[726], Fresh[725], Fresh[724], Fresh[723], Fresh[722], Fresh[721], Fresh[720]}), .O ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[11].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I3 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .clk (CLK), .r ({Fresh[751], Fresh[750], Fresh[749], Fresh[748], Fresh[747], Fresh[746], Fresh[745], Fresh[744], Fresh[743], Fresh[742], Fresh[741], Fresh[740], Fresh[739], Fresh[738], Fresh[737], Fresh[736]}), .O ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[11].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I3 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .clk (CLK), .r ({Fresh[767], Fresh[766], Fresh[765], Fresh[764], Fresh[763], Fresh[762], Fresh[761], Fresh[760], Fresh[759], Fresh[758], Fresh[757], Fresh[756], Fresh[755], Fresh[754], Fresh[753], Fresh[752]}), .O ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[12].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}), .I1 ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}), .I2 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I3 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .clk (CLK), .r ({Fresh[783], Fresh[782], Fresh[781], Fresh[780], Fresh[779], Fresh[778], Fresh[777], Fresh[776], Fresh[775], Fresh[774], Fresh[773], Fresh[772], Fresh[771], Fresh[770], Fresh[769], Fresh[768]}), .O ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[12].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}), .I1 ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}), .I2 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I3 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .clk (CLK), .r ({Fresh[799], Fresh[798], Fresh[797], Fresh[796], Fresh[795], Fresh[794], Fresh[793], Fresh[792], Fresh[791], Fresh[790], Fresh[789], Fresh[788], Fresh[787], Fresh[786], Fresh[785], Fresh[784]}), .O ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[12].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}), .I1 ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}), .I2 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I3 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .clk (CLK), .r ({Fresh[815], Fresh[814], Fresh[813], Fresh[812], Fresh[811], Fresh[810], Fresh[809], Fresh[808], Fresh[807], Fresh[806], Fresh[805], Fresh[804], Fresh[803], Fresh[802], Fresh[801], Fresh[800]}), .O ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[12].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1129, \LED_128_Instance/addconst_out [48]}), .I1 ({new_AGEMA_signal_1128, \LED_128_Instance/addconst_out [49]}), .I2 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I3 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .clk (CLK), .r ({Fresh[831], Fresh[830], Fresh[829], Fresh[828], Fresh[827], Fresh[826], Fresh[825], Fresh[824], Fresh[823], Fresh[822], Fresh[821], Fresh[820], Fresh[819], Fresh[818], Fresh[817], Fresh[816]}), .O ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[13].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}), .I1 ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}), .I2 ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}), .I3 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .clk (CLK), .r ({Fresh[847], Fresh[846], Fresh[845], Fresh[844], Fresh[843], Fresh[842], Fresh[841], Fresh[840], Fresh[839], Fresh[838], Fresh[837], Fresh[836], Fresh[835], Fresh[834], Fresh[833], Fresh[832]}), .O ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[13].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}), .I1 ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}), .I2 ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}), .I3 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .clk (CLK), .r ({Fresh[863], Fresh[862], Fresh[861], Fresh[860], Fresh[859], Fresh[858], Fresh[857], Fresh[856], Fresh[855], Fresh[854], Fresh[853], Fresh[852], Fresh[851], Fresh[850], Fresh[849], Fresh[848]}), .O ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[13].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}), .I1 ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}), .I2 ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}), .I3 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .clk (CLK), .r ({Fresh[879], Fresh[878], Fresh[877], Fresh[876], Fresh[875], Fresh[874], Fresh[873], Fresh[872], Fresh[871], Fresh[870], Fresh[869], Fresh[868], Fresh[867], Fresh[866], Fresh[865], Fresh[864]}), .O ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[13].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_1132, \LED_128_Instance/addconst_out [52]}), .I1 ({new_AGEMA_signal_1131, \LED_128_Instance/addconst_out [53]}), .I2 ({new_AGEMA_signal_1130, \LED_128_Instance/addconst_out [54]}), .I3 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .clk (CLK), .r ({Fresh[895], Fresh[894], Fresh[893], Fresh[892], Fresh[891], Fresh[890], Fresh[889], Fresh[888], Fresh[887], Fresh[886], Fresh[885], Fresh[884], Fresh[883], Fresh[882], Fresh[881], Fresh[880]}), .O ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[14].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I3 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .clk (CLK), .r ({Fresh[911], Fresh[910], Fresh[909], Fresh[908], Fresh[907], Fresh[906], Fresh[905], Fresh[904], Fresh[903], Fresh[902], Fresh[901], Fresh[900], Fresh[899], Fresh[898], Fresh[897], Fresh[896]}), .O ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[14].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I3 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .clk (CLK), .r ({Fresh[927], Fresh[926], Fresh[925], Fresh[924], Fresh[923], Fresh[922], Fresh[921], Fresh[920], Fresh[919], Fresh[918], Fresh[917], Fresh[916], Fresh[915], Fresh[914], Fresh[913], Fresh[912]}), .O ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[14].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I3 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .clk (CLK), .r ({Fresh[943], Fresh[942], Fresh[941], Fresh[940], Fresh[939], Fresh[938], Fresh[937], Fresh[936], Fresh[935], Fresh[934], Fresh[933], Fresh[932], Fresh[931], Fresh[930], Fresh[929], Fresh[928]}), .O ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[14].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I3 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .clk (CLK), .r ({Fresh[959], Fresh[958], Fresh[957], Fresh[956], Fresh[955], Fresh[954], Fresh[953], Fresh[952], Fresh[951], Fresh[950], Fresh[949], Fresh[948], Fresh[947], Fresh[946], Fresh[945], Fresh[944]}), .O ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h659A ) ) \LED_128_Instance/sub_loop[15].SBox_Instance/y_0 ( .I0 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I3 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .clk (CLK), .r ({Fresh[975], Fresh[974], Fresh[973], Fresh[972], Fresh[971], Fresh[970], Fresh[969], Fresh[968], Fresh[967], Fresh[966], Fresh[965], Fresh[964], Fresh[963], Fresh[962], Fresh[961], Fresh[960]}), .O ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'hA74C ) ) \LED_128_Instance/sub_loop[15].SBox_Instance/y_1 ( .I0 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I3 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .clk (CLK), .r ({Fresh[991], Fresh[990], Fresh[989], Fresh[988], Fresh[987], Fresh[986], Fresh[985], Fresh[984], Fresh[983], Fresh[982], Fresh[981], Fresh[980], Fresh[979], Fresh[978], Fresh[977], Fresh[976]}), .O ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h3687 ) ) \LED_128_Instance/sub_loop[15].SBox_Instance/y_2 ( .I0 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I3 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .clk (CLK), .r ({Fresh[1007], Fresh[1006], Fresh[1005], Fresh[1004], Fresh[1003], Fresh[1002], Fresh[1001], Fresh[1000], Fresh[999], Fresh[998], Fresh[997], Fresh[996], Fresh[995], Fresh[994], Fresh[993], Fresh[992]}), .O ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}) ) ;
    LUT4_GHPC #(.low_latency(1), .pipeline(0),  .INIT ( 16'h0ED9 ) ) \LED_128_Instance/sub_loop[15].SBox_Instance/y_3 ( .I0 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I3 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .clk (CLK), .r ({Fresh[1023], Fresh[1022], Fresh[1021], Fresh[1020], Fresh[1019], Fresh[1018], Fresh[1017], Fresh[1016], Fresh[1015], Fresh[1014], Fresh[1013], Fresh[1012], Fresh[1011], Fresh[1010], Fresh[1009], Fresh[1008]}), .O ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[0].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1203, \LED_128_Instance/mixcolumns_out [0]}), .I1 ({new_AGEMA_signal_1045, \LED_128_Instance/addroundkey_out [0]}), .I2 ({IN_plaintext_s1[0], IN_plaintext_s0[0]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1265, \LED_128_Instance/state [0]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[1].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1334, \LED_128_Instance/mixcolumns_out [1]}), .I1 ({new_AGEMA_signal_1009, \LED_128_Instance/addroundkey_out [1]}), .I2 ({IN_plaintext_s1[1], IN_plaintext_s0[1]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1345, \LED_128_Instance/state [1]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[2].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1200, \LED_128_Instance/mixcolumns_out [2]}), .I1 ({new_AGEMA_signal_977, \LED_128_Instance/addroundkey_out [2]}), .I2 ({IN_plaintext_s1[2], IN_plaintext_s0[2]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1267, \LED_128_Instance/state [2]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[3].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1202, \LED_128_Instance/mixcolumns_out [3]}), .I1 ({new_AGEMA_signal_1081, \LED_128_Instance/addroundkey_out [3]}), .I2 ({IN_plaintext_s1[3], IN_plaintext_s0[3]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1269, \LED_128_Instance/state [3]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[4].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1207, \LED_128_Instance/mixcolumns_out [4]}), .I1 ({new_AGEMA_signal_1069, \LED_128_Instance/addroundkey_out [4]}), .I2 ({IN_plaintext_s1[4], IN_plaintext_s0[4]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1271, \LED_128_Instance/state [4]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[5].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1336, \LED_128_Instance/mixcolumns_out [5]}), .I1 ({new_AGEMA_signal_1053, \LED_128_Instance/addroundkey_out [5]}), .I2 ({IN_plaintext_s1[5], IN_plaintext_s0[5]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1347, \LED_128_Instance/state [5]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[6].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1204, \LED_128_Instance/mixcolumns_out [6]}), .I1 ({new_AGEMA_signal_1049, \LED_128_Instance/addroundkey_out [6]}), .I2 ({IN_plaintext_s1[6], IN_plaintext_s0[6]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1273, \LED_128_Instance/state [6]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[7].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1206, \LED_128_Instance/mixcolumns_out [7]}), .I1 ({new_AGEMA_signal_873, \LED_128_Instance/addroundkey_out [7]}), .I2 ({IN_plaintext_s1[7], IN_plaintext_s0[7]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1275, \LED_128_Instance/state [7]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[8].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1210, \LED_128_Instance/mixcolumns_out [8]}), .I1 ({new_AGEMA_signal_869, \LED_128_Instance/addroundkey_out [8]}), .I2 ({IN_plaintext_s1[8], IN_plaintext_s0[8]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1277, \LED_128_Instance/state [8]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[9].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1338, \LED_128_Instance/mixcolumns_out [9]}), .I1 ({new_AGEMA_signal_865, \LED_128_Instance/addroundkey_out [9]}), .I2 ({IN_plaintext_s1[9], IN_plaintext_s0[9]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1349, \LED_128_Instance/state [9]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[10].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1209, \LED_128_Instance/mixcolumns_out [10]}), .I1 ({new_AGEMA_signal_1041, \LED_128_Instance/addroundkey_out [10]}), .I2 ({IN_plaintext_s1[10], IN_plaintext_s0[10]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1279, \LED_128_Instance/state [10]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[11].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1211, \LED_128_Instance/mixcolumns_out [11]}), .I1 ({new_AGEMA_signal_1037, \LED_128_Instance/addroundkey_out [11]}), .I2 ({IN_plaintext_s1[11], IN_plaintext_s0[11]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1281, \LED_128_Instance/state [11]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[12].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1215, \LED_128_Instance/mixcolumns_out [12]}), .I1 ({new_AGEMA_signal_1033, \LED_128_Instance/addroundkey_out [12]}), .I2 ({IN_plaintext_s1[12], IN_plaintext_s0[12]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1283, \LED_128_Instance/state [12]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[13].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1332, \LED_128_Instance/mixcolumns_out [13]}), .I1 ({new_AGEMA_signal_1029, \LED_128_Instance/addroundkey_out [13]}), .I2 ({IN_plaintext_s1[13], IN_plaintext_s0[13]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1351, \LED_128_Instance/state [13]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[14].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1213, \LED_128_Instance/mixcolumns_out [14]}), .I1 ({new_AGEMA_signal_1025, \LED_128_Instance/addroundkey_out [14]}), .I2 ({IN_plaintext_s1[14], IN_plaintext_s0[14]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1285, \LED_128_Instance/state [14]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[15].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1214, \LED_128_Instance/mixcolumns_out [15]}), .I1 ({new_AGEMA_signal_1021, \LED_128_Instance/addroundkey_out [15]}), .I2 ({IN_plaintext_s1[15], IN_plaintext_s0[15]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1287, \LED_128_Instance/state [15]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[16].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1297, \LED_128_Instance/mixcolumns_out [16]}), .I1 ({new_AGEMA_signal_1117, \LED_128_Instance/addroundkey_out [16]}), .I2 ({IN_plaintext_s1[16], IN_plaintext_s0[16]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1353, \LED_128_Instance/state [16]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[17].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1304, \LED_128_Instance/mixcolumns_out [17]}), .I1 ({new_AGEMA_signal_1017, \LED_128_Instance/addroundkey_out [17]}), .I2 ({IN_plaintext_s1[17], IN_plaintext_s0[17]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1355, \LED_128_Instance/state [17]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[18].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1340, \LED_128_Instance/mixcolumns_out [18]}), .I1 ({new_AGEMA_signal_1013, \LED_128_Instance/addroundkey_out [18]}), .I2 ({IN_plaintext_s1[18], IN_plaintext_s0[18]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1357, \LED_128_Instance/state [18]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[19].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1296, \LED_128_Instance/mixcolumns_out [19]}), .I1 ({new_AGEMA_signal_1113, \LED_128_Instance/addroundkey_out [19]}), .I2 ({IN_plaintext_s1[19], IN_plaintext_s0[19]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1359, \LED_128_Instance/state [19]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[20].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1306, \LED_128_Instance/mixcolumns_out [20]}), .I1 ({new_AGEMA_signal_1109, \LED_128_Instance/addroundkey_out [20]}), .I2 ({IN_plaintext_s1[20], IN_plaintext_s0[20]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1361, \LED_128_Instance/state [20]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[21].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1313, \LED_128_Instance/mixcolumns_out [21]}), .I1 ({new_AGEMA_signal_1105, \LED_128_Instance/addroundkey_out [21]}), .I2 ({IN_plaintext_s1[21], IN_plaintext_s0[21]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1363, \LED_128_Instance/state [21]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[22].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1341, \LED_128_Instance/mixcolumns_out [22]}), .I1 ({new_AGEMA_signal_1101, \LED_128_Instance/addroundkey_out [22]}), .I2 ({IN_plaintext_s1[22], IN_plaintext_s0[22]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1365, \LED_128_Instance/state [22]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[23].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1305, \LED_128_Instance/mixcolumns_out [23]}), .I1 ({new_AGEMA_signal_1005, \LED_128_Instance/addroundkey_out [23]}), .I2 ({IN_plaintext_s1[23], IN_plaintext_s0[23]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1367, \LED_128_Instance/state [23]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[24].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1314, \LED_128_Instance/mixcolumns_out [24]}), .I1 ({new_AGEMA_signal_1001, \LED_128_Instance/addroundkey_out [24]}), .I2 ({IN_plaintext_s1[24], IN_plaintext_s0[24]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1369, \LED_128_Instance/state [24]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[25].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1322, \LED_128_Instance/mixcolumns_out [25]}), .I1 ({new_AGEMA_signal_997, \LED_128_Instance/addroundkey_out [25]}), .I2 ({IN_plaintext_s1[25], IN_plaintext_s0[25]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1371, \LED_128_Instance/state [25]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[26].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1342, \LED_128_Instance/mixcolumns_out [26]}), .I1 ({new_AGEMA_signal_993, \LED_128_Instance/addroundkey_out [26]}), .I2 ({IN_plaintext_s1[26], IN_plaintext_s0[26]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1373, \LED_128_Instance/state [26]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[27].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1315, \LED_128_Instance/mixcolumns_out [27]}), .I1 ({new_AGEMA_signal_989, \LED_128_Instance/addroundkey_out [27]}), .I2 ({IN_plaintext_s1[27], IN_plaintext_s0[27]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1375, \LED_128_Instance/state [27]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[28].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1323, \LED_128_Instance/mixcolumns_out [28]}), .I1 ({new_AGEMA_signal_985, \LED_128_Instance/addroundkey_out [28]}), .I2 ({IN_plaintext_s1[28], IN_plaintext_s0[28]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1377, \LED_128_Instance/state [28]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[29].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1331, \LED_128_Instance/mixcolumns_out [29]}), .I1 ({new_AGEMA_signal_981, \LED_128_Instance/addroundkey_out [29]}), .I2 ({IN_plaintext_s1[29], IN_plaintext_s0[29]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1379, \LED_128_Instance/state [29]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[30].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1343, \LED_128_Instance/mixcolumns_out [30]}), .I1 ({new_AGEMA_signal_973, \LED_128_Instance/addroundkey_out [30]}), .I2 ({IN_plaintext_s1[30], IN_plaintext_s0[30]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1381, \LED_128_Instance/state [30]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[31].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1324, \LED_128_Instance/mixcolumns_out [31]}), .I1 ({new_AGEMA_signal_969, \LED_128_Instance/addroundkey_out [31]}), .I2 ({IN_plaintext_s1[31], IN_plaintext_s0[31]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1383, \LED_128_Instance/state [31]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[32].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1303, \LED_128_Instance/mixcolumns_out [32]}), .I1 ({new_AGEMA_signal_965, \LED_128_Instance/addroundkey_out [32]}), .I2 ({IN_plaintext_s1[32], IN_plaintext_s0[32]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1385, \LED_128_Instance/state [32]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[33].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1299, \LED_128_Instance/mixcolumns_out [33]}), .I1 ({new_AGEMA_signal_1097, \LED_128_Instance/addroundkey_out [33]}), .I2 ({IN_plaintext_s1[33], IN_plaintext_s0[33]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1387, \LED_128_Instance/state [33]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[34].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1302, \LED_128_Instance/mixcolumns_out [34]}), .I1 ({new_AGEMA_signal_961, \LED_128_Instance/addroundkey_out [34]}), .I2 ({IN_plaintext_s1[34], IN_plaintext_s0[34]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1389, \LED_128_Instance/state [34]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[35].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1298, \LED_128_Instance/mixcolumns_out [35]}), .I1 ({new_AGEMA_signal_957, \LED_128_Instance/addroundkey_out [35]}), .I2 ({IN_plaintext_s1[35], IN_plaintext_s0[35]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1391, \LED_128_Instance/state [35]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[36].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1312, \LED_128_Instance/mixcolumns_out [36]}), .I1 ({new_AGEMA_signal_1093, \LED_128_Instance/addroundkey_out [36]}), .I2 ({IN_plaintext_s1[36], IN_plaintext_s0[36]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1393, \LED_128_Instance/state [36]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[37].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1308, \LED_128_Instance/mixcolumns_out [37]}), .I1 ({new_AGEMA_signal_1089, \LED_128_Instance/addroundkey_out [37]}), .I2 ({IN_plaintext_s1[37], IN_plaintext_s0[37]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1395, \LED_128_Instance/state [37]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[38].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1311, \LED_128_Instance/mixcolumns_out [38]}), .I1 ({new_AGEMA_signal_1085, \LED_128_Instance/addroundkey_out [38]}), .I2 ({IN_plaintext_s1[38], IN_plaintext_s0[38]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1397, \LED_128_Instance/state [38]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[39].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1307, \LED_128_Instance/mixcolumns_out [39]}), .I1 ({new_AGEMA_signal_953, \LED_128_Instance/addroundkey_out [39]}), .I2 ({IN_plaintext_s1[39], IN_plaintext_s0[39]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1399, \LED_128_Instance/state [39]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[40].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1321, \LED_128_Instance/mixcolumns_out [40]}), .I1 ({new_AGEMA_signal_949, \LED_128_Instance/addroundkey_out [40]}), .I2 ({IN_plaintext_s1[40], IN_plaintext_s0[40]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1401, \LED_128_Instance/state [40]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[41].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1317, \LED_128_Instance/mixcolumns_out [41]}), .I1 ({new_AGEMA_signal_945, \LED_128_Instance/addroundkey_out [41]}), .I2 ({IN_plaintext_s1[41], IN_plaintext_s0[41]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1403, \LED_128_Instance/state [41]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[42].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1320, \LED_128_Instance/mixcolumns_out [42]}), .I1 ({new_AGEMA_signal_941, \LED_128_Instance/addroundkey_out [42]}), .I2 ({IN_plaintext_s1[42], IN_plaintext_s0[42]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1405, \LED_128_Instance/state [42]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[43].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1316, \LED_128_Instance/mixcolumns_out [43]}), .I1 ({new_AGEMA_signal_937, \LED_128_Instance/addroundkey_out [43]}), .I2 ({IN_plaintext_s1[43], IN_plaintext_s0[43]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1407, \LED_128_Instance/state [43]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[44].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1330, \LED_128_Instance/mixcolumns_out [44]}), .I1 ({new_AGEMA_signal_933, \LED_128_Instance/addroundkey_out [44]}), .I2 ({IN_plaintext_s1[44], IN_plaintext_s0[44]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1409, \LED_128_Instance/state [44]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[45].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1326, \LED_128_Instance/mixcolumns_out [45]}), .I1 ({new_AGEMA_signal_929, \LED_128_Instance/addroundkey_out [45]}), .I2 ({IN_plaintext_s1[45], IN_plaintext_s0[45]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1411, \LED_128_Instance/state [45]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[46].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1329, \LED_128_Instance/mixcolumns_out [46]}), .I1 ({new_AGEMA_signal_925, \LED_128_Instance/addroundkey_out [46]}), .I2 ({IN_plaintext_s1[46], IN_plaintext_s0[46]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1413, \LED_128_Instance/state [46]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[47].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1325, \LED_128_Instance/mixcolumns_out [47]}), .I1 ({new_AGEMA_signal_921, \LED_128_Instance/addroundkey_out [47]}), .I2 ({IN_plaintext_s1[47], IN_plaintext_s0[47]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1415, \LED_128_Instance/state [47]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[48].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1301, \LED_128_Instance/mixcolumns_out [48]}), .I1 ({new_AGEMA_signal_1077, \LED_128_Instance/addroundkey_out [48]}), .I2 ({IN_plaintext_s1[48], IN_plaintext_s0[48]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1417, \LED_128_Instance/state [48]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[49].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1300, \LED_128_Instance/mixcolumns_out [49]}), .I1 ({new_AGEMA_signal_1073, \LED_128_Instance/addroundkey_out [49]}), .I2 ({IN_plaintext_s1[49], IN_plaintext_s0[49]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1419, \LED_128_Instance/state [49]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[50].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1201, \LED_128_Instance/mixcolumns_out [50]}), .I1 ({new_AGEMA_signal_917, \LED_128_Instance/addroundkey_out [50]}), .I2 ({IN_plaintext_s1[50], IN_plaintext_s0[50]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1289, \LED_128_Instance/state [50]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[51].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1335, \LED_128_Instance/mixcolumns_out [51]}), .I1 ({new_AGEMA_signal_913, \LED_128_Instance/addroundkey_out [51]}), .I2 ({IN_plaintext_s1[51], IN_plaintext_s0[51]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1421, \LED_128_Instance/state [51]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[52].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1310, \LED_128_Instance/mixcolumns_out [52]}), .I1 ({new_AGEMA_signal_1065, \LED_128_Instance/addroundkey_out [52]}), .I2 ({IN_plaintext_s1[52], IN_plaintext_s0[52]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1423, \LED_128_Instance/state [52]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[53].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1309, \LED_128_Instance/mixcolumns_out [53]}), .I1 ({new_AGEMA_signal_1061, \LED_128_Instance/addroundkey_out [53]}), .I2 ({IN_plaintext_s1[53], IN_plaintext_s0[53]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1425, \LED_128_Instance/state [53]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[54].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1205, \LED_128_Instance/mixcolumns_out [54]}), .I1 ({new_AGEMA_signal_1057, \LED_128_Instance/addroundkey_out [54]}), .I2 ({IN_plaintext_s1[54], IN_plaintext_s0[54]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1291, \LED_128_Instance/state [54]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[55].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1337, \LED_128_Instance/mixcolumns_out [55]}), .I1 ({new_AGEMA_signal_909, \LED_128_Instance/addroundkey_out [55]}), .I2 ({IN_plaintext_s1[55], IN_plaintext_s0[55]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1427, \LED_128_Instance/state [55]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[56].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1319, \LED_128_Instance/mixcolumns_out [56]}), .I1 ({new_AGEMA_signal_905, \LED_128_Instance/addroundkey_out [56]}), .I2 ({IN_plaintext_s1[56], IN_plaintext_s0[56]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1429, \LED_128_Instance/state [56]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[57].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1318, \LED_128_Instance/mixcolumns_out [57]}), .I1 ({new_AGEMA_signal_901, \LED_128_Instance/addroundkey_out [57]}), .I2 ({IN_plaintext_s1[57], IN_plaintext_s0[57]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1431, \LED_128_Instance/state [57]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[58].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1208, \LED_128_Instance/mixcolumns_out [58]}), .I1 ({new_AGEMA_signal_897, \LED_128_Instance/addroundkey_out [58]}), .I2 ({IN_plaintext_s1[58], IN_plaintext_s0[58]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1293, \LED_128_Instance/state [58]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[59].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1339, \LED_128_Instance/mixcolumns_out [59]}), .I1 ({new_AGEMA_signal_893, \LED_128_Instance/addroundkey_out [59]}), .I2 ({IN_plaintext_s1[59], IN_plaintext_s0[59]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1433, \LED_128_Instance/state [59]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[60].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1328, \LED_128_Instance/mixcolumns_out [60]}), .I1 ({new_AGEMA_signal_889, \LED_128_Instance/addroundkey_out [60]}), .I2 ({IN_plaintext_s1[60], IN_plaintext_s0[60]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1435, \LED_128_Instance/state [60]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[61].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1327, \LED_128_Instance/mixcolumns_out [61]}), .I1 ({new_AGEMA_signal_885, \LED_128_Instance/addroundkey_out [61]}), .I2 ({IN_plaintext_s1[61], IN_plaintext_s0[61]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1437, \LED_128_Instance/state [61]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[62].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1212, \LED_128_Instance/mixcolumns_out [62]}), .I1 ({new_AGEMA_signal_881, \LED_128_Instance/addroundkey_out [62]}), .I2 ({IN_plaintext_s1[62], IN_plaintext_s0[62]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1295, \LED_128_Instance/state [62]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'hF0F0CCAA ) , .MASK ( 5'b11000 ), .INIT2 ( 32'hF0F0CCAA ) ) \LED_128_Instance/MUX_state/gen_mux[63].mux_inst/LUTINST ( .I0 ({new_AGEMA_signal_1333, \LED_128_Instance/mixcolumns_out [63]}), .I1 ({new_AGEMA_signal_877, \LED_128_Instance/addroundkey_out [63]}), .I2 ({IN_plaintext_s1[63], IN_plaintext_s0[63]}), .I3 ({1'b0, \LED_128_Instance/roundconstant_001001 }), .I4 ({1'b0, IN_reset}), .O ({new_AGEMA_signal_1439, \LED_128_Instance/state [63]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<2>1 ( .I0 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I1 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I2 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I3 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I4 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .O ({new_AGEMA_signal_1200, \LED_128_Instance/mixcolumns_out [2]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<50>1 ( .I0 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I1 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I2 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I4 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .I5 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .O ({new_AGEMA_signal_1201, \LED_128_Instance/mixcolumns_out [50]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<3>1 ( .I0 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I1 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I2 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I3 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .O ({new_AGEMA_signal_1202, \LED_128_Instance/mixcolumns_out [3]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<0>1 ( .I0 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I3 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .O ({new_AGEMA_signal_1203, \LED_128_Instance/mixcolumns_out [0]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<6>1 ( .I0 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I1 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I2 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I3 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I4 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .O ({new_AGEMA_signal_1204, \LED_128_Instance/mixcolumns_out [6]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<54>1 ( .I0 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I1 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I2 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I3 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I4 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I5 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .O ({new_AGEMA_signal_1205, \LED_128_Instance/mixcolumns_out [54]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<7>1 ( .I0 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I1 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I2 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I3 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .O ({new_AGEMA_signal_1206, \LED_128_Instance/mixcolumns_out [7]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<4>1 ( .I0 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I1 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I3 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .O ({new_AGEMA_signal_1207, \LED_128_Instance/mixcolumns_out [4]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<58>1 ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I2 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .I3 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I4 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I5 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .O ({new_AGEMA_signal_1208, \LED_128_Instance/mixcolumns_out [58]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<10>1 ( .I0 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I1 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I2 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I3 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I4 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .O ({new_AGEMA_signal_1209, \LED_128_Instance/mixcolumns_out [10]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<8>1 ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I2 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I3 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .O ({new_AGEMA_signal_1210, \LED_128_Instance/mixcolumns_out [8]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<11>1 ( .I0 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I1 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I2 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I3 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .O ({new_AGEMA_signal_1211, \LED_128_Instance/mixcolumns_out [11]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<62>1 ( .I0 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I1 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I2 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I3 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I4 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I5 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1212, \LED_128_Instance/mixcolumns_out [62]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h96696996 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<14>1 ( .I0 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I1 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I2 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I3 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I4 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1213, \LED_128_Instance/mixcolumns_out [14]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<15>1 ( .I0 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I1 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I2 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I3 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1214, \LED_128_Instance/mixcolumns_out [15]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<12>1 ( .I0 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I1 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I2 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I3 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .O ({new_AGEMA_signal_1215, \LED_128_Instance/mixcolumns_out [12]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<19>_SW0 ( .I0 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I1 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I2 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .O ({new_AGEMA_signal_1216, N2}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<19> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I2 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I3 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I4 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I5 ({new_AGEMA_signal_1216, N2}), .O ({new_AGEMA_signal_1296, \LED_128_Instance/mixcolumns_out [19]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<16>_SW0 ( .I0 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I1 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1217, N4}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<16> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I2 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .I3 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I4 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I5 ({new_AGEMA_signal_1217, N4}), .O ({new_AGEMA_signal_1297, \LED_128_Instance/mixcolumns_out [16]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<35>_SW0 ( .I0 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I1 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I2 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I3 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I4 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1218, N6}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<35> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I2 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I3 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I4 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I5 ({new_AGEMA_signal_1218, N6}), .O ({new_AGEMA_signal_1298, \LED_128_Instance/mixcolumns_out [35]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<33>_SW0 ( .I0 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I4 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1219, N8}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<33> ( .I0 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I1 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I2 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I3 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I4 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I5 ({new_AGEMA_signal_1219, N8}), .O ({new_AGEMA_signal_1299, \LED_128_Instance/mixcolumns_out [33]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<49>_SW0 ( .I0 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I1 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I2 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1220, N12}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<49> ( .I0 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I1 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I2 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I3 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I4 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I5 ({new_AGEMA_signal_1220, N12}), .O ({new_AGEMA_signal_1300, \LED_128_Instance/mixcolumns_out [49]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<48>_SW0 ( .I0 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I1 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .I2 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I3 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .O ({new_AGEMA_signal_1221, N14}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<48> ( .I0 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I1 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I2 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I3 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I4 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I5 ({new_AGEMA_signal_1221, N14}), .O ({new_AGEMA_signal_1301, \LED_128_Instance/mixcolumns_out [48]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<34>_SW0 ( .I0 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .O ({new_AGEMA_signal_1222, N16}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<34> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I2 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I3 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I4 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .I5 ({new_AGEMA_signal_1222, N16}), .O ({new_AGEMA_signal_1302, \LED_128_Instance/mixcolumns_out [34]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<32>_SW0 ( .I0 ({new_AGEMA_signal_1136, \LED_128_Instance/subcells_out [0]}), .I1 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I2 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I4 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .O ({new_AGEMA_signal_1223, N18}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<32> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I2 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I3 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I4 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .I5 ({new_AGEMA_signal_1223, N18}), .O ({new_AGEMA_signal_1303, \LED_128_Instance/mixcolumns_out [32]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<17>_SW0 ( .I0 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I3 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .O ({new_AGEMA_signal_1224, N20}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<17> ( .I0 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I1 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I2 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I3 ({new_AGEMA_signal_1137, \LED_128_Instance/subcells_out [1]}), .I4 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I5 ({new_AGEMA_signal_1224, N20}), .O ({new_AGEMA_signal_1304, \LED_128_Instance/mixcolumns_out [17]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<23>_SW0 ( .I0 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I1 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I2 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1225, N22}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<23> ( .I0 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I1 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I2 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I3 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I4 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I5 ({new_AGEMA_signal_1225, N22}), .O ({new_AGEMA_signal_1305, \LED_128_Instance/mixcolumns_out [23]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<20>_SW0 ( .I0 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I1 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .O ({new_AGEMA_signal_1226, N24}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<20> ( .I0 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .I1 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I2 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I3 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I4 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I5 ({new_AGEMA_signal_1226, N24}), .O ({new_AGEMA_signal_1306, \LED_128_Instance/mixcolumns_out [20]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<39>_SW0 ( .I0 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I1 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I3 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1227, N26}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<39> ( .I0 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I1 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I2 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I3 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I4 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I5 ({new_AGEMA_signal_1227, N26}), .O ({new_AGEMA_signal_1307, \LED_128_Instance/mixcolumns_out [39]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<37>_SW0 ( .I0 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I1 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I3 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1228, N28}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<37> ( .I0 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I1 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I2 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I3 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I4 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I5 ({new_AGEMA_signal_1228, N28}), .O ({new_AGEMA_signal_1308, \LED_128_Instance/mixcolumns_out [37]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<53>_SW0 ( .I0 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I1 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .O ({new_AGEMA_signal_1229, N32}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<53> ( .I0 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I1 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I2 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I3 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I4 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I5 ({new_AGEMA_signal_1229, N32}), .O ({new_AGEMA_signal_1309, \LED_128_Instance/mixcolumns_out [53]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<52>_SW0 ( .I0 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I1 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I2 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I3 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1230, N34}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<52> ( .I0 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I1 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I2 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I3 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I4 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I5 ({new_AGEMA_signal_1230, N34}), .O ({new_AGEMA_signal_1310, \LED_128_Instance/mixcolumns_out [52]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<38>_SW0 ( .I0 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I1 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I2 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I3 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1231, N36}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<38> ( .I0 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .I1 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I2 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I3 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I4 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I5 ({new_AGEMA_signal_1231, N36}), .O ({new_AGEMA_signal_1311, \LED_128_Instance/mixcolumns_out [38]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<36>_SW0 ( .I0 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I1 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I2 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I3 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1232, N38}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<36> ( .I0 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .I1 ({new_AGEMA_signal_1140, \LED_128_Instance/subcells_out [4]}), .I2 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I3 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I4 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I5 ({new_AGEMA_signal_1232, N38}), .O ({new_AGEMA_signal_1312, \LED_128_Instance/mixcolumns_out [36]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<21>_SW0 ( .I0 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I1 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .I2 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I3 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .O ({new_AGEMA_signal_1233, N40}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<21> ( .I0 ({new_AGEMA_signal_1141, \LED_128_Instance/subcells_out [5]}), .I1 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I2 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I3 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I4 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I5 ({new_AGEMA_signal_1233, N40}), .O ({new_AGEMA_signal_1313, \LED_128_Instance/mixcolumns_out [21]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<24>_SW0 ( .I0 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I1 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .O ({new_AGEMA_signal_1234, N42}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<24> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I2 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I3 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I4 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .I5 ({new_AGEMA_signal_1234, N42}), .O ({new_AGEMA_signal_1314, \LED_128_Instance/mixcolumns_out [24]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<27>_SW0 ( .I0 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I1 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I2 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1235, N44}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<27> ( .I0 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I1 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I2 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I3 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I4 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I5 ({new_AGEMA_signal_1235, N44}), .O ({new_AGEMA_signal_1315, \LED_128_Instance/mixcolumns_out [27]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<43>_SW0 ( .I0 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I1 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I2 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .I3 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I4 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1236, N46}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<43> ( .I0 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I1 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I2 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I3 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I4 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I5 ({new_AGEMA_signal_1236, N46}), .O ({new_AGEMA_signal_1316, \LED_128_Instance/mixcolumns_out [43]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<41>_SW0 ( .I0 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I1 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I2 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I3 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .I4 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1237, N48}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<41> ( .I0 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I1 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I2 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I3 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I4 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I5 ({new_AGEMA_signal_1237, N48}), .O ({new_AGEMA_signal_1317, \LED_128_Instance/mixcolumns_out [41]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<57>_SW0 ( .I0 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I1 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I2 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .O ({new_AGEMA_signal_1238, N52}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<57> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I2 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I3 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I4 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I5 ({new_AGEMA_signal_1238, N52}), .O ({new_AGEMA_signal_1318, \LED_128_Instance/mixcolumns_out [57]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<56>_SW0 ( .I0 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I1 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I2 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I3 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .O ({new_AGEMA_signal_1239, N54}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<56> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I2 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I3 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I4 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I5 ({new_AGEMA_signal_1239, N54}), .O ({new_AGEMA_signal_1319, \LED_128_Instance/mixcolumns_out [56]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<42>_SW0 ( .I0 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I1 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I2 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I3 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1240, N56}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<42> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I2 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I3 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I4 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .I5 ({new_AGEMA_signal_1240, N56}), .O ({new_AGEMA_signal_1320, \LED_128_Instance/mixcolumns_out [42]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<40>_SW0 ( .I0 ({new_AGEMA_signal_1144, \LED_128_Instance/subcells_out [8]}), .I1 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I2 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I3 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I4 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .O ({new_AGEMA_signal_1241, N58}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<40> ( .I0 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I1 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I2 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I3 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I4 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .I5 ({new_AGEMA_signal_1241, N58}), .O ({new_AGEMA_signal_1321, \LED_128_Instance/mixcolumns_out [40]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<25>_SW0 ( .I0 ({new_AGEMA_signal_1145, \LED_128_Instance/subcells_out [9]}), .I1 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I2 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .I3 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .O ({new_AGEMA_signal_1242, N60}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<25> ( .I0 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I1 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I2 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I3 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I4 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I5 ({new_AGEMA_signal_1242, N60}), .O ({new_AGEMA_signal_1322, \LED_128_Instance/mixcolumns_out [25]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<28>_SW0 ( .I0 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I1 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1243, N62}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<28> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I2 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I3 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I4 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I5 ({new_AGEMA_signal_1243, N62}), .O ({new_AGEMA_signal_1323, \LED_128_Instance/mixcolumns_out [28]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<31>_SW0 ( .I0 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I1 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I2 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1244, N64}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<31> ( .I0 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I1 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I2 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I3 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I4 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I5 ({new_AGEMA_signal_1244, N64}), .O ({new_AGEMA_signal_1324, \LED_128_Instance/mixcolumns_out [31]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<47>_SW0 ( .I0 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I1 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I2 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I3 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .I4 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1245, N66}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<47> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I4 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I5 ({new_AGEMA_signal_1245, N66}), .O ({new_AGEMA_signal_1325, \LED_128_Instance/mixcolumns_out [47]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<45>_SW0 ( .I0 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I1 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I2 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I3 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .I4 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1246, N68}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<45> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I4 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I5 ({new_AGEMA_signal_1246, N68}), .O ({new_AGEMA_signal_1326, \LED_128_Instance/mixcolumns_out [45]}) ) ;
    LUT3_masked #(.low_latency(1), .pipeline(0),  .INIT ( 8'h69 ) , .MASK ( 3'b000 ), .INIT2 ( 8'h96 ) ) \LED_128_Instance/mixcolumns_out<61>_SW0 ( .I0 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I1 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I2 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1247, N72}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<61> ( .I0 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I1 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I2 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I3 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I4 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I5 ({new_AGEMA_signal_1247, N72}), .O ({new_AGEMA_signal_1327, \LED_128_Instance/mixcolumns_out [61]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<60>_SW0 ( .I0 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I1 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I2 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I3 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .O ({new_AGEMA_signal_1248, N74}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<60> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I4 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I5 ({new_AGEMA_signal_1248, N74}), .O ({new_AGEMA_signal_1328, \LED_128_Instance/mixcolumns_out [60]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<46>_SW0 ( .I0 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I1 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I2 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I3 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1249, N76}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<46> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I2 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I3 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I4 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I5 ({new_AGEMA_signal_1249, N76}), .O ({new_AGEMA_signal_1329, \LED_128_Instance/mixcolumns_out [46]}) ) ;
    LUT5_masked #(.low_latency(1), .pipeline(0),  .INIT ( 32'h69969669 ) , .MASK ( 5'b00000 ), .INIT2 ( 32'h96696996 ) ) \LED_128_Instance/mixcolumns_out<44>_SW0 ( .I0 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I1 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I2 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I3 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .I4 ({new_AGEMA_signal_1148, \LED_128_Instance/subcells_out [12]}), .O ({new_AGEMA_signal_1250, N78}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h9669699669969669 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<44> ( .I0 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I1 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I2 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I3 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I4 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I5 ({new_AGEMA_signal_1250, N78}), .O ({new_AGEMA_signal_1330, \LED_128_Instance/mixcolumns_out [44]}) ) ;
    LUT4_masked #(.low_latency(1), .pipeline(0),  .INIT ( 16'h6996 ) , .MASK ( 4'b0000 ), .INIT2 ( 16'h6996 ) ) \LED_128_Instance/mixcolumns_out<29>_SW0 ( .I0 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I1 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I2 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .I3 ({new_AGEMA_signal_1149, \LED_128_Instance/subcells_out [13]}), .O ({new_AGEMA_signal_1251, N80}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<29> ( .I0 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I1 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I2 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I3 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .I4 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I5 ({new_AGEMA_signal_1251, N80}), .O ({new_AGEMA_signal_1331, \LED_128_Instance/mixcolumns_out [29]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<13>31_SW0 ( .I0 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I1 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .O ({new_AGEMA_signal_1252, N82}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<13>1 ( .I0 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I1 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I4 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I5 ({new_AGEMA_signal_1252, N82}), .O ({new_AGEMA_signal_1332, \LED_128_Instance/mixcolumns_out [13]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<13>31_SW1 ( .I0 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I1 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .O ({new_AGEMA_signal_1253, N84}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<63>1 ( .I0 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I1 ({new_AGEMA_signal_1154, \LED_128_Instance/subcells_out [18]}), .I2 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I3 ({new_AGEMA_signal_1173, \LED_128_Instance/subcells_out [37]}), .I4 ({new_AGEMA_signal_1194, \LED_128_Instance/subcells_out [58]}), .I5 ({new_AGEMA_signal_1253, N84}), .O ({new_AGEMA_signal_1333, \LED_128_Instance/mixcolumns_out [63]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<18>41_SW0 ( .I0 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I1 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1254, N86}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<1>1 ( .I0 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I1 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .I2 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I3 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I4 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I5 ({new_AGEMA_signal_1254, N86}), .O ({new_AGEMA_signal_1334, \LED_128_Instance/mixcolumns_out [1]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<18>41_SW1 ( .I0 ({new_AGEMA_signal_1177, \LED_128_Instance/subcells_out [41]}), .I1 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .O ({new_AGEMA_signal_1255, N88}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<51>1 ( .I0 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I1 ({new_AGEMA_signal_1158, \LED_128_Instance/subcells_out [22]}), .I2 ({new_AGEMA_signal_1198, \LED_128_Instance/subcells_out [62]}), .I3 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I4 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I5 ({new_AGEMA_signal_1255, N88}), .O ({new_AGEMA_signal_1335, \LED_128_Instance/mixcolumns_out [51]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<22>41_SW0 ( .I0 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I1 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .O ({new_AGEMA_signal_1256, N90}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<5>1 ( .I0 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I1 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .I2 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I3 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .I5 ({new_AGEMA_signal_1256, N90}), .O ({new_AGEMA_signal_1336, \LED_128_Instance/mixcolumns_out [5]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<22>41_SW1 ( .I0 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I1 ({new_AGEMA_signal_1162, \LED_128_Instance/subcells_out [26]}), .O ({new_AGEMA_signal_1257, N92}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<55>1 ( .I0 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I1 ({new_AGEMA_signal_1186, \LED_128_Instance/subcells_out [50]}), .I2 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I3 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I4 ({new_AGEMA_signal_1181, \LED_128_Instance/subcells_out [45]}), .I5 ({new_AGEMA_signal_1257, N92}), .O ({new_AGEMA_signal_1337, \LED_128_Instance/mixcolumns_out [55]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<26>41_SW0 ( .I0 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I1 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .O ({new_AGEMA_signal_1258, N94}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<9>1 ( .I0 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I1 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I2 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I3 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I4 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .I5 ({new_AGEMA_signal_1258, N94}), .O ({new_AGEMA_signal_1338, \LED_128_Instance/mixcolumns_out [9]}) ) ;
    LUT2_masked #(.low_latency(1), .pipeline(0),  .INIT ( 4'h6 ) , .MASK ( 2'b00 ), .INIT2 ( 4'h6 ) ) \LED_128_Instance/mixcolumns_out<26>41_SW1 ( .I0 ({new_AGEMA_signal_1166, \LED_128_Instance/subcells_out [30]}), .I1 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .O ({new_AGEMA_signal_1259, N96}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<59>1 ( .I0 ({new_AGEMA_signal_1169, \LED_128_Instance/subcells_out [33]}), .I1 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I2 ({new_AGEMA_signal_1190, \LED_128_Instance/subcells_out [54]}), .I3 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I4 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .I5 ({new_AGEMA_signal_1259, N96}), .O ({new_AGEMA_signal_1339, \LED_128_Instance/mixcolumns_out [59]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<18>_SW1 ( .I0 ({new_AGEMA_signal_1196, \LED_128_Instance/subcells_out [60]}), .I1 ({new_AGEMA_signal_1179, \LED_128_Instance/subcells_out [43]}), .I2 ({new_AGEMA_signal_1178, \LED_128_Instance/subcells_out [42]}), .I3 ({new_AGEMA_signal_1176, \LED_128_Instance/subcells_out [40]}), .I4 ({new_AGEMA_signal_1138, \LED_128_Instance/subcells_out [2]}), .I5 ({new_AGEMA_signal_1139, \LED_128_Instance/subcells_out [3]}), .O ({new_AGEMA_signal_1260, N98}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<18> ( .I0 ({new_AGEMA_signal_1159, \LED_128_Instance/subcells_out [23]}), .I1 ({new_AGEMA_signal_1157, \LED_128_Instance/subcells_out [21]}), .I2 ({new_AGEMA_signal_1156, \LED_128_Instance/subcells_out [20]}), .I3 ({new_AGEMA_signal_1199, \LED_128_Instance/subcells_out [63]}), .I4 ({new_AGEMA_signal_1197, \LED_128_Instance/subcells_out [61]}), .I5 ({new_AGEMA_signal_1260, N98}), .O ({new_AGEMA_signal_1340, \LED_128_Instance/mixcolumns_out [18]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<22>_SW1 ( .I0 ({new_AGEMA_signal_1182, \LED_128_Instance/subcells_out [46]}), .I1 ({new_AGEMA_signal_1180, \LED_128_Instance/subcells_out [44]}), .I2 ({new_AGEMA_signal_1163, \LED_128_Instance/subcells_out [27]}), .I3 ({new_AGEMA_signal_1161, \LED_128_Instance/subcells_out [25]}), .I4 ({new_AGEMA_signal_1160, \LED_128_Instance/subcells_out [24]}), .I5 ({new_AGEMA_signal_1143, \LED_128_Instance/subcells_out [7]}), .O ({new_AGEMA_signal_1261, N100}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<22> ( .I0 ({new_AGEMA_signal_1187, \LED_128_Instance/subcells_out [51]}), .I1 ({new_AGEMA_signal_1185, \LED_128_Instance/subcells_out [49]}), .I2 ({new_AGEMA_signal_1184, \LED_128_Instance/subcells_out [48]}), .I3 ({new_AGEMA_signal_1142, \LED_128_Instance/subcells_out [6]}), .I4 ({new_AGEMA_signal_1183, \LED_128_Instance/subcells_out [47]}), .I5 ({new_AGEMA_signal_1261, N100}), .O ({new_AGEMA_signal_1341, \LED_128_Instance/mixcolumns_out [22]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<26>_SW1 ( .I0 ({new_AGEMA_signal_1167, \LED_128_Instance/subcells_out [31]}), .I1 ({new_AGEMA_signal_1165, \LED_128_Instance/subcells_out [29]}), .I2 ({new_AGEMA_signal_1164, \LED_128_Instance/subcells_out [28]}), .I3 ({new_AGEMA_signal_1147, \LED_128_Instance/subcells_out [11]}), .I4 ({new_AGEMA_signal_1146, \LED_128_Instance/subcells_out [10]}), .I5 ({new_AGEMA_signal_1170, \LED_128_Instance/subcells_out [34]}), .O ({new_AGEMA_signal_1262, N102}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<26> ( .I0 ({new_AGEMA_signal_1191, \LED_128_Instance/subcells_out [55]}), .I1 ({new_AGEMA_signal_1189, \LED_128_Instance/subcells_out [53]}), .I2 ({new_AGEMA_signal_1188, \LED_128_Instance/subcells_out [52]}), .I3 ({new_AGEMA_signal_1171, \LED_128_Instance/subcells_out [35]}), .I4 ({new_AGEMA_signal_1168, \LED_128_Instance/subcells_out [32]}), .I5 ({new_AGEMA_signal_1262, N102}), .O ({new_AGEMA_signal_1342, \LED_128_Instance/mixcolumns_out [26]}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<30>_SW1 ( .I0 ({new_AGEMA_signal_1151, \LED_128_Instance/subcells_out [15]}), .I1 ({new_AGEMA_signal_1150, \LED_128_Instance/subcells_out [14]}), .I2 ({new_AGEMA_signal_1175, \LED_128_Instance/subcells_out [39]}), .I3 ({new_AGEMA_signal_1174, \LED_128_Instance/subcells_out [38]}), .I4 ({new_AGEMA_signal_1155, \LED_128_Instance/subcells_out [19]}), .I5 ({new_AGEMA_signal_1152, \LED_128_Instance/subcells_out [16]}), .O ({new_AGEMA_signal_1263, N104}) ) ;
    LUT6_masked #(.low_latency(1), .pipeline(0),  .INIT ( 64'h6996966996696996 ) , .MASK ( 6'b000000 ), .INIT2 ( 64'h6996966996696996 ) ) \LED_128_Instance/mixcolumns_out<30> ( .I0 ({new_AGEMA_signal_1195, \LED_128_Instance/subcells_out [59]}), .I1 ({new_AGEMA_signal_1193, \LED_128_Instance/subcells_out [57]}), .I2 ({new_AGEMA_signal_1192, \LED_128_Instance/subcells_out [56]}), .I3 ({new_AGEMA_signal_1172, \LED_128_Instance/subcells_out [36]}), .I4 ({new_AGEMA_signal_1153, \LED_128_Instance/subcells_out [17]}), .I5 ({new_AGEMA_signal_1263, N104}), .O ({new_AGEMA_signal_1343, \LED_128_Instance/mixcolumns_out [30]}) ) ;

    /* register cells */
    FDR \LED_128_Instance/roundconstant_5 ( .D (\LED_128_Instance/roundconstant [4]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [5]) ) ;
    FDR \LED_128_Instance/roundconstant_4 ( .D (\LED_128_Instance/roundconstant [3]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [4]) ) ;
    FDR \LED_128_Instance/roundconstant_3 ( .D (\LED_128_Instance/roundconstant [2]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [3]) ) ;
    FDR \LED_128_Instance/roundconstant_2 ( .D (\LED_128_Instance/roundconstant [1]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [2]) ) ;
    FDR \LED_128_Instance/roundconstant_1 ( .D (\LED_128_Instance/roundconstant [0]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/roundconstant [1]) ) ;
    FDS \LED_128_Instance/roundconstant_0 ( .D (\LED_128_Instance/roundconstant[5]_roundconstant[4]_XOR_7_o ), .C (clk_gated), .S (IN_reset), .Q (\LED_128_Instance/roundconstant [0]) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_63 ( .D ({new_AGEMA_signal_1439, \LED_128_Instance/state [63]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[63], OUT_ciphertext_s0[63]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_62 ( .D ({new_AGEMA_signal_1295, \LED_128_Instance/state [62]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[62], OUT_ciphertext_s0[62]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_61 ( .D ({new_AGEMA_signal_1437, \LED_128_Instance/state [61]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[61], OUT_ciphertext_s0[61]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_60 ( .D ({new_AGEMA_signal_1435, \LED_128_Instance/state [60]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[60], OUT_ciphertext_s0[60]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_59 ( .D ({new_AGEMA_signal_1433, \LED_128_Instance/state [59]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[59], OUT_ciphertext_s0[59]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_58 ( .D ({new_AGEMA_signal_1293, \LED_128_Instance/state [58]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[58], OUT_ciphertext_s0[58]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_57 ( .D ({new_AGEMA_signal_1431, \LED_128_Instance/state [57]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[57], OUT_ciphertext_s0[57]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_56 ( .D ({new_AGEMA_signal_1429, \LED_128_Instance/state [56]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[56], OUT_ciphertext_s0[56]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_55 ( .D ({new_AGEMA_signal_1427, \LED_128_Instance/state [55]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[55], OUT_ciphertext_s0[55]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_54 ( .D ({new_AGEMA_signal_1291, \LED_128_Instance/state [54]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[54], OUT_ciphertext_s0[54]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_53 ( .D ({new_AGEMA_signal_1425, \LED_128_Instance/state [53]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[53], OUT_ciphertext_s0[53]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_52 ( .D ({new_AGEMA_signal_1423, \LED_128_Instance/state [52]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[52], OUT_ciphertext_s0[52]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_51 ( .D ({new_AGEMA_signal_1421, \LED_128_Instance/state [51]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[51], OUT_ciphertext_s0[51]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_50 ( .D ({new_AGEMA_signal_1289, \LED_128_Instance/state [50]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[50], OUT_ciphertext_s0[50]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_49 ( .D ({new_AGEMA_signal_1419, \LED_128_Instance/state [49]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[49], OUT_ciphertext_s0[49]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_48 ( .D ({new_AGEMA_signal_1417, \LED_128_Instance/state [48]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[48], OUT_ciphertext_s0[48]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_47 ( .D ({new_AGEMA_signal_1415, \LED_128_Instance/state [47]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[47], OUT_ciphertext_s0[47]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_46 ( .D ({new_AGEMA_signal_1413, \LED_128_Instance/state [46]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[46], OUT_ciphertext_s0[46]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_45 ( .D ({new_AGEMA_signal_1411, \LED_128_Instance/state [45]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[45], OUT_ciphertext_s0[45]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_44 ( .D ({new_AGEMA_signal_1409, \LED_128_Instance/state [44]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[44], OUT_ciphertext_s0[44]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_43 ( .D ({new_AGEMA_signal_1407, \LED_128_Instance/state [43]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[43], OUT_ciphertext_s0[43]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_42 ( .D ({new_AGEMA_signal_1405, \LED_128_Instance/state [42]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[42], OUT_ciphertext_s0[42]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_41 ( .D ({new_AGEMA_signal_1403, \LED_128_Instance/state [41]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[41], OUT_ciphertext_s0[41]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_40 ( .D ({new_AGEMA_signal_1401, \LED_128_Instance/state [40]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[40], OUT_ciphertext_s0[40]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_39 ( .D ({new_AGEMA_signal_1399, \LED_128_Instance/state [39]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[39], OUT_ciphertext_s0[39]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_38 ( .D ({new_AGEMA_signal_1397, \LED_128_Instance/state [38]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[38], OUT_ciphertext_s0[38]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_37 ( .D ({new_AGEMA_signal_1395, \LED_128_Instance/state [37]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[37], OUT_ciphertext_s0[37]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_36 ( .D ({new_AGEMA_signal_1393, \LED_128_Instance/state [36]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[36], OUT_ciphertext_s0[36]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_35 ( .D ({new_AGEMA_signal_1391, \LED_128_Instance/state [35]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[35], OUT_ciphertext_s0[35]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_34 ( .D ({new_AGEMA_signal_1389, \LED_128_Instance/state [34]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[34], OUT_ciphertext_s0[34]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_33 ( .D ({new_AGEMA_signal_1387, \LED_128_Instance/state [33]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[33], OUT_ciphertext_s0[33]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_32 ( .D ({new_AGEMA_signal_1385, \LED_128_Instance/state [32]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[32], OUT_ciphertext_s0[32]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_31 ( .D ({new_AGEMA_signal_1383, \LED_128_Instance/state [31]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[31], OUT_ciphertext_s0[31]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_30 ( .D ({new_AGEMA_signal_1381, \LED_128_Instance/state [30]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[30], OUT_ciphertext_s0[30]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_29 ( .D ({new_AGEMA_signal_1379, \LED_128_Instance/state [29]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[29], OUT_ciphertext_s0[29]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_28 ( .D ({new_AGEMA_signal_1377, \LED_128_Instance/state [28]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[28], OUT_ciphertext_s0[28]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_27 ( .D ({new_AGEMA_signal_1375, \LED_128_Instance/state [27]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[27], OUT_ciphertext_s0[27]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_26 ( .D ({new_AGEMA_signal_1373, \LED_128_Instance/state [26]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[26], OUT_ciphertext_s0[26]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_25 ( .D ({new_AGEMA_signal_1371, \LED_128_Instance/state [25]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[25], OUT_ciphertext_s0[25]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_24 ( .D ({new_AGEMA_signal_1369, \LED_128_Instance/state [24]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[24], OUT_ciphertext_s0[24]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_23 ( .D ({new_AGEMA_signal_1367, \LED_128_Instance/state [23]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[23], OUT_ciphertext_s0[23]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_22 ( .D ({new_AGEMA_signal_1365, \LED_128_Instance/state [22]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[22], OUT_ciphertext_s0[22]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_21 ( .D ({new_AGEMA_signal_1363, \LED_128_Instance/state [21]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[21], OUT_ciphertext_s0[21]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_20 ( .D ({new_AGEMA_signal_1361, \LED_128_Instance/state [20]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[20], OUT_ciphertext_s0[20]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_19 ( .D ({new_AGEMA_signal_1359, \LED_128_Instance/state [19]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[19], OUT_ciphertext_s0[19]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_18 ( .D ({new_AGEMA_signal_1357, \LED_128_Instance/state [18]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[18], OUT_ciphertext_s0[18]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_17 ( .D ({new_AGEMA_signal_1355, \LED_128_Instance/state [17]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[17], OUT_ciphertext_s0[17]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_16 ( .D ({new_AGEMA_signal_1353, \LED_128_Instance/state [16]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[16], OUT_ciphertext_s0[16]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_15 ( .D ({new_AGEMA_signal_1287, \LED_128_Instance/state [15]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[15], OUT_ciphertext_s0[15]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_14 ( .D ({new_AGEMA_signal_1285, \LED_128_Instance/state [14]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[14], OUT_ciphertext_s0[14]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_13 ( .D ({new_AGEMA_signal_1351, \LED_128_Instance/state [13]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[13], OUT_ciphertext_s0[13]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_12 ( .D ({new_AGEMA_signal_1283, \LED_128_Instance/state [12]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[12], OUT_ciphertext_s0[12]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_11 ( .D ({new_AGEMA_signal_1281, \LED_128_Instance/state [11]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[11], OUT_ciphertext_s0[11]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_10 ( .D ({new_AGEMA_signal_1279, \LED_128_Instance/state [10]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[10], OUT_ciphertext_s0[10]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_9 ( .D ({new_AGEMA_signal_1349, \LED_128_Instance/state [9]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[9], OUT_ciphertext_s0[9]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_8 ( .D ({new_AGEMA_signal_1277, \LED_128_Instance/state [8]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[8], OUT_ciphertext_s0[8]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_7 ( .D ({new_AGEMA_signal_1275, \LED_128_Instance/state [7]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[7], OUT_ciphertext_s0[7]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_6 ( .D ({new_AGEMA_signal_1273, \LED_128_Instance/state [6]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[6], OUT_ciphertext_s0[6]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_5 ( .D ({new_AGEMA_signal_1347, \LED_128_Instance/state [5]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[5], OUT_ciphertext_s0[5]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_4 ( .D ({new_AGEMA_signal_1271, \LED_128_Instance/state [4]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[4], OUT_ciphertext_s0[4]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_3 ( .D ({new_AGEMA_signal_1269, \LED_128_Instance/state [3]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[3], OUT_ciphertext_s0[3]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_2 ( .D ({new_AGEMA_signal_1267, \LED_128_Instance/state [2]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[2], OUT_ciphertext_s0[2]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_1 ( .D ({new_AGEMA_signal_1345, \LED_128_Instance/state [1]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[1], OUT_ciphertext_s0[1]}) ) ;
    FD_masked #(.low_latency(1), .pipeline(0)) \LED_128_Instance/cipherstate_0 ( .D ({new_AGEMA_signal_1265, \LED_128_Instance/state [0]}), .clk (clk_gated), .Q ({OUT_ciphertext_s1[0], OUT_ciphertext_s0[0]}) ) ;
    FDR \LED_128_Instance/ks_3 ( .D (\LED_128_Instance/ks [2]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/ks [3]) ) ;
    FDR \LED_128_Instance/ks_2 ( .D (\LED_128_Instance/ks [1]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/ks [2]) ) ;
    FDR \LED_128_Instance/ks_1 ( .D (\LED_128_Instance/ks [0]), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/ks [1]) ) ;
    FDR \LED_128_Instance/ks_0 ( .D (\LED_128_Instance/ks[3]_INV_6_o ), .C (clk_gated), .R (IN_reset), .Q (\LED_128_Instance/ks [0]) ) ;
    FDR internal_done ( .D (internal_done_glue_set_843), .C (clk_gated), .R (IN_reset), .Q (OUT_done) ) ;
endmodule
